magic
tech sky130A
magscale 1 2
timestamp 1638470712
<< locali >>
rect 15577 5559 15611 5797
rect 213 3587 247 4029
rect 5089 2907 5123 3009
rect 4905 2499 4939 2601
rect 12265 1751 12299 1989
<< viali >>
rect 6837 10761 6871 10795
rect 10057 10761 10091 10795
rect 13737 10761 13771 10795
rect 18245 10761 18279 10795
rect 7481 10693 7515 10727
rect 8309 10693 8343 10727
rect 12817 10693 12851 10727
rect 17969 10693 18003 10727
rect 2329 10625 2363 10659
rect 2605 10625 2639 10659
rect 3157 10625 3191 10659
rect 5273 10625 5307 10659
rect 5457 10625 5491 10659
rect 6653 10625 6687 10659
rect 6929 10625 6963 10659
rect 7297 10625 7331 10659
rect 8861 10625 8895 10659
rect 10241 10625 10275 10659
rect 13921 10625 13955 10659
rect 17601 10625 17635 10659
rect 17877 10625 17911 10659
rect 18061 10625 18095 10659
rect 2881 10557 2915 10591
rect 8309 10557 8343 10591
rect 8401 10557 8435 10591
rect 12541 10557 12575 10591
rect 12725 10557 12759 10591
rect 3065 10489 3099 10523
rect 7849 10489 7883 10523
rect 17785 10489 17819 10523
rect 2237 10421 2271 10455
rect 2513 10421 2547 10455
rect 2973 10421 3007 10455
rect 5273 10421 5307 10455
rect 7113 10421 7147 10455
rect 8585 10421 8619 10455
rect 9505 10421 9539 10455
rect 11345 10421 11379 10455
rect 13185 10421 13219 10455
rect 14013 10421 14047 10455
rect 14933 10421 14967 10455
rect 1869 10217 1903 10251
rect 8585 10217 8619 10251
rect 10609 10217 10643 10251
rect 18015 10217 18049 10251
rect 9137 10149 9171 10183
rect 1685 10081 1719 10115
rect 2053 10081 2087 10115
rect 2421 10081 2455 10115
rect 4445 10081 4479 10115
rect 4721 10081 4755 10115
rect 5825 10081 5859 10115
rect 14013 10081 14047 10115
rect 16221 10081 16255 10115
rect 1961 10013 1995 10047
rect 4353 10013 4387 10047
rect 4813 10013 4847 10047
rect 5089 10013 5123 10047
rect 5641 10013 5675 10047
rect 5917 10013 5951 10047
rect 7205 10013 7239 10047
rect 7461 10013 7495 10047
rect 9321 10013 9355 10047
rect 11253 10013 11287 10047
rect 14381 10013 14415 10047
rect 15807 10013 15841 10047
rect 16589 10013 16623 10047
rect 11529 9945 11563 9979
rect 1685 9877 1719 9911
rect 3847 9877 3881 9911
rect 5365 9877 5399 9911
rect 6285 9877 6319 9911
rect 13001 9877 13035 9911
rect 13185 9877 13219 9911
rect 13921 9877 13955 9911
rect 16037 9877 16071 9911
rect 2513 9673 2547 9707
rect 3065 9673 3099 9707
rect 3249 9673 3283 9707
rect 6745 9673 6779 9707
rect 11529 9673 11563 9707
rect 14611 9673 14645 9707
rect 949 9605 983 9639
rect 2973 9605 3007 9639
rect 5641 9605 5675 9639
rect 10885 9605 10919 9639
rect 12449 9605 12483 9639
rect 12633 9605 12667 9639
rect 673 9537 707 9571
rect 2513 9537 2547 9571
rect 2697 9537 2731 9571
rect 2881 9537 2915 9571
rect 3157 9537 3191 9571
rect 3249 9537 3283 9571
rect 3433 9537 3467 9571
rect 3801 9537 3835 9571
rect 4721 9537 4755 9571
rect 4813 9537 4847 9571
rect 5733 9537 5767 9571
rect 6653 9537 6687 9571
rect 8760 9537 8794 9571
rect 11897 9537 11931 9571
rect 12817 9537 12851 9571
rect 18245 9537 18279 9571
rect 18521 9537 18555 9571
rect 2421 9469 2455 9503
rect 4997 9469 5031 9503
rect 5825 9469 5859 9503
rect 6469 9469 6503 9503
rect 8493 9469 8527 9503
rect 10609 9469 10643 9503
rect 10793 9469 10827 9503
rect 11989 9469 12023 9503
rect 12173 9469 12207 9503
rect 13185 9469 13219 9503
rect 14841 9469 14875 9503
rect 16589 9469 16623 9503
rect 16865 9469 16899 9503
rect 4353 9401 4387 9435
rect 5273 9401 5307 9435
rect 11253 9401 11287 9435
rect 3709 9333 3743 9367
rect 4077 9333 4111 9367
rect 4169 9333 4203 9367
rect 7113 9333 7147 9367
rect 9873 9333 9907 9367
rect 18337 9333 18371 9367
rect 1133 9129 1167 9163
rect 6469 9129 6503 9163
rect 10609 9129 10643 9163
rect 15853 9129 15887 9163
rect 1225 8993 1259 9027
rect 7021 8993 7055 9027
rect 8861 8993 8895 9027
rect 14105 8993 14139 9027
rect 16037 8993 16071 9027
rect 1409 8925 1443 8959
rect 1501 8925 1535 8959
rect 1685 8925 1719 8959
rect 3341 8925 3375 8959
rect 4077 8925 4111 8959
rect 4261 8925 4295 8959
rect 7297 8925 7331 8959
rect 11253 8925 11287 8959
rect 16405 8925 16439 8959
rect 2881 8857 2915 8891
rect 6837 8857 6871 8891
rect 7564 8857 7598 8891
rect 9137 8857 9171 8891
rect 11529 8857 11563 8891
rect 13277 8857 13311 8891
rect 14381 8857 14415 8891
rect 1225 8789 1259 8823
rect 3249 8789 3283 8823
rect 4169 8789 4203 8823
rect 6929 8789 6963 8823
rect 8677 8789 8711 8823
rect 11069 8789 11103 8823
rect 14013 8789 14047 8823
rect 18153 8789 18187 8823
rect 2881 8585 2915 8619
rect 4445 8585 4479 8619
rect 8217 8585 8251 8619
rect 8769 8585 8803 8619
rect 9597 8585 9631 8619
rect 11529 8585 11563 8619
rect 16635 8585 16669 8619
rect 949 8517 983 8551
rect 6101 8517 6135 8551
rect 18245 8517 18279 8551
rect 673 8449 707 8483
rect 2881 8449 2915 8483
rect 3065 8449 3099 8483
rect 3157 8449 3191 8483
rect 3433 8449 3467 8483
rect 5365 8449 5399 8483
rect 5549 8449 5583 8483
rect 5825 8449 5859 8483
rect 5917 8449 5951 8483
rect 6191 8471 6225 8505
rect 6285 8449 6319 8483
rect 6377 8449 6411 8483
rect 6561 8449 6595 8483
rect 8309 8449 8343 8483
rect 8861 8449 8895 8483
rect 9045 8449 9079 8483
rect 9321 8449 9355 8483
rect 9689 8449 9723 8483
rect 9873 8449 9907 8483
rect 10425 8449 10459 8483
rect 10977 8449 11011 8483
rect 11713 8449 11747 8483
rect 13838 8449 13872 8483
rect 14841 8449 14875 8483
rect 17969 8449 18003 8483
rect 2421 8381 2455 8415
rect 4261 8381 4295 8415
rect 4353 8381 4387 8415
rect 9597 8381 9631 8415
rect 10885 8381 10919 8415
rect 11989 8381 12023 8415
rect 14105 8381 14139 8415
rect 15209 8381 15243 8415
rect 2605 8313 2639 8347
rect 6193 8313 6227 8347
rect 6469 8313 6503 8347
rect 9229 8313 9263 8347
rect 9413 8313 9447 8347
rect 9873 8313 9907 8347
rect 16773 8313 16807 8347
rect 17785 8313 17819 8347
rect 18521 8313 18555 8347
rect 4813 8245 4847 8279
rect 5549 8245 5583 8279
rect 10517 8245 10551 8279
rect 11253 8245 11287 8279
rect 11437 8245 11471 8279
rect 11897 8245 11931 8279
rect 12725 8245 12759 8279
rect 14657 8245 14691 8279
rect 18153 8245 18187 8279
rect 4077 8041 4111 8075
rect 4905 8041 4939 8075
rect 5273 8041 5307 8075
rect 5641 8041 5675 8075
rect 2789 7973 2823 8007
rect 6285 7973 6319 8007
rect 14289 7973 14323 8007
rect 3801 7905 3835 7939
rect 4721 7905 4755 7939
rect 4997 7905 5031 7939
rect 5089 7905 5123 7939
rect 5457 7905 5491 7939
rect 7205 7905 7239 7939
rect 11253 7905 11287 7939
rect 14749 7905 14783 7939
rect 15669 7905 15703 7939
rect 16221 7905 16255 7939
rect 2053 7837 2087 7871
rect 2237 7837 2271 7871
rect 2605 7837 2639 7871
rect 2789 7837 2823 7871
rect 3709 7837 3743 7871
rect 4445 7837 4479 7871
rect 5365 7837 5399 7871
rect 5733 7837 5767 7871
rect 6837 7837 6871 7871
rect 11069 7837 11103 7871
rect 11621 7837 11655 7871
rect 13047 7837 13081 7871
rect 13645 7837 13679 7871
rect 14013 7837 14047 7871
rect 14197 7837 14231 7871
rect 14841 7837 14875 7871
rect 16037 7837 16071 7871
rect 4537 7769 4571 7803
rect 5457 7769 5491 7803
rect 5917 7769 5951 7803
rect 6469 7769 6503 7803
rect 6653 7769 6687 7803
rect 13277 7769 13311 7803
rect 13461 7769 13495 7803
rect 15577 7769 15611 7803
rect 16497 7769 16531 7803
rect 18245 7769 18279 7803
rect 2237 7701 2271 7735
rect 6009 7701 6043 7735
rect 8631 7701 8665 7735
rect 9781 7701 9815 7735
rect 13737 7701 13771 7735
rect 15117 7701 15151 7735
rect 15485 7701 15519 7735
rect 2605 7497 2639 7531
rect 2973 7497 3007 7531
rect 6561 7497 6595 7531
rect 7757 7497 7791 7531
rect 8861 7497 8895 7531
rect 9873 7497 9907 7531
rect 10885 7497 10919 7531
rect 11437 7497 11471 7531
rect 11897 7497 11931 7531
rect 13185 7497 13219 7531
rect 14565 7497 14599 7531
rect 14933 7497 14967 7531
rect 15301 7497 15335 7531
rect 7297 7429 7331 7463
rect 11161 7429 11195 7463
rect 11989 7429 12023 7463
rect 673 7361 707 7395
rect 2513 7361 2547 7395
rect 3065 7361 3099 7395
rect 3249 7361 3283 7395
rect 4905 7361 4939 7395
rect 5089 7361 5123 7395
rect 5641 7361 5675 7395
rect 6837 7361 6871 7395
rect 7021 7361 7055 7395
rect 7849 7361 7883 7395
rect 8769 7361 8803 7395
rect 9505 7361 9539 7395
rect 9689 7361 9723 7395
rect 10149 7361 10183 7395
rect 10241 7361 10275 7395
rect 10333 7361 10367 7395
rect 10609 7361 10643 7395
rect 10793 7361 10827 7395
rect 11345 7361 11379 7395
rect 11437 7361 11471 7395
rect 11713 7361 11747 7395
rect 11805 7361 11839 7395
rect 12817 7361 12851 7395
rect 14105 7361 14139 7395
rect 14197 7361 14231 7395
rect 14381 7361 14415 7395
rect 14473 7361 14507 7395
rect 14841 7361 14875 7395
rect 15025 7361 15059 7395
rect 17049 7361 17083 7395
rect 17417 7361 17451 7395
rect 949 7293 983 7327
rect 3801 7293 3835 7327
rect 5733 7293 5767 7327
rect 5825 7293 5859 7327
rect 6101 7293 6135 7327
rect 9045 7293 9079 7327
rect 9413 7293 9447 7327
rect 10517 7293 10551 7327
rect 12725 7293 12759 7327
rect 16773 7293 16807 7327
rect 3525 7225 3559 7259
rect 4905 7225 4939 7259
rect 7481 7225 7515 7259
rect 11069 7225 11103 7259
rect 2421 7157 2455 7191
rect 3341 7157 3375 7191
rect 5273 7157 5307 7191
rect 7021 7157 7055 7191
rect 8401 7157 8435 7191
rect 11621 7157 11655 7191
rect 14105 7157 14139 7191
rect 15117 7157 15151 7191
rect 17233 7157 17267 7191
rect 2421 6953 2455 6987
rect 9045 6953 9079 6987
rect 11253 6953 11287 6987
rect 1409 6885 1443 6919
rect 2881 6885 2915 6919
rect 3065 6885 3099 6919
rect 10885 6885 10919 6919
rect 15439 6885 15473 6919
rect 1225 6817 1259 6851
rect 5365 6817 5399 6851
rect 6745 6817 6779 6851
rect 7021 6817 7055 6851
rect 8125 6817 8159 6851
rect 9597 6817 9631 6851
rect 13645 6817 13679 6851
rect 16773 6817 16807 6851
rect 18199 6817 18233 6851
rect 949 6749 983 6783
rect 1501 6749 1535 6783
rect 1961 6749 1995 6783
rect 2053 6749 2087 6783
rect 2513 6749 2547 6783
rect 2973 6749 3007 6783
rect 3341 6749 3375 6783
rect 3525 6749 3559 6783
rect 3617 6749 3651 6783
rect 3801 6749 3835 6783
rect 4261 6749 4295 6783
rect 4353 6749 4387 6783
rect 4445 6749 4479 6783
rect 4905 6749 4939 6783
rect 5457 6749 5491 6783
rect 6653 6749 6687 6783
rect 7113 6749 7147 6783
rect 7665 6749 7699 6783
rect 8217 6749 8251 6783
rect 10699 6759 10733 6793
rect 10793 6751 10827 6785
rect 12265 6749 12299 6783
rect 14013 6749 14047 6783
rect 15853 6749 15887 6783
rect 16221 6749 16255 6783
rect 16405 6749 16439 6783
rect 3709 6681 3743 6715
rect 7389 6681 7423 6715
rect 7573 6681 7607 6715
rect 10425 6681 10459 6715
rect 10589 6681 10623 6715
rect 857 6613 891 6647
rect 1225 6613 1259 6647
rect 2237 6613 2271 6647
rect 3249 6613 3283 6647
rect 4077 6613 4111 6647
rect 4721 6613 4755 6647
rect 5181 6613 5215 6647
rect 5825 6613 5859 6647
rect 7205 6613 7239 6647
rect 7665 6613 7699 6647
rect 7757 6613 7791 6647
rect 8401 6613 8435 6647
rect 9413 6613 9447 6647
rect 9505 6613 9539 6647
rect 10701 6613 10735 6647
rect 12265 6613 12299 6647
rect 13369 6613 13403 6647
rect 15761 6613 15795 6647
rect 16221 6613 16255 6647
rect 3525 6409 3559 6443
rect 5733 6409 5767 6443
rect 5917 6409 5951 6443
rect 6285 6409 6319 6443
rect 6745 6409 6779 6443
rect 7113 6409 7147 6443
rect 8861 6409 8895 6443
rect 10701 6409 10735 6443
rect 11805 6409 11839 6443
rect 12449 6409 12483 6443
rect 12817 6409 12851 6443
rect 12909 6409 12943 6443
rect 14013 6409 14047 6443
rect 14565 6409 14599 6443
rect 16589 6409 16623 6443
rect 16681 6409 16715 6443
rect 17049 6409 17083 6443
rect 17601 6409 17635 6443
rect 17693 6409 17727 6443
rect 18337 6409 18371 6443
rect 5641 6341 5675 6375
rect 8769 6341 8803 6375
rect 9137 6341 9171 6375
rect 14933 6341 14967 6375
rect 673 6273 707 6307
rect 1041 6273 1075 6307
rect 3157 6273 3191 6307
rect 5549 6273 5583 6307
rect 5825 6273 5859 6307
rect 6377 6273 6411 6307
rect 8677 6273 8711 6307
rect 8953 6273 8987 6307
rect 9045 6273 9079 6307
rect 11161 6273 11195 6307
rect 11897 6273 11931 6307
rect 13921 6273 13955 6307
rect 14105 6273 14139 6307
rect 14381 6273 14415 6307
rect 14657 6273 14691 6307
rect 15025 6273 15059 6307
rect 15577 6273 15611 6307
rect 18245 6273 18279 6307
rect 18521 6273 18555 6307
rect 2697 6205 2731 6239
rect 3065 6205 3099 6239
rect 6561 6205 6595 6239
rect 7205 6205 7239 6239
rect 7297 6205 7331 6239
rect 11069 6205 11103 6239
rect 12081 6205 12115 6239
rect 13001 6205 13035 6239
rect 14197 6205 14231 6239
rect 15669 6205 15703 6239
rect 15761 6205 15795 6239
rect 16405 6205 16439 6239
rect 17877 6205 17911 6239
rect 2467 6137 2501 6171
rect 11345 6137 11379 6171
rect 15209 6137 15243 6171
rect 17233 6137 17267 6171
rect 2881 6069 2915 6103
rect 4169 6069 4203 6103
rect 11437 6069 11471 6103
rect 16129 6069 16163 6103
rect 2316 5865 2350 5899
rect 3801 5865 3835 5899
rect 6561 5865 6595 5899
rect 10793 5865 10827 5899
rect 6009 5797 6043 5831
rect 6883 5797 6917 5831
rect 13001 5797 13035 5831
rect 15485 5797 15519 5831
rect 15577 5797 15611 5831
rect 16313 5797 16347 5831
rect 2053 5729 2087 5763
rect 4261 5729 4295 5763
rect 8861 5729 8895 5763
rect 11253 5729 11287 5763
rect 14749 5729 14783 5763
rect 15209 5729 15243 5763
rect 6653 5661 6687 5695
rect 8309 5661 8343 5695
rect 8677 5661 8711 5695
rect 10609 5661 10643 5695
rect 13829 5661 13863 5695
rect 14473 5661 14507 5695
rect 15117 5661 15151 5695
rect 4537 5593 4571 5627
rect 11529 5593 11563 5627
rect 14565 5593 14599 5627
rect 16504 5729 16538 5763
rect 16405 5661 16439 5695
rect 16129 5593 16163 5627
rect 16773 5593 16807 5627
rect 4169 5525 4203 5559
rect 6285 5525 6319 5559
rect 10977 5525 11011 5559
rect 13645 5525 13679 5559
rect 14105 5525 14139 5559
rect 15577 5525 15611 5559
rect 15761 5525 15795 5559
rect 16405 5525 16439 5559
rect 18245 5525 18279 5559
rect 4077 5321 4111 5355
rect 5549 5321 5583 5355
rect 8677 5321 8711 5355
rect 9413 5321 9447 5355
rect 14657 5321 14691 5355
rect 16313 5321 16347 5355
rect 9689 5253 9723 5287
rect 9873 5253 9907 5287
rect 12725 5253 12759 5287
rect 5641 5185 5675 5219
rect 8585 5185 8619 5219
rect 8769 5185 8803 5219
rect 9045 5185 9079 5219
rect 11805 5185 11839 5219
rect 12909 5185 12943 5219
rect 15761 5185 15795 5219
rect 16221 5185 16255 5219
rect 16681 5185 16715 5219
rect 17049 5185 17083 5219
rect 18245 5185 18279 5219
rect 18521 5185 18555 5219
rect 6009 5117 6043 5151
rect 8953 5117 8987 5151
rect 10057 5117 10091 5151
rect 11529 5117 11563 5151
rect 13185 5117 13219 5151
rect 15853 5117 15887 5151
rect 16129 5117 16163 5151
rect 7389 4981 7423 5015
rect 18337 4981 18371 5015
rect 4905 4777 4939 4811
rect 5917 4777 5951 4811
rect 7941 4777 7975 4811
rect 12743 4777 12777 4811
rect 3893 4709 3927 4743
rect 6469 4709 6503 4743
rect 949 4641 983 4675
rect 1225 4641 1259 4675
rect 2145 4641 2179 4675
rect 4721 4641 4755 4675
rect 6929 4641 6963 4675
rect 7113 4641 7147 4675
rect 9965 4641 9999 4675
rect 11069 4641 11103 4675
rect 14105 4641 14139 4675
rect 1317 4573 1351 4607
rect 4537 4573 4571 4607
rect 4905 4573 4939 4607
rect 4997 4573 5031 4607
rect 6101 4573 6135 4607
rect 13001 4573 13035 4607
rect 13921 4573 13955 4607
rect 17877 4573 17911 4607
rect 18245 4573 18279 4607
rect 2421 4505 2455 4539
rect 5181 4505 5215 4539
rect 6837 4505 6871 4539
rect 13737 4505 13771 4539
rect 14350 4505 14384 4539
rect 4077 4437 4111 4471
rect 4445 4437 4479 4471
rect 11253 4437 11287 4471
rect 15485 4437 15519 4471
rect 16221 4437 16255 4471
rect 16451 4437 16485 4471
rect 2973 4233 3007 4267
rect 5549 4233 5583 4267
rect 7113 4233 7147 4267
rect 10701 4233 10735 4267
rect 18337 4233 18371 4267
rect 949 4165 983 4199
rect 6745 4165 6779 4199
rect 3157 4097 3191 4131
rect 3893 4097 3927 4131
rect 4077 4097 4111 4131
rect 4721 4097 4755 4131
rect 5917 4097 5951 4131
rect 7297 4097 7331 4131
rect 7757 4097 7791 4131
rect 8033 4097 8067 4131
rect 10609 4097 10643 4131
rect 11069 4097 11103 4131
rect 11253 4097 11287 4131
rect 15485 4097 15519 4131
rect 16037 4097 16071 4131
rect 18245 4097 18279 4131
rect 18521 4097 18555 4131
rect 213 4029 247 4063
rect 673 4029 707 4063
rect 2421 4029 2455 4063
rect 4813 4029 4847 4063
rect 6009 4029 6043 4063
rect 6193 4029 6227 4063
rect 6469 4029 6503 4063
rect 6653 4029 6687 4063
rect 7205 4029 7239 4063
rect 8401 4029 8435 4063
rect 10885 4029 10919 4063
rect 11161 4029 11195 4063
rect 12449 4029 12483 4063
rect 12725 4029 12759 4063
rect 14473 4029 14507 4063
rect 5089 3961 5123 3995
rect 15025 3961 15059 3995
rect 2605 3893 2639 3927
rect 4077 3893 4111 3927
rect 7849 3893 7883 3927
rect 9827 3893 9861 3927
rect 10241 3893 10275 3927
rect 12265 3893 12299 3927
rect 15209 3893 15243 3927
rect 15577 3893 15611 3927
rect 15761 3893 15795 3927
rect 4445 3689 4479 3723
rect 6561 3689 6595 3723
rect 8217 3689 8251 3723
rect 10241 3621 10275 3655
rect 12725 3621 12759 3655
rect 13185 3621 13219 3655
rect 13737 3621 13771 3655
rect 213 3553 247 3587
rect 2145 3553 2179 3587
rect 3893 3553 3927 3587
rect 7941 3553 7975 3587
rect 8401 3553 8435 3587
rect 11345 3553 11379 3587
rect 13369 3553 13403 3587
rect 13921 3553 13955 3587
rect 14197 3553 14231 3587
rect 18245 3553 18279 3587
rect 949 3485 983 3519
rect 4077 3485 4111 3519
rect 5273 3485 5307 3519
rect 5457 3485 5491 3519
rect 6469 3485 6503 3519
rect 6653 3485 6687 3519
rect 7537 3485 7571 3519
rect 7655 3485 7689 3519
rect 7757 3495 7791 3529
rect 8493 3485 8527 3519
rect 8861 3485 8895 3519
rect 9965 3485 9999 3519
rect 11601 3485 11635 3519
rect 12909 3485 12943 3519
rect 13001 3485 13035 3519
rect 13277 3485 13311 3519
rect 13461 3485 13495 3519
rect 13645 3485 13679 3519
rect 17877 3485 17911 3519
rect 2421 3417 2455 3451
rect 14464 3417 14498 3451
rect 857 3349 891 3383
rect 4261 3349 4295 3383
rect 5365 3349 5399 3383
rect 9321 3349 9355 3383
rect 10425 3349 10459 3383
rect 13921 3349 13955 3383
rect 15577 3349 15611 3383
rect 15761 3349 15795 3383
rect 16129 3349 16163 3383
rect 3433 3145 3467 3179
rect 6837 3145 6871 3179
rect 13093 3145 13127 3179
rect 15393 3145 15427 3179
rect 16497 3145 16531 3179
rect 4353 3077 4387 3111
rect 10333 3077 10367 3111
rect 15485 3077 15519 3111
rect 15669 3077 15703 3111
rect 673 3009 707 3043
rect 3157 3009 3191 3043
rect 3617 3009 3651 3043
rect 3709 3009 3743 3043
rect 3985 3009 4019 3043
rect 4445 3009 4479 3043
rect 4721 3009 4755 3043
rect 5089 3009 5123 3043
rect 5273 3009 5307 3043
rect 5457 3009 5491 3043
rect 5825 3009 5859 3043
rect 5917 3009 5951 3043
rect 6193 3009 6227 3043
rect 7665 3009 7699 3043
rect 9459 3009 9493 3043
rect 9781 3009 9815 3043
rect 10149 3009 10183 3043
rect 10425 3009 10459 3043
rect 10793 3009 10827 3043
rect 11161 3009 11195 3043
rect 12725 3009 12759 3043
rect 13277 3009 13311 3043
rect 13553 3009 13587 3043
rect 15025 3009 15059 3043
rect 15209 3009 15243 3043
rect 15301 3009 15335 3043
rect 15393 3009 15427 3043
rect 16405 3009 16439 3043
rect 1041 2941 1075 2975
rect 4169 2941 4203 2975
rect 4537 2941 4571 2975
rect 7481 2941 7515 2975
rect 8033 2941 8067 2975
rect 9689 2941 9723 2975
rect 10885 2941 10919 2975
rect 3985 2873 4019 2907
rect 4813 2873 4847 2907
rect 5089 2873 5123 2907
rect 5365 2873 5399 2907
rect 6101 2873 6135 2907
rect 2467 2805 2501 2839
rect 2697 2805 2731 2839
rect 3249 2805 3283 2839
rect 5825 2805 5859 2839
rect 7021 2805 7055 2839
rect 12817 2805 12851 2839
rect 13461 2805 13495 2839
rect 14841 2805 14875 2839
rect 1501 2601 1535 2635
rect 4905 2601 4939 2635
rect 11299 2601 11333 2635
rect 13645 2601 13679 2635
rect 16037 2601 16071 2635
rect 1409 2533 1443 2567
rect 6653 2533 6687 2567
rect 6929 2533 6963 2567
rect 7297 2533 7331 2567
rect 10241 2533 10275 2567
rect 13185 2533 13219 2567
rect 1041 2465 1075 2499
rect 1869 2465 1903 2499
rect 3341 2465 3375 2499
rect 4169 2465 4203 2499
rect 4905 2465 4939 2499
rect 5549 2465 5583 2499
rect 8125 2465 8159 2499
rect 9965 2465 9999 2499
rect 11069 2465 11103 2499
rect 14105 2465 14139 2499
rect 16221 2465 16255 2499
rect 18245 2465 18279 2499
rect 1961 2397 1995 2431
rect 2605 2397 2639 2431
rect 3249 2397 3283 2431
rect 3893 2397 3927 2431
rect 4721 2397 4755 2431
rect 5365 2397 5399 2431
rect 5825 2397 5859 2431
rect 6009 2397 6043 2431
rect 6469 2397 6503 2431
rect 6587 2397 6621 2431
rect 7021 2397 7055 2431
rect 7205 2397 7239 2431
rect 7297 2397 7331 2431
rect 7849 2397 7883 2431
rect 8033 2397 8067 2431
rect 9045 2397 9079 2431
rect 9597 2397 9631 2431
rect 9873 2397 9907 2431
rect 12725 2397 12759 2431
rect 13093 2397 13127 2431
rect 13201 2397 13235 2431
rect 13829 2397 13863 2431
rect 2329 2329 2363 2363
rect 7389 2329 7423 2363
rect 8861 2329 8895 2363
rect 13277 2329 13311 2363
rect 13461 2329 13495 2363
rect 15853 2329 15887 2363
rect 17969 2329 18003 2363
rect 1685 2261 1719 2295
rect 4997 2261 5031 2295
rect 5457 2261 5491 2295
rect 5825 2261 5859 2295
rect 10609 2261 10643 2295
rect 673 2057 707 2091
rect 2605 2057 2639 2091
rect 2973 2057 3007 2091
rect 7665 2057 7699 2091
rect 12817 2057 12851 2091
rect 13553 2057 13587 2091
rect 15669 2057 15703 2091
rect 17233 2057 17267 2091
rect 17693 2057 17727 2091
rect 18153 2057 18187 2091
rect 7757 1989 7791 2023
rect 8585 1989 8619 2023
rect 12265 1989 12299 2023
rect 14565 1989 14599 2023
rect 15761 1989 15795 2023
rect 17601 1989 17635 2023
rect 2421 1921 2455 1955
rect 2513 1921 2547 1955
rect 2697 1921 2731 1955
rect 3065 1921 3099 1955
rect 3433 1921 3467 1955
rect 3525 1921 3559 1955
rect 3617 1921 3651 1955
rect 4169 1921 4203 1955
rect 4261 1921 4295 1955
rect 5273 1921 5307 1955
rect 5457 1921 5491 1955
rect 5549 1921 5583 1955
rect 7665 1921 7699 1955
rect 7941 1921 7975 1955
rect 8217 1921 8251 1955
rect 8401 1921 8435 1955
rect 8769 1921 8803 1955
rect 9873 1921 9907 1955
rect 10333 1921 10367 1955
rect 10793 1921 10827 1955
rect 2145 1853 2179 1887
rect 4077 1853 4111 1887
rect 5825 1853 5859 1887
rect 10241 1853 10275 1887
rect 10977 1853 11011 1887
rect 3249 1785 3283 1819
rect 13001 1921 13035 1955
rect 13093 1921 13127 1955
rect 13221 1921 13255 1955
rect 13645 1921 13679 1955
rect 13829 1921 13863 1955
rect 14289 1921 14323 1955
rect 14381 1921 14415 1955
rect 16497 1921 16531 1955
rect 18061 1921 18095 1955
rect 18521 1921 18555 1955
rect 13369 1853 13403 1887
rect 15853 1853 15887 1887
rect 16589 1853 16623 1887
rect 16681 1853 16715 1887
rect 17877 1853 17911 1887
rect 16129 1785 16163 1819
rect 3893 1717 3927 1751
rect 4353 1717 4387 1751
rect 5365 1717 5399 1751
rect 8861 1717 8895 1751
rect 9413 1717 9447 1751
rect 11253 1717 11287 1751
rect 12265 1717 12299 1751
rect 14473 1717 14507 1751
rect 15301 1717 15335 1751
rect 18337 1717 18371 1751
rect 5365 1513 5399 1547
rect 18061 1513 18095 1547
rect 18521 1513 18555 1547
rect 4537 1445 4571 1479
rect 11253 1445 11287 1479
rect 2145 1377 2179 1411
rect 2421 1377 2455 1411
rect 4445 1377 4479 1411
rect 5825 1377 5859 1411
rect 6009 1377 6043 1411
rect 7757 1377 7791 1411
rect 8493 1377 8527 1411
rect 9781 1377 9815 1411
rect 9873 1377 9907 1411
rect 12265 1377 12299 1411
rect 13093 1377 13127 1411
rect 13277 1377 13311 1411
rect 14013 1377 14047 1411
rect 16589 1377 16623 1411
rect 4629 1309 4663 1343
rect 4721 1309 4755 1343
rect 4997 1309 5031 1343
rect 6469 1309 6503 1343
rect 6653 1309 6687 1343
rect 6929 1309 6963 1343
rect 8401 1309 8435 1343
rect 10609 1309 10643 1343
rect 10701 1309 10735 1343
rect 11069 1309 11103 1343
rect 11253 1309 11287 1343
rect 11529 1309 11563 1343
rect 12081 1309 12115 1343
rect 13645 1309 13679 1343
rect 14381 1309 14415 1343
rect 16313 1309 16347 1343
rect 4905 1241 4939 1275
rect 5733 1241 5767 1275
rect 7481 1241 7515 1275
rect 8309 1241 8343 1275
rect 11345 1241 11379 1275
rect 13001 1241 13035 1275
rect 13737 1241 13771 1275
rect 13921 1241 13955 1275
rect 15807 1241 15841 1275
rect 3893 1173 3927 1207
rect 4169 1173 4203 1207
rect 6469 1173 6503 1207
rect 6837 1173 6871 1207
rect 7113 1173 7147 1207
rect 7573 1173 7607 1207
rect 7941 1173 7975 1207
rect 9321 1173 9355 1207
rect 9689 1173 9723 1207
rect 10425 1173 10459 1207
rect 11621 1173 11655 1207
rect 11989 1173 12023 1207
rect 12633 1173 12667 1207
rect 13645 1173 13679 1207
rect 16129 1173 16163 1207
rect 2927 969 2961 1003
rect 7297 969 7331 1003
rect 8677 969 8711 1003
rect 9413 969 9447 1003
rect 9505 969 9539 1003
rect 10333 969 10367 1003
rect 12173 969 12207 1003
rect 12633 969 12667 1003
rect 13369 969 13403 1003
rect 13645 969 13679 1003
rect 14657 969 14691 1003
rect 15117 969 15151 1003
rect 17233 969 17267 1003
rect 18245 969 18279 1003
rect 10701 901 10735 935
rect 13921 901 13955 935
rect 14841 901 14875 935
rect 15025 901 15059 935
rect 4721 833 4755 867
rect 5089 833 5123 867
rect 5273 833 5307 867
rect 5549 833 5583 867
rect 7849 833 7883 867
rect 8033 833 8067 867
rect 8125 833 8159 867
rect 8401 833 8435 867
rect 8953 833 8987 867
rect 12541 833 12575 867
rect 13277 833 13311 867
rect 13737 833 13771 867
rect 15101 823 15135 857
rect 17601 833 17635 867
rect 18061 833 18095 867
rect 2697 765 2731 799
rect 4353 765 4387 799
rect 4813 765 4847 799
rect 5825 765 5859 799
rect 9597 765 9631 799
rect 10425 765 10459 799
rect 14197 765 14231 799
rect 14289 765 14323 799
rect 15209 765 15243 799
rect 15485 765 15519 799
rect 17693 765 17727 799
rect 17877 765 17911 799
rect 4905 697 4939 731
rect 16957 697 16991 731
rect 4997 629 5031 663
rect 5365 629 5399 663
rect 8033 629 8067 663
rect 9045 629 9079 663
rect 14013 629 14047 663
rect 4997 425 5031 459
rect 5825 425 5859 459
rect 5917 425 5951 459
rect 6561 425 6595 459
rect 8401 425 8435 459
rect 13001 425 13035 459
rect 15025 425 15059 459
rect 15761 425 15795 459
rect 17693 425 17727 459
rect 18061 425 18095 459
rect 18521 425 18555 459
rect 9413 357 9447 391
rect 5733 289 5767 323
rect 8125 289 8159 323
rect 8953 289 8987 323
rect 12725 289 12759 323
rect 13277 289 13311 323
rect 15117 289 15151 323
rect 15485 289 15519 323
rect 17325 289 17359 323
rect 4905 221 4939 255
rect 5089 221 5123 255
rect 5457 221 5491 255
rect 6009 221 6043 255
rect 6745 221 6779 255
rect 8033 221 8067 255
rect 9045 221 9079 255
rect 12633 221 12667 255
rect 13185 221 13219 255
rect 13369 221 13403 255
rect 15577 221 15611 255
rect 17417 221 17451 255
rect 18245 221 18279 255
rect 6469 153 6503 187
rect 6653 153 6687 187
<< metal1 >>
rect 368 10906 18860 10928
rect 368 10854 5028 10906
rect 5080 10854 5092 10906
rect 5144 10854 5156 10906
rect 5208 10854 5220 10906
rect 5272 10854 5284 10906
rect 5336 10854 8128 10906
rect 8180 10854 8192 10906
rect 8244 10854 8256 10906
rect 8308 10854 8320 10906
rect 8372 10854 8384 10906
rect 8436 10854 11228 10906
rect 11280 10854 11292 10906
rect 11344 10854 11356 10906
rect 11408 10854 11420 10906
rect 11472 10854 11484 10906
rect 11536 10854 14328 10906
rect 14380 10854 14392 10906
rect 14444 10854 14456 10906
rect 14508 10854 14520 10906
rect 14572 10854 14584 10906
rect 14636 10854 17428 10906
rect 17480 10854 17492 10906
rect 17544 10854 17556 10906
rect 17608 10854 17620 10906
rect 17672 10854 17684 10906
rect 17736 10854 18860 10906
rect 368 10832 18860 10854
rect 6822 10792 6828 10804
rect 6783 10764 6828 10792
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 7392 10764 9904 10792
rect 7392 10724 7420 10764
rect 6656 10696 7420 10724
rect 7469 10727 7527 10733
rect 658 10616 664 10668
rect 716 10656 722 10668
rect 2317 10659 2375 10665
rect 2317 10656 2329 10659
rect 716 10628 2329 10656
rect 716 10616 722 10628
rect 2317 10625 2329 10628
rect 2363 10625 2375 10659
rect 2317 10619 2375 10625
rect 2406 10616 2412 10668
rect 2464 10656 2470 10668
rect 2593 10659 2651 10665
rect 2593 10656 2605 10659
rect 2464 10628 2605 10656
rect 2464 10616 2470 10628
rect 2593 10625 2605 10628
rect 2639 10625 2651 10659
rect 2593 10619 2651 10625
rect 3050 10616 3056 10668
rect 3108 10656 3114 10668
rect 3145 10659 3203 10665
rect 3145 10656 3157 10659
rect 3108 10628 3157 10656
rect 3108 10616 3114 10628
rect 3145 10625 3157 10628
rect 3191 10625 3203 10659
rect 5258 10656 5264 10668
rect 5219 10628 5264 10656
rect 3145 10619 3203 10625
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 5442 10656 5448 10668
rect 5403 10628 5448 10656
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 6656 10665 6684 10696
rect 7469 10693 7481 10727
rect 7515 10724 7527 10727
rect 8297 10727 8355 10733
rect 8297 10724 8309 10727
rect 7515 10696 8309 10724
rect 7515 10693 7527 10696
rect 7469 10687 7527 10693
rect 8297 10693 8309 10696
rect 8343 10693 8355 10727
rect 9876 10724 9904 10764
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10045 10795 10103 10801
rect 10045 10792 10057 10795
rect 10008 10764 10057 10792
rect 10008 10752 10014 10764
rect 10045 10761 10057 10764
rect 10091 10761 10103 10795
rect 10045 10755 10103 10761
rect 12894 10752 12900 10804
rect 12952 10792 12958 10804
rect 13725 10795 13783 10801
rect 13725 10792 13737 10795
rect 12952 10764 13737 10792
rect 12952 10752 12958 10764
rect 13725 10761 13737 10764
rect 13771 10761 13783 10795
rect 18233 10795 18291 10801
rect 18233 10792 18245 10795
rect 13725 10755 13783 10761
rect 17604 10764 18245 10792
rect 9876 10696 12434 10724
rect 8297 10687 8355 10693
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10656 7343 10659
rect 8754 10656 8760 10668
rect 7331 10628 8760 10656
rect 7331 10625 7343 10628
rect 7285 10619 7343 10625
rect 2869 10591 2927 10597
rect 2869 10557 2881 10591
rect 2915 10588 2927 10591
rect 3234 10588 3240 10600
rect 2915 10560 3240 10588
rect 2915 10557 2927 10560
rect 2869 10551 2927 10557
rect 3234 10548 3240 10560
rect 3292 10548 3298 10600
rect 6932 10588 6960 10619
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10625 8907 10659
rect 8849 10619 8907 10625
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10656 10287 10659
rect 11146 10656 11152 10668
rect 10275 10628 11152 10656
rect 10275 10625 10287 10628
rect 10229 10619 10287 10625
rect 8297 10591 8355 10597
rect 6932 10560 7880 10588
rect 2682 10480 2688 10532
rect 2740 10520 2746 10532
rect 7852 10529 7880 10560
rect 8297 10557 8309 10591
rect 8343 10557 8355 10591
rect 8297 10551 8355 10557
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10588 8447 10591
rect 8570 10588 8576 10600
rect 8435 10560 8576 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 3053 10523 3111 10529
rect 3053 10520 3065 10523
rect 2740 10492 3065 10520
rect 2740 10480 2746 10492
rect 3053 10489 3065 10492
rect 3099 10489 3111 10523
rect 3053 10483 3111 10489
rect 7837 10523 7895 10529
rect 7837 10489 7849 10523
rect 7883 10489 7895 10523
rect 8312 10520 8340 10551
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 8478 10520 8484 10532
rect 8312 10492 8484 10520
rect 7837 10483 7895 10489
rect 8478 10480 8484 10492
rect 8536 10520 8542 10532
rect 8864 10520 8892 10619
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 12406 10656 12434 10696
rect 12526 10684 12532 10736
rect 12584 10724 12590 10736
rect 12805 10727 12863 10733
rect 12805 10724 12817 10727
rect 12584 10696 12817 10724
rect 12584 10684 12590 10696
rect 12805 10693 12817 10696
rect 12851 10693 12863 10727
rect 12805 10687 12863 10693
rect 13170 10656 13176 10668
rect 12406 10628 13176 10656
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 17604 10665 17632 10764
rect 18233 10761 18245 10764
rect 18279 10792 18291 10795
rect 18782 10792 18788 10804
rect 18279 10764 18788 10792
rect 18279 10761 18291 10764
rect 18233 10755 18291 10761
rect 18782 10752 18788 10764
rect 18840 10752 18846 10804
rect 17957 10727 18015 10733
rect 17957 10724 17969 10727
rect 17696 10696 17969 10724
rect 13909 10659 13967 10665
rect 13909 10625 13921 10659
rect 13955 10625 13967 10659
rect 13909 10619 13967 10625
rect 17589 10659 17647 10665
rect 17589 10625 17601 10659
rect 17635 10625 17647 10659
rect 17589 10619 17647 10625
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12529 10591 12587 10597
rect 12529 10588 12541 10591
rect 12492 10560 12541 10588
rect 12492 10548 12498 10560
rect 12529 10557 12541 10560
rect 12575 10557 12587 10591
rect 12529 10551 12587 10557
rect 12713 10591 12771 10597
rect 12713 10557 12725 10591
rect 12759 10588 12771 10591
rect 13262 10588 13268 10600
rect 12759 10560 13268 10588
rect 12759 10557 12771 10560
rect 12713 10551 12771 10557
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 13924 10588 13952 10619
rect 17696 10588 17724 10696
rect 17957 10693 17969 10696
rect 18003 10693 18015 10727
rect 17957 10687 18015 10693
rect 17865 10659 17923 10665
rect 17865 10656 17877 10659
rect 13924 10560 17724 10588
rect 17788 10628 17877 10656
rect 17788 10529 17816 10628
rect 17865 10625 17877 10628
rect 17911 10625 17923 10659
rect 18046 10656 18052 10668
rect 18007 10628 18052 10656
rect 17865 10619 17923 10625
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 8536 10492 8892 10520
rect 17773 10523 17831 10529
rect 8536 10480 8542 10492
rect 17773 10489 17785 10523
rect 17819 10489 17831 10523
rect 17773 10483 17831 10489
rect 2038 10412 2044 10464
rect 2096 10452 2102 10464
rect 2225 10455 2283 10461
rect 2225 10452 2237 10455
rect 2096 10424 2237 10452
rect 2096 10412 2102 10424
rect 2225 10421 2237 10424
rect 2271 10421 2283 10455
rect 2225 10415 2283 10421
rect 2501 10455 2559 10461
rect 2501 10421 2513 10455
rect 2547 10452 2559 10455
rect 2590 10452 2596 10464
rect 2547 10424 2596 10452
rect 2547 10421 2559 10424
rect 2501 10415 2559 10421
rect 2590 10412 2596 10424
rect 2648 10412 2654 10464
rect 2958 10452 2964 10464
rect 2919 10424 2964 10452
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 4430 10412 4436 10464
rect 4488 10452 4494 10464
rect 5261 10455 5319 10461
rect 5261 10452 5273 10455
rect 4488 10424 5273 10452
rect 4488 10412 4494 10424
rect 5261 10421 5273 10424
rect 5307 10421 5319 10455
rect 5261 10415 5319 10421
rect 7101 10455 7159 10461
rect 7101 10421 7113 10455
rect 7147 10452 7159 10455
rect 7282 10452 7288 10464
rect 7147 10424 7288 10452
rect 7147 10421 7159 10424
rect 7101 10415 7159 10421
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 8570 10452 8576 10464
rect 8531 10424 8576 10452
rect 8570 10412 8576 10424
rect 8628 10412 8634 10464
rect 9122 10412 9128 10464
rect 9180 10452 9186 10464
rect 9493 10455 9551 10461
rect 9493 10452 9505 10455
rect 9180 10424 9505 10452
rect 9180 10412 9186 10424
rect 9493 10421 9505 10424
rect 9539 10421 9551 10455
rect 9493 10415 9551 10421
rect 11333 10455 11391 10461
rect 11333 10421 11345 10455
rect 11379 10452 11391 10455
rect 11974 10452 11980 10464
rect 11379 10424 11980 10452
rect 11379 10421 11391 10424
rect 11333 10415 11391 10421
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 13170 10452 13176 10464
rect 13131 10424 13176 10452
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 13998 10452 14004 10464
rect 13959 10424 14004 10452
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 14921 10455 14979 10461
rect 14921 10421 14933 10455
rect 14967 10452 14979 10455
rect 15286 10452 15292 10464
rect 14967 10424 15292 10452
rect 14967 10421 14979 10424
rect 14921 10415 14979 10421
rect 15286 10412 15292 10424
rect 15344 10412 15350 10464
rect 368 10362 18860 10384
rect 368 10310 3478 10362
rect 3530 10310 3542 10362
rect 3594 10310 3606 10362
rect 3658 10310 3670 10362
rect 3722 10310 3734 10362
rect 3786 10310 6578 10362
rect 6630 10310 6642 10362
rect 6694 10310 6706 10362
rect 6758 10310 6770 10362
rect 6822 10310 6834 10362
rect 6886 10310 9678 10362
rect 9730 10310 9742 10362
rect 9794 10310 9806 10362
rect 9858 10310 9870 10362
rect 9922 10310 9934 10362
rect 9986 10310 12778 10362
rect 12830 10310 12842 10362
rect 12894 10310 12906 10362
rect 12958 10310 12970 10362
rect 13022 10310 13034 10362
rect 13086 10310 15878 10362
rect 15930 10310 15942 10362
rect 15994 10310 16006 10362
rect 16058 10310 16070 10362
rect 16122 10310 16134 10362
rect 16186 10310 18860 10362
rect 368 10288 18860 10310
rect 1857 10251 1915 10257
rect 1857 10217 1869 10251
rect 1903 10248 1915 10251
rect 2682 10248 2688 10260
rect 1903 10220 2688 10248
rect 1903 10217 1915 10220
rect 1857 10211 1915 10217
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 4246 10208 4252 10260
rect 4304 10248 4310 10260
rect 4304 10220 8340 10248
rect 4304 10208 4310 10220
rect 5258 10180 5264 10192
rect 3160 10152 5264 10180
rect 3160 10124 3188 10152
rect 5258 10140 5264 10152
rect 5316 10180 5322 10192
rect 8312 10180 8340 10220
rect 8478 10208 8484 10260
rect 8536 10248 8542 10260
rect 8573 10251 8631 10257
rect 8573 10248 8585 10251
rect 8536 10220 8585 10248
rect 8536 10208 8542 10220
rect 8573 10217 8585 10220
rect 8619 10217 8631 10251
rect 8573 10211 8631 10217
rect 8754 10208 8760 10260
rect 8812 10248 8818 10260
rect 10597 10251 10655 10257
rect 10597 10248 10609 10251
rect 8812 10220 10609 10248
rect 8812 10208 8818 10220
rect 10597 10217 10609 10220
rect 10643 10248 10655 10251
rect 12618 10248 12624 10260
rect 10643 10220 12624 10248
rect 10643 10217 10655 10220
rect 10597 10211 10655 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 18046 10257 18052 10260
rect 18003 10251 18052 10257
rect 18003 10217 18015 10251
rect 18049 10217 18052 10251
rect 18003 10211 18052 10217
rect 18046 10208 18052 10211
rect 18104 10208 18110 10260
rect 9125 10183 9183 10189
rect 9125 10180 9137 10183
rect 5316 10152 5672 10180
rect 8312 10152 9137 10180
rect 5316 10140 5322 10152
rect 1670 10112 1676 10124
rect 1631 10084 1676 10112
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 2038 10112 2044 10124
rect 1999 10084 2044 10112
rect 2038 10072 2044 10084
rect 2096 10072 2102 10124
rect 2409 10115 2467 10121
rect 2409 10081 2421 10115
rect 2455 10112 2467 10115
rect 2958 10112 2964 10124
rect 2455 10084 2964 10112
rect 2455 10081 2467 10084
rect 2409 10075 2467 10081
rect 2958 10072 2964 10084
rect 3016 10072 3022 10124
rect 3142 10072 3148 10124
rect 3200 10072 3206 10124
rect 4430 10112 4436 10124
rect 4391 10084 4436 10112
rect 4430 10072 4436 10084
rect 4488 10072 4494 10124
rect 4709 10115 4767 10121
rect 4709 10081 4721 10115
rect 4755 10112 4767 10115
rect 5534 10112 5540 10124
rect 4755 10084 5540 10112
rect 4755 10081 4767 10084
rect 4709 10075 4767 10081
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 5644 10112 5672 10152
rect 9125 10149 9137 10152
rect 9171 10149 9183 10183
rect 9125 10143 9183 10149
rect 5813 10115 5871 10121
rect 5813 10112 5825 10115
rect 5644 10084 5825 10112
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10044 2007 10047
rect 2498 10044 2504 10056
rect 1995 10016 2504 10044
rect 1995 10013 2007 10016
rect 1949 10007 2007 10013
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 5644 10053 5672 10084
rect 5813 10081 5825 10084
rect 5859 10081 5871 10115
rect 5813 10075 5871 10081
rect 4341 10047 4399 10053
rect 4341 10044 4353 10047
rect 3712 10016 4353 10044
rect 2774 9936 2780 9988
rect 2832 9936 2838 9988
rect 934 9868 940 9920
rect 992 9908 998 9920
rect 1673 9911 1731 9917
rect 1673 9908 1685 9911
rect 992 9880 1685 9908
rect 992 9868 998 9880
rect 1673 9877 1685 9880
rect 1719 9877 1731 9911
rect 1673 9871 1731 9877
rect 2406 9868 2412 9920
rect 2464 9908 2470 9920
rect 3712 9908 3740 10016
rect 4341 10013 4353 10016
rect 4387 10044 4399 10047
rect 4801 10047 4859 10053
rect 4801 10044 4813 10047
rect 4387 10016 4813 10044
rect 4387 10013 4399 10016
rect 4341 10007 4399 10013
rect 4801 10013 4813 10016
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10013 5135 10047
rect 5077 10007 5135 10013
rect 5629 10047 5687 10053
rect 5629 10013 5641 10047
rect 5675 10013 5687 10047
rect 5629 10007 5687 10013
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 7190 10044 7196 10056
rect 7151 10016 7196 10044
rect 5905 10007 5963 10013
rect 5092 9976 5120 10007
rect 5442 9976 5448 9988
rect 4816 9948 5448 9976
rect 2464 9880 3740 9908
rect 2464 9868 2470 9880
rect 3786 9868 3792 9920
rect 3844 9917 3850 9920
rect 3844 9911 3893 9917
rect 3844 9877 3847 9911
rect 3881 9908 3893 9911
rect 4816 9908 4844 9948
rect 5442 9936 5448 9948
rect 5500 9976 5506 9988
rect 5920 9976 5948 10007
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 7282 10004 7288 10056
rect 7340 10044 7346 10056
rect 7449 10047 7507 10053
rect 7449 10044 7461 10047
rect 7340 10016 7461 10044
rect 7340 10004 7346 10016
rect 7449 10013 7461 10016
rect 7495 10013 7507 10047
rect 9140 10044 9168 10143
rect 11974 10072 11980 10124
rect 12032 10112 12038 10124
rect 12032 10084 13124 10112
rect 12032 10072 12038 10084
rect 9309 10047 9367 10053
rect 9309 10044 9321 10047
rect 9140 10016 9321 10044
rect 7449 10007 7507 10013
rect 9309 10013 9321 10016
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11241 10047 11299 10053
rect 11241 10044 11253 10047
rect 11112 10016 11253 10044
rect 11112 10004 11118 10016
rect 11241 10013 11253 10016
rect 11287 10013 11299 10047
rect 13096 10044 13124 10084
rect 13170 10072 13176 10124
rect 13228 10112 13234 10124
rect 14001 10115 14059 10121
rect 14001 10112 14013 10115
rect 13228 10084 14013 10112
rect 13228 10072 13234 10084
rect 14001 10081 14013 10084
rect 14047 10112 14059 10115
rect 16209 10115 16267 10121
rect 16209 10112 16221 10115
rect 14047 10084 16221 10112
rect 14047 10081 14059 10084
rect 14001 10075 14059 10081
rect 16209 10081 16221 10084
rect 16255 10081 16267 10115
rect 16209 10075 16267 10081
rect 13096 10016 13216 10044
rect 11241 10007 11299 10013
rect 5500 9948 5948 9976
rect 11517 9979 11575 9985
rect 5500 9936 5506 9948
rect 11517 9945 11529 9979
rect 11563 9976 11575 9979
rect 11606 9976 11612 9988
rect 11563 9948 11612 9976
rect 11563 9945 11575 9948
rect 11517 9939 11575 9945
rect 11606 9936 11612 9948
rect 11664 9936 11670 9988
rect 11974 9936 11980 9988
rect 12032 9936 12038 9988
rect 5350 9908 5356 9920
rect 3881 9880 4844 9908
rect 5311 9880 5356 9908
rect 3881 9877 3893 9880
rect 3844 9871 3893 9877
rect 3844 9868 3850 9871
rect 5350 9868 5356 9880
rect 5408 9868 5414 9920
rect 6270 9908 6276 9920
rect 6231 9880 6276 9908
rect 6270 9868 6276 9880
rect 6328 9868 6334 9920
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 12802 9908 12808 9920
rect 12492 9880 12808 9908
rect 12492 9868 12498 9880
rect 12802 9868 12808 9880
rect 12860 9908 12866 9920
rect 13188 9917 13216 10016
rect 14090 10004 14096 10056
rect 14148 10044 14154 10056
rect 14369 10047 14427 10053
rect 14369 10044 14381 10047
rect 14148 10016 14381 10044
rect 14148 10004 14154 10016
rect 14369 10013 14381 10016
rect 14415 10013 14427 10047
rect 14369 10007 14427 10013
rect 15795 10047 15853 10053
rect 15795 10013 15807 10047
rect 15841 10044 15853 10047
rect 16577 10047 16635 10053
rect 16577 10044 16589 10047
rect 15841 10016 16589 10044
rect 15841 10013 15853 10016
rect 15795 10007 15853 10013
rect 16577 10013 16589 10016
rect 16623 10013 16635 10047
rect 16577 10007 16635 10013
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 12860 9880 13001 9908
rect 12860 9868 12866 9880
rect 12989 9877 13001 9880
rect 13035 9877 13047 9911
rect 12989 9871 13047 9877
rect 13173 9911 13231 9917
rect 13173 9877 13185 9911
rect 13219 9908 13231 9911
rect 13909 9911 13967 9917
rect 13909 9908 13921 9911
rect 13219 9880 13921 9908
rect 13219 9877 13231 9880
rect 13173 9871 13231 9877
rect 13909 9877 13921 9880
rect 13955 9908 13967 9911
rect 15212 9908 15240 9962
rect 15286 9908 15292 9920
rect 13955 9880 15292 9908
rect 13955 9877 13967 9880
rect 13909 9871 13967 9877
rect 15286 9868 15292 9880
rect 15344 9908 15350 9920
rect 16025 9911 16083 9917
rect 16025 9908 16037 9911
rect 15344 9880 16037 9908
rect 15344 9868 15350 9880
rect 16025 9877 16037 9880
rect 16071 9908 16083 9911
rect 16960 9908 16988 9962
rect 16071 9880 16988 9908
rect 16071 9877 16083 9880
rect 16025 9871 16083 9877
rect 368 9818 18860 9840
rect 368 9766 5028 9818
rect 5080 9766 5092 9818
rect 5144 9766 5156 9818
rect 5208 9766 5220 9818
rect 5272 9766 5284 9818
rect 5336 9766 8128 9818
rect 8180 9766 8192 9818
rect 8244 9766 8256 9818
rect 8308 9766 8320 9818
rect 8372 9766 8384 9818
rect 8436 9766 11228 9818
rect 11280 9766 11292 9818
rect 11344 9766 11356 9818
rect 11408 9766 11420 9818
rect 11472 9766 11484 9818
rect 11536 9766 14328 9818
rect 14380 9766 14392 9818
rect 14444 9766 14456 9818
rect 14508 9766 14520 9818
rect 14572 9766 14584 9818
rect 14636 9766 17428 9818
rect 17480 9766 17492 9818
rect 17544 9766 17556 9818
rect 17608 9766 17620 9818
rect 17672 9766 17684 9818
rect 17736 9766 18860 9818
rect 368 9744 18860 9766
rect 1670 9664 1676 9716
rect 1728 9704 1734 9716
rect 2501 9707 2559 9713
rect 2501 9704 2513 9707
rect 1728 9676 2513 9704
rect 1728 9664 1734 9676
rect 2501 9673 2513 9676
rect 2547 9673 2559 9707
rect 2501 9667 2559 9673
rect 3053 9707 3111 9713
rect 3053 9673 3065 9707
rect 3099 9673 3111 9707
rect 3234 9704 3240 9716
rect 3195 9676 3240 9704
rect 3053 9667 3111 9673
rect 934 9636 940 9648
rect 895 9608 940 9636
rect 934 9596 940 9608
rect 992 9596 998 9648
rect 2590 9596 2596 9648
rect 2648 9636 2654 9648
rect 2958 9636 2964 9648
rect 2648 9608 2820 9636
rect 2919 9608 2964 9636
rect 2648 9596 2654 9608
rect 658 9568 664 9580
rect 619 9540 664 9568
rect 658 9528 664 9540
rect 716 9528 722 9580
rect 2498 9568 2504 9580
rect 2056 9500 2084 9554
rect 2459 9540 2504 9568
rect 2498 9528 2504 9540
rect 2556 9528 2562 9580
rect 2685 9571 2743 9577
rect 2685 9537 2697 9571
rect 2731 9537 2743 9571
rect 2792 9568 2820 9608
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 3068 9636 3096 9667
rect 3234 9664 3240 9676
rect 3292 9664 3298 9716
rect 6270 9664 6276 9716
rect 6328 9704 6334 9716
rect 6733 9707 6791 9713
rect 6733 9704 6745 9707
rect 6328 9676 6745 9704
rect 6328 9664 6334 9676
rect 6733 9673 6745 9676
rect 6779 9673 6791 9707
rect 6733 9667 6791 9673
rect 11146 9664 11152 9716
rect 11204 9704 11210 9716
rect 11517 9707 11575 9713
rect 11517 9704 11529 9707
rect 11204 9676 11529 9704
rect 11204 9664 11210 9676
rect 11517 9673 11529 9676
rect 11563 9673 11575 9707
rect 11517 9667 11575 9673
rect 14090 9664 14096 9716
rect 14148 9704 14154 9716
rect 14599 9707 14657 9713
rect 14599 9704 14611 9707
rect 14148 9676 14611 9704
rect 14148 9664 14154 9676
rect 14599 9673 14611 9676
rect 14645 9673 14657 9707
rect 14599 9667 14657 9673
rect 5258 9636 5264 9648
rect 3068 9608 5264 9636
rect 5258 9596 5264 9608
rect 5316 9596 5322 9648
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 5629 9639 5687 9645
rect 5629 9636 5641 9639
rect 5592 9608 5641 9636
rect 5592 9596 5598 9608
rect 5629 9605 5641 9608
rect 5675 9605 5687 9639
rect 5629 9599 5687 9605
rect 10873 9639 10931 9645
rect 10873 9605 10885 9639
rect 10919 9636 10931 9639
rect 12437 9639 12495 9645
rect 12437 9636 12449 9639
rect 10919 9608 12449 9636
rect 10919 9605 10931 9608
rect 10873 9599 10931 9605
rect 12437 9605 12449 9608
rect 12483 9605 12495 9639
rect 12618 9636 12624 9648
rect 12579 9608 12624 9636
rect 12437 9599 12495 9605
rect 12618 9596 12624 9608
rect 12676 9596 12682 9648
rect 14182 9596 14188 9648
rect 14240 9596 14246 9648
rect 15562 9596 15568 9648
rect 15620 9596 15626 9648
rect 2869 9571 2927 9577
rect 2869 9568 2881 9571
rect 2792 9540 2881 9568
rect 2685 9531 2743 9537
rect 2869 9537 2881 9540
rect 2915 9537 2927 9571
rect 3142 9568 3148 9580
rect 3103 9540 3148 9568
rect 2869 9531 2927 9537
rect 2406 9500 2412 9512
rect 2056 9472 2268 9500
rect 2367 9472 2412 9500
rect 2240 9364 2268 9472
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 2700 9500 2728 9531
rect 3142 9528 3148 9540
rect 3200 9528 3206 9580
rect 3234 9528 3240 9580
rect 3292 9568 3298 9580
rect 3421 9571 3479 9577
rect 3292 9540 3337 9568
rect 3292 9528 3298 9540
rect 3421 9537 3433 9571
rect 3467 9537 3479 9571
rect 3786 9568 3792 9580
rect 3747 9540 3792 9568
rect 3421 9531 3479 9537
rect 3436 9500 3464 9531
rect 3786 9528 3792 9540
rect 3844 9528 3850 9580
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9537 4767 9571
rect 4709 9531 4767 9537
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9568 4859 9571
rect 5721 9571 5779 9577
rect 5721 9568 5733 9571
rect 4847 9540 5733 9568
rect 4847 9537 4859 9540
rect 4801 9531 4859 9537
rect 5721 9537 5733 9540
rect 5767 9568 5779 9571
rect 5994 9568 6000 9580
rect 5767 9540 6000 9568
rect 5767 9537 5779 9540
rect 5721 9531 5779 9537
rect 4614 9500 4620 9512
rect 2700 9472 3372 9500
rect 3436 9472 4620 9500
rect 2498 9392 2504 9444
rect 2556 9432 2562 9444
rect 2682 9432 2688 9444
rect 2556 9404 2688 9432
rect 2556 9392 2562 9404
rect 2682 9392 2688 9404
rect 2740 9432 2746 9444
rect 3234 9432 3240 9444
rect 2740 9404 3240 9432
rect 2740 9392 2746 9404
rect 3234 9392 3240 9404
rect 3292 9392 3298 9444
rect 3344 9432 3372 9472
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 4341 9435 4399 9441
rect 4341 9432 4353 9435
rect 3344 9404 4353 9432
rect 4341 9401 4353 9404
rect 4387 9401 4399 9435
rect 4724 9432 4752 9531
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 6362 9528 6368 9580
rect 6420 9568 6426 9580
rect 8754 9577 8760 9580
rect 6641 9571 6699 9577
rect 6641 9568 6653 9571
rect 6420 9540 6653 9568
rect 6420 9528 6426 9540
rect 6641 9537 6653 9540
rect 6687 9537 6699 9571
rect 6641 9531 6699 9537
rect 8748 9531 8760 9577
rect 8812 9568 8818 9580
rect 11606 9568 11612 9580
rect 8812 9540 8848 9568
rect 10612 9540 11612 9568
rect 8754 9528 8760 9531
rect 8812 9528 8818 9540
rect 4985 9503 5043 9509
rect 4985 9469 4997 9503
rect 5031 9500 5043 9503
rect 5813 9503 5871 9509
rect 5031 9472 5396 9500
rect 5031 9469 5043 9472
rect 4985 9463 5043 9469
rect 5261 9435 5319 9441
rect 5261 9432 5273 9435
rect 4724 9404 5273 9432
rect 4341 9395 4399 9401
rect 5261 9401 5273 9404
rect 5307 9401 5319 9435
rect 5261 9395 5319 9401
rect 2866 9364 2872 9376
rect 2240 9336 2872 9364
rect 2866 9324 2872 9336
rect 2924 9324 2930 9376
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 3697 9367 3755 9373
rect 3697 9364 3709 9367
rect 3108 9336 3709 9364
rect 3108 9324 3114 9336
rect 3697 9333 3709 9336
rect 3743 9333 3755 9367
rect 4062 9364 4068 9376
rect 4023 9336 4068 9364
rect 3697 9327 3755 9333
rect 4062 9324 4068 9336
rect 4120 9364 4126 9376
rect 4157 9367 4215 9373
rect 4157 9364 4169 9367
rect 4120 9336 4169 9364
rect 4120 9324 4126 9336
rect 4157 9333 4169 9336
rect 4203 9333 4215 9367
rect 5368 9364 5396 9472
rect 5813 9469 5825 9503
rect 5859 9500 5871 9503
rect 6457 9503 6515 9509
rect 6457 9500 6469 9503
rect 5859 9472 6469 9500
rect 5859 9469 5871 9472
rect 5813 9463 5871 9469
rect 6457 9469 6469 9472
rect 6503 9469 6515 9503
rect 6457 9463 6515 9469
rect 8481 9503 8539 9509
rect 8481 9469 8493 9503
rect 8527 9469 8539 9503
rect 8481 9463 8539 9469
rect 5442 9392 5448 9444
rect 5500 9432 5506 9444
rect 5828 9432 5856 9463
rect 8496 9432 8524 9463
rect 10318 9460 10324 9512
rect 10376 9500 10382 9512
rect 10612 9509 10640 9540
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9568 11943 9571
rect 12526 9568 12532 9580
rect 11931 9540 12532 9568
rect 11931 9537 11943 9540
rect 11885 9531 11943 9537
rect 10597 9503 10655 9509
rect 10597 9500 10609 9503
rect 10376 9472 10609 9500
rect 10376 9460 10382 9472
rect 10597 9469 10609 9472
rect 10643 9469 10655 9503
rect 10778 9500 10784 9512
rect 10739 9472 10784 9500
rect 10597 9463 10655 9469
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 5500 9404 5856 9432
rect 6472 9404 8524 9432
rect 11241 9435 11299 9441
rect 5500 9392 5506 9404
rect 6472 9376 6500 9404
rect 11241 9401 11253 9435
rect 11287 9432 11299 9435
rect 11900 9432 11928 9531
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12805 9571 12863 9577
rect 12805 9537 12817 9571
rect 12851 9568 12863 9571
rect 13078 9568 13084 9580
rect 12851 9540 13084 9568
rect 12851 9537 12863 9540
rect 12805 9531 12863 9537
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 18233 9571 18291 9577
rect 18233 9537 18245 9571
rect 18279 9568 18291 9571
rect 18509 9571 18567 9577
rect 18509 9568 18521 9571
rect 18279 9540 18521 9568
rect 18279 9537 18291 9540
rect 18233 9531 18291 9537
rect 18509 9537 18521 9540
rect 18555 9568 18567 9571
rect 18690 9568 18696 9580
rect 18555 9540 18696 9568
rect 18555 9537 18567 9540
rect 18509 9531 18567 9537
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 11977 9503 12035 9509
rect 11977 9469 11989 9503
rect 12023 9469 12035 9503
rect 11977 9463 12035 9469
rect 12161 9503 12219 9509
rect 12161 9469 12173 9503
rect 12207 9469 12219 9503
rect 12161 9463 12219 9469
rect 13173 9503 13231 9509
rect 13173 9469 13185 9503
rect 13219 9500 13231 9503
rect 13998 9500 14004 9512
rect 13219 9472 14004 9500
rect 13219 9469 13231 9472
rect 13173 9463 13231 9469
rect 11287 9404 11928 9432
rect 11287 9401 11299 9404
rect 11241 9395 11299 9401
rect 6270 9364 6276 9376
rect 5368 9336 6276 9364
rect 4157 9327 4215 9333
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 6454 9324 6460 9376
rect 6512 9324 6518 9376
rect 7098 9364 7104 9376
rect 7059 9336 7104 9364
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 9861 9367 9919 9373
rect 9861 9333 9873 9367
rect 9907 9364 9919 9367
rect 10502 9364 10508 9376
rect 9907 9336 10508 9364
rect 9907 9333 9919 9336
rect 9861 9327 9919 9333
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 11992 9364 12020 9463
rect 12176 9432 12204 9463
rect 13998 9460 14004 9472
rect 14056 9460 14062 9512
rect 14826 9500 14832 9512
rect 14787 9472 14832 9500
rect 14826 9460 14832 9472
rect 14884 9460 14890 9512
rect 16574 9500 16580 9512
rect 16535 9472 16580 9500
rect 16574 9460 16580 9472
rect 16632 9460 16638 9512
rect 16850 9500 16856 9512
rect 16811 9472 16856 9500
rect 16850 9460 16856 9472
rect 16908 9460 16914 9512
rect 12802 9432 12808 9444
rect 12176 9404 12808 9432
rect 12802 9392 12808 9404
rect 12860 9392 12866 9444
rect 14090 9364 14096 9376
rect 11992 9336 14096 9364
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 14366 9324 14372 9376
rect 14424 9364 14430 9376
rect 18325 9367 18383 9373
rect 18325 9364 18337 9367
rect 14424 9336 18337 9364
rect 14424 9324 14430 9336
rect 18325 9333 18337 9336
rect 18371 9333 18383 9367
rect 18325 9327 18383 9333
rect 368 9274 18860 9296
rect 368 9222 3478 9274
rect 3530 9222 3542 9274
rect 3594 9222 3606 9274
rect 3658 9222 3670 9274
rect 3722 9222 3734 9274
rect 3786 9222 6578 9274
rect 6630 9222 6642 9274
rect 6694 9222 6706 9274
rect 6758 9222 6770 9274
rect 6822 9222 6834 9274
rect 6886 9222 9678 9274
rect 9730 9222 9742 9274
rect 9794 9222 9806 9274
rect 9858 9222 9870 9274
rect 9922 9222 9934 9274
rect 9986 9222 12778 9274
rect 12830 9222 12842 9274
rect 12894 9222 12906 9274
rect 12958 9222 12970 9274
rect 13022 9222 13034 9274
rect 13086 9222 15878 9274
rect 15930 9222 15942 9274
rect 15994 9222 16006 9274
rect 16058 9222 16070 9274
rect 16122 9222 16134 9274
rect 16186 9222 18860 9274
rect 368 9200 18860 9222
rect 1121 9163 1179 9169
rect 1121 9129 1133 9163
rect 1167 9160 1179 9163
rect 1394 9160 1400 9172
rect 1167 9132 1400 9160
rect 1167 9129 1179 9132
rect 1121 9123 1179 9129
rect 1394 9120 1400 9132
rect 1452 9120 1458 9172
rect 4614 9120 4620 9172
rect 4672 9160 4678 9172
rect 6457 9163 6515 9169
rect 6457 9160 6469 9163
rect 4672 9132 6469 9160
rect 4672 9120 4678 9132
rect 6457 9129 6469 9132
rect 6503 9129 6515 9163
rect 6457 9123 6515 9129
rect 9582 9120 9588 9172
rect 9640 9160 9646 9172
rect 10597 9163 10655 9169
rect 9640 9132 10180 9160
rect 9640 9120 9646 9132
rect 1213 9027 1271 9033
rect 1213 8993 1225 9027
rect 1259 9024 1271 9027
rect 1302 9024 1308 9036
rect 1259 8996 1308 9024
rect 1259 8993 1271 8996
rect 1213 8987 1271 8993
rect 1302 8984 1308 8996
rect 1360 8984 1366 9036
rect 1412 9024 1440 9120
rect 1486 9052 1492 9104
rect 1544 9092 1550 9104
rect 2498 9092 2504 9104
rect 1544 9064 2504 9092
rect 1544 9052 1550 9064
rect 2498 9052 2504 9064
rect 2556 9052 2562 9104
rect 10152 9092 10180 9132
rect 10597 9129 10609 9163
rect 10643 9160 10655 9163
rect 10778 9160 10784 9172
rect 10643 9132 10784 9160
rect 10643 9129 10655 9132
rect 10597 9123 10655 9129
rect 10778 9120 10784 9132
rect 10836 9120 10842 9172
rect 14826 9160 14832 9172
rect 13924 9132 14832 9160
rect 10152 9064 11192 9092
rect 1412 8996 1716 9024
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 1688 8965 1716 8996
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 3142 9024 3148 9036
rect 2832 8996 3148 9024
rect 2832 8984 2838 8996
rect 3142 8984 3148 8996
rect 3200 9024 3206 9036
rect 3200 8996 3372 9024
rect 3200 8984 3206 8996
rect 3344 8965 3372 8996
rect 6270 8984 6276 9036
rect 6328 9024 6334 9036
rect 7009 9027 7067 9033
rect 7009 9024 7021 9027
rect 6328 8996 7021 9024
rect 6328 8984 6334 8996
rect 7009 8993 7021 8996
rect 7055 8993 7067 9027
rect 7009 8987 7067 8993
rect 8849 9027 8907 9033
rect 8849 8993 8861 9027
rect 8895 9024 8907 9027
rect 10134 9024 10140 9036
rect 8895 8996 10140 9024
rect 8895 8993 8907 8996
rect 8849 8987 8907 8993
rect 10134 8984 10140 8996
rect 10192 9024 10198 9036
rect 11054 9024 11060 9036
rect 10192 8996 11060 9024
rect 10192 8984 10198 8996
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 11164 9024 11192 9064
rect 13924 9024 13952 9132
rect 14826 9120 14832 9132
rect 14884 9120 14890 9172
rect 15841 9163 15899 9169
rect 15841 9129 15853 9163
rect 15887 9160 15899 9163
rect 16574 9160 16580 9172
rect 15887 9132 16580 9160
rect 15887 9129 15899 9132
rect 15841 9123 15899 9129
rect 16574 9120 16580 9132
rect 16632 9120 16638 9172
rect 14090 9024 14096 9036
rect 11164 8996 13952 9024
rect 14051 8996 14096 9024
rect 14090 8984 14096 8996
rect 14148 9024 14154 9036
rect 16025 9027 16083 9033
rect 16025 9024 16037 9027
rect 14148 8996 16037 9024
rect 14148 8984 14154 8996
rect 16025 8993 16037 8996
rect 16071 9024 16083 9027
rect 16850 9024 16856 9036
rect 16071 8996 16856 9024
rect 16071 8993 16083 8996
rect 16025 8987 16083 8993
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 1489 8959 1547 8965
rect 1489 8925 1501 8959
rect 1535 8925 1547 8959
rect 1489 8919 1547 8925
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8956 4123 8959
rect 4154 8956 4160 8968
rect 4111 8928 4160 8956
rect 4111 8925 4123 8928
rect 4065 8919 4123 8925
rect 1210 8820 1216 8832
rect 1171 8792 1216 8820
rect 1210 8780 1216 8792
rect 1268 8780 1274 8832
rect 1504 8820 1532 8919
rect 4154 8916 4160 8928
rect 4212 8916 4218 8968
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 4890 8956 4896 8968
rect 4295 8928 4896 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 4890 8916 4896 8928
rect 4948 8916 4954 8968
rect 6454 8916 6460 8968
rect 6512 8956 6518 8968
rect 7285 8959 7343 8965
rect 7285 8956 7297 8959
rect 6512 8928 7297 8956
rect 6512 8916 6518 8928
rect 7285 8925 7297 8928
rect 7331 8925 7343 8959
rect 7285 8919 7343 8925
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 11241 8959 11299 8965
rect 11241 8956 11253 8959
rect 11204 8928 11253 8956
rect 11204 8916 11210 8928
rect 11241 8925 11253 8928
rect 11287 8925 11299 8959
rect 16390 8956 16396 8968
rect 16351 8928 16396 8956
rect 11241 8919 11299 8925
rect 16390 8916 16396 8928
rect 16448 8916 16454 8968
rect 2866 8888 2872 8900
rect 2779 8860 2872 8888
rect 2866 8848 2872 8860
rect 2924 8888 2930 8900
rect 3970 8888 3976 8900
rect 2924 8860 3976 8888
rect 2924 8848 2930 8860
rect 3970 8848 3976 8860
rect 4028 8848 4034 8900
rect 6825 8891 6883 8897
rect 6825 8857 6837 8891
rect 6871 8888 6883 8891
rect 7098 8888 7104 8900
rect 6871 8860 7104 8888
rect 6871 8857 6883 8860
rect 6825 8851 6883 8857
rect 7098 8848 7104 8860
rect 7156 8848 7162 8900
rect 7552 8891 7610 8897
rect 7552 8857 7564 8891
rect 7598 8888 7610 8891
rect 9122 8888 9128 8900
rect 7598 8860 8984 8888
rect 9083 8860 9128 8888
rect 7598 8857 7610 8860
rect 7552 8851 7610 8857
rect 3234 8820 3240 8832
rect 1504 8792 3240 8820
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 3326 8780 3332 8832
rect 3384 8820 3390 8832
rect 4157 8823 4215 8829
rect 4157 8820 4169 8823
rect 3384 8792 4169 8820
rect 3384 8780 3390 8792
rect 4157 8789 4169 8792
rect 4203 8789 4215 8823
rect 4157 8783 4215 8789
rect 6362 8780 6368 8832
rect 6420 8820 6426 8832
rect 6917 8823 6975 8829
rect 6917 8820 6929 8823
rect 6420 8792 6929 8820
rect 6420 8780 6426 8792
rect 6917 8789 6929 8792
rect 6963 8789 6975 8823
rect 6917 8783 6975 8789
rect 8665 8823 8723 8829
rect 8665 8789 8677 8823
rect 8711 8820 8723 8823
rect 8846 8820 8852 8832
rect 8711 8792 8852 8820
rect 8711 8789 8723 8792
rect 8665 8783 8723 8789
rect 8846 8780 8852 8792
rect 8904 8780 8910 8832
rect 8956 8820 8984 8860
rect 9122 8848 9128 8860
rect 9180 8848 9186 8900
rect 11517 8891 11575 8897
rect 9214 8820 9220 8832
rect 8956 8792 9220 8820
rect 9214 8780 9220 8792
rect 9272 8780 9278 8832
rect 9306 8780 9312 8832
rect 9364 8820 9370 8832
rect 10336 8820 10364 8874
rect 11517 8857 11529 8891
rect 11563 8888 11575 8891
rect 11606 8888 11612 8900
rect 11563 8860 11612 8888
rect 11563 8857 11575 8860
rect 11517 8851 11575 8857
rect 11606 8848 11612 8860
rect 11664 8848 11670 8900
rect 12066 8848 12072 8900
rect 12124 8848 12130 8900
rect 13265 8891 13323 8897
rect 13265 8857 13277 8891
rect 13311 8857 13323 8891
rect 14366 8888 14372 8900
rect 14327 8860 14372 8888
rect 13265 8851 13323 8857
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 9364 8792 11069 8820
rect 9364 8780 9370 8792
rect 11057 8789 11069 8792
rect 11103 8820 11115 8823
rect 12084 8820 12112 8848
rect 11103 8792 12112 8820
rect 11103 8789 11115 8792
rect 11057 8783 11115 8789
rect 12158 8780 12164 8832
rect 12216 8820 12222 8832
rect 13280 8820 13308 8851
rect 14366 8848 14372 8860
rect 14424 8848 14430 8900
rect 12216 8792 13308 8820
rect 14001 8823 14059 8829
rect 12216 8780 12222 8792
rect 14001 8789 14013 8823
rect 14047 8820 14059 8823
rect 14182 8820 14188 8832
rect 14047 8792 14188 8820
rect 14047 8789 14059 8792
rect 14001 8783 14059 8789
rect 14182 8780 14188 8792
rect 14240 8820 14246 8832
rect 14844 8820 14872 8874
rect 17126 8848 17132 8900
rect 17184 8848 17190 8900
rect 18138 8820 18144 8832
rect 14240 8792 14872 8820
rect 18099 8792 18144 8820
rect 14240 8780 14246 8792
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 368 8730 18860 8752
rect 368 8678 5028 8730
rect 5080 8678 5092 8730
rect 5144 8678 5156 8730
rect 5208 8678 5220 8730
rect 5272 8678 5284 8730
rect 5336 8678 8128 8730
rect 8180 8678 8192 8730
rect 8244 8678 8256 8730
rect 8308 8678 8320 8730
rect 8372 8678 8384 8730
rect 8436 8678 11228 8730
rect 11280 8678 11292 8730
rect 11344 8678 11356 8730
rect 11408 8678 11420 8730
rect 11472 8678 11484 8730
rect 11536 8678 14328 8730
rect 14380 8678 14392 8730
rect 14444 8678 14456 8730
rect 14508 8678 14520 8730
rect 14572 8678 14584 8730
rect 14636 8678 17428 8730
rect 17480 8678 17492 8730
rect 17544 8678 17556 8730
rect 17608 8678 17620 8730
rect 17672 8678 17684 8730
rect 17736 8678 18860 8730
rect 368 8656 18860 8678
rect 1302 8576 1308 8628
rect 1360 8616 1366 8628
rect 2869 8619 2927 8625
rect 2869 8616 2881 8619
rect 1360 8588 2881 8616
rect 1360 8576 1366 8588
rect 2869 8585 2881 8588
rect 2915 8585 2927 8619
rect 2869 8579 2927 8585
rect 3234 8576 3240 8628
rect 3292 8616 3298 8628
rect 4433 8619 4491 8625
rect 4433 8616 4445 8619
rect 3292 8588 4445 8616
rect 3292 8576 3298 8588
rect 4433 8585 4445 8588
rect 4479 8585 4491 8619
rect 5442 8616 5448 8628
rect 4433 8579 4491 8585
rect 4816 8588 5448 8616
rect 937 8551 995 8557
rect 937 8517 949 8551
rect 983 8548 995 8551
rect 1210 8548 1216 8560
rect 983 8520 1216 8548
rect 983 8517 995 8520
rect 937 8511 995 8517
rect 1210 8508 1216 8520
rect 1268 8508 1274 8560
rect 2498 8508 2504 8560
rect 2556 8548 2562 8560
rect 2556 8520 3464 8548
rect 2556 8508 2562 8520
rect 658 8480 664 8492
rect 619 8452 664 8480
rect 658 8440 664 8452
rect 716 8440 722 8492
rect 2869 8483 2927 8489
rect 2056 8344 2084 8466
rect 2869 8449 2881 8483
rect 2915 8449 2927 8483
rect 3050 8480 3056 8492
rect 3011 8452 3056 8480
rect 2869 8443 2927 8449
rect 2409 8415 2467 8421
rect 2409 8381 2421 8415
rect 2455 8412 2467 8415
rect 2774 8412 2780 8424
rect 2455 8384 2780 8412
rect 2455 8381 2467 8384
rect 2409 8375 2467 8381
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 2884 8412 2912 8443
rect 3050 8440 3056 8452
rect 3108 8440 3114 8492
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8480 3203 8483
rect 3326 8480 3332 8492
rect 3191 8452 3332 8480
rect 3191 8449 3203 8452
rect 3145 8443 3203 8449
rect 3160 8412 3188 8443
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 3436 8489 3464 8520
rect 3421 8483 3479 8489
rect 3421 8449 3433 8483
rect 3467 8449 3479 8483
rect 4816 8480 4844 8588
rect 5442 8576 5448 8588
rect 5500 8616 5506 8628
rect 8205 8619 8263 8625
rect 8205 8616 8217 8619
rect 5500 8588 5764 8616
rect 5500 8576 5506 8588
rect 4890 8508 4896 8560
rect 4948 8548 4954 8560
rect 4948 8520 5580 8548
rect 4948 8508 4954 8520
rect 5350 8480 5356 8492
rect 3421 8443 3479 8449
rect 4264 8452 4844 8480
rect 5311 8452 5356 8480
rect 4264 8421 4292 8452
rect 5350 8440 5356 8452
rect 5408 8440 5414 8492
rect 5552 8489 5580 8520
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8449 5595 8483
rect 5537 8443 5595 8449
rect 2884 8384 3188 8412
rect 4249 8415 4307 8421
rect 4249 8381 4261 8415
rect 4295 8381 4307 8415
rect 4249 8375 4307 8381
rect 4338 8372 4344 8424
rect 4396 8412 4402 8424
rect 5736 8412 5764 8588
rect 6104 8588 8217 8616
rect 6104 8557 6132 8588
rect 8205 8585 8217 8588
rect 8251 8585 8263 8619
rect 8205 8579 8263 8585
rect 8757 8619 8815 8625
rect 8757 8585 8769 8619
rect 8803 8616 8815 8619
rect 9306 8616 9312 8628
rect 8803 8588 9312 8616
rect 8803 8585 8815 8588
rect 8757 8579 8815 8585
rect 6089 8551 6147 8557
rect 6089 8548 6101 8551
rect 5828 8520 6101 8548
rect 5828 8489 5856 8520
rect 6089 8517 6101 8520
rect 6135 8517 6147 8551
rect 6089 8511 6147 8517
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8449 5963 8483
rect 6178 8474 6184 8526
rect 6236 8474 6242 8526
rect 8386 8508 8392 8560
rect 8444 8548 8450 8560
rect 8570 8548 8576 8560
rect 8444 8520 8576 8548
rect 8444 8508 8450 8520
rect 8570 8508 8576 8520
rect 8628 8548 8634 8560
rect 8772 8548 8800 8579
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 9585 8619 9643 8625
rect 9585 8585 9597 8619
rect 9631 8616 9643 8619
rect 11517 8619 11575 8625
rect 9631 8588 10180 8616
rect 9631 8585 9643 8588
rect 9585 8579 9643 8585
rect 8628 8520 8800 8548
rect 8864 8520 9720 8548
rect 8628 8508 8634 8520
rect 8864 8492 8892 8520
rect 6273 8483 6331 8489
rect 6179 8471 6191 8474
rect 6225 8471 6237 8474
rect 6179 8465 6237 8471
rect 5905 8443 5963 8449
rect 6273 8449 6285 8483
rect 6319 8449 6331 8483
rect 6273 8443 6331 8449
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 7558 8480 7564 8492
rect 6595 8452 7564 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 5920 8412 5948 8443
rect 4396 8384 4441 8412
rect 5736 8384 5948 8412
rect 4396 8372 4402 8384
rect 2593 8347 2651 8353
rect 2593 8344 2605 8347
rect 2056 8316 2605 8344
rect 2593 8313 2605 8316
rect 2639 8344 2651 8347
rect 2866 8344 2872 8356
rect 2639 8316 2872 8344
rect 2639 8313 2651 8316
rect 2593 8307 2651 8313
rect 2866 8304 2872 8316
rect 2924 8304 2930 8356
rect 6181 8347 6239 8353
rect 6181 8313 6193 8347
rect 6227 8344 6239 8347
rect 6288 8344 6316 8443
rect 6227 8316 6316 8344
rect 6227 8313 6239 8316
rect 6181 8307 6239 8313
rect 4798 8276 4804 8288
rect 4759 8248 4804 8276
rect 4798 8236 4804 8248
rect 4856 8236 4862 8288
rect 5537 8279 5595 8285
rect 5537 8245 5549 8279
rect 5583 8276 5595 8279
rect 6380 8276 6408 8443
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8480 8355 8483
rect 8478 8480 8484 8492
rect 8343 8452 8484 8480
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 8478 8440 8484 8452
rect 8536 8440 8542 8492
rect 8846 8480 8852 8492
rect 8807 8452 8852 8480
rect 8846 8440 8852 8452
rect 8904 8440 8910 8492
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8480 9091 8483
rect 9214 8480 9220 8492
rect 9079 8452 9220 8480
rect 9079 8449 9091 8452
rect 9033 8443 9091 8449
rect 9214 8440 9220 8452
rect 9272 8440 9278 8492
rect 9692 8489 9720 8520
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8480 9367 8483
rect 9677 8483 9735 8489
rect 9355 8452 9536 8480
rect 9355 8449 9367 8452
rect 9309 8443 9367 8449
rect 6457 8347 6515 8353
rect 6457 8313 6469 8347
rect 6503 8344 6515 8347
rect 7098 8344 7104 8356
rect 6503 8316 7104 8344
rect 6503 8313 6515 8316
rect 6457 8307 6515 8313
rect 7098 8304 7104 8316
rect 7156 8304 7162 8356
rect 9217 8347 9275 8353
rect 9217 8313 9229 8347
rect 9263 8344 9275 8347
rect 9401 8347 9459 8353
rect 9401 8344 9413 8347
rect 9263 8316 9413 8344
rect 9263 8313 9275 8316
rect 9217 8307 9275 8313
rect 9401 8313 9413 8316
rect 9447 8313 9459 8347
rect 9508 8344 9536 8452
rect 9677 8449 9689 8483
rect 9723 8449 9735 8483
rect 9677 8443 9735 8449
rect 9766 8440 9772 8492
rect 9824 8480 9830 8492
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 9824 8452 9873 8480
rect 9824 8440 9830 8452
rect 9861 8449 9873 8452
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8412 9643 8415
rect 10042 8412 10048 8424
rect 9631 8384 10048 8412
rect 9631 8381 9643 8384
rect 9585 8375 9643 8381
rect 10042 8372 10048 8384
rect 10100 8372 10106 8424
rect 9861 8347 9919 8353
rect 9861 8344 9873 8347
rect 9508 8316 9873 8344
rect 9401 8307 9459 8313
rect 9861 8313 9873 8316
rect 9907 8313 9919 8347
rect 10152 8344 10180 8588
rect 11517 8585 11529 8619
rect 11563 8616 11575 8619
rect 11606 8616 11612 8628
rect 11563 8588 11612 8616
rect 11563 8585 11575 8588
rect 11517 8579 11575 8585
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 11716 8588 16344 8616
rect 11716 8548 11744 8588
rect 10428 8520 11744 8548
rect 10428 8492 10456 8520
rect 14090 8508 14096 8560
rect 14148 8548 14154 8560
rect 14148 8520 14872 8548
rect 14148 8508 14154 8520
rect 10410 8480 10416 8492
rect 10323 8452 10416 8480
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10778 8440 10784 8492
rect 10836 8480 10842 8492
rect 10965 8483 11023 8489
rect 10965 8480 10977 8483
rect 10836 8452 10977 8480
rect 10836 8440 10842 8452
rect 10965 8449 10977 8452
rect 11011 8449 11023 8483
rect 10965 8443 11023 8449
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 11296 8452 11713 8480
rect 11296 8440 11302 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 13814 8440 13820 8492
rect 13872 8489 13878 8492
rect 14844 8489 14872 8520
rect 15562 8508 15568 8560
rect 15620 8508 15626 8560
rect 16316 8548 16344 8588
rect 16390 8576 16396 8628
rect 16448 8616 16454 8628
rect 16623 8619 16681 8625
rect 16623 8616 16635 8619
rect 16448 8588 16635 8616
rect 16448 8576 16454 8588
rect 16623 8585 16635 8588
rect 16669 8585 16681 8619
rect 16623 8579 16681 8585
rect 18138 8548 18144 8560
rect 16316 8520 18144 8548
rect 18138 8508 18144 8520
rect 18196 8548 18202 8560
rect 18233 8551 18291 8557
rect 18233 8548 18245 8551
rect 18196 8520 18245 8548
rect 18196 8508 18202 8520
rect 18233 8517 18245 8520
rect 18279 8517 18291 8551
rect 18233 8511 18291 8517
rect 13872 8480 13884 8489
rect 14829 8483 14887 8489
rect 13872 8452 13917 8480
rect 13872 8443 13884 8452
rect 14829 8449 14841 8483
rect 14875 8449 14887 8483
rect 14829 8443 14887 8449
rect 17957 8483 18015 8489
rect 17957 8449 17969 8483
rect 18003 8449 18015 8483
rect 17957 8443 18015 8449
rect 13872 8440 13878 8443
rect 10873 8415 10931 8421
rect 10873 8381 10885 8415
rect 10919 8412 10931 8415
rect 11606 8412 11612 8424
rect 10919 8384 11612 8412
rect 10919 8381 10931 8384
rect 10873 8375 10931 8381
rect 11606 8372 11612 8384
rect 11664 8372 11670 8424
rect 11882 8372 11888 8424
rect 11940 8412 11946 8424
rect 11977 8415 12035 8421
rect 11977 8412 11989 8415
rect 11940 8384 11989 8412
rect 11940 8372 11946 8384
rect 11977 8381 11989 8384
rect 12023 8381 12035 8415
rect 11977 8375 12035 8381
rect 14093 8415 14151 8421
rect 14093 8381 14105 8415
rect 14139 8381 14151 8415
rect 14093 8375 14151 8381
rect 15197 8415 15255 8421
rect 15197 8381 15209 8415
rect 15243 8412 15255 8415
rect 17972 8412 18000 8443
rect 15243 8384 17816 8412
rect 17972 8384 18552 8412
rect 15243 8381 15255 8384
rect 15197 8375 15255 8381
rect 10152 8316 11928 8344
rect 9861 8307 9919 8313
rect 5583 8248 6408 8276
rect 5583 8245 5595 8248
rect 5537 8239 5595 8245
rect 6914 8236 6920 8288
rect 6972 8276 6978 8288
rect 8202 8276 8208 8288
rect 6972 8248 8208 8276
rect 6972 8236 6978 8248
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 10502 8276 10508 8288
rect 10463 8248 10508 8276
rect 10502 8236 10508 8248
rect 10560 8276 10566 8288
rect 10778 8276 10784 8288
rect 10560 8248 10784 8276
rect 10560 8236 10566 8248
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 10962 8236 10968 8288
rect 11020 8276 11026 8288
rect 11241 8279 11299 8285
rect 11241 8276 11253 8279
rect 11020 8248 11253 8276
rect 11020 8236 11026 8248
rect 11241 8245 11253 8248
rect 11287 8276 11299 8279
rect 11330 8276 11336 8288
rect 11287 8248 11336 8276
rect 11287 8245 11299 8248
rect 11241 8239 11299 8245
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 11425 8279 11483 8285
rect 11425 8245 11437 8279
rect 11471 8276 11483 8279
rect 11790 8276 11796 8288
rect 11471 8248 11796 8276
rect 11471 8245 11483 8248
rect 11425 8239 11483 8245
rect 11790 8236 11796 8248
rect 11848 8236 11854 8288
rect 11900 8285 11928 8316
rect 11885 8279 11943 8285
rect 11885 8245 11897 8279
rect 11931 8245 11943 8279
rect 11885 8239 11943 8245
rect 12066 8236 12072 8288
rect 12124 8276 12130 8288
rect 12713 8279 12771 8285
rect 12713 8276 12725 8279
rect 12124 8248 12725 8276
rect 12124 8236 12130 8248
rect 12713 8245 12725 8248
rect 12759 8245 12771 8279
rect 12713 8239 12771 8245
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 14108 8276 14136 8375
rect 16761 8347 16819 8353
rect 16761 8313 16773 8347
rect 16807 8344 16819 8347
rect 17126 8344 17132 8356
rect 16807 8316 17132 8344
rect 16807 8313 16819 8316
rect 16761 8307 16819 8313
rect 17126 8304 17132 8316
rect 17184 8304 17190 8356
rect 17788 8353 17816 8384
rect 18524 8353 18552 8384
rect 17773 8347 17831 8353
rect 17773 8313 17785 8347
rect 17819 8313 17831 8347
rect 17773 8307 17831 8313
rect 18509 8347 18567 8353
rect 18509 8313 18521 8347
rect 18555 8344 18567 8347
rect 18598 8344 18604 8356
rect 18555 8316 18604 8344
rect 18555 8313 18567 8316
rect 18509 8307 18567 8313
rect 18598 8304 18604 8316
rect 18656 8304 18662 8356
rect 13504 8248 14136 8276
rect 13504 8236 13510 8248
rect 14182 8236 14188 8288
rect 14240 8276 14246 8288
rect 14645 8279 14703 8285
rect 14645 8276 14657 8279
rect 14240 8248 14657 8276
rect 14240 8236 14246 8248
rect 14645 8245 14657 8248
rect 14691 8276 14703 8279
rect 15378 8276 15384 8288
rect 14691 8248 15384 8276
rect 14691 8245 14703 8248
rect 14645 8239 14703 8245
rect 15378 8236 15384 8248
rect 15436 8236 15442 8288
rect 16850 8236 16856 8288
rect 16908 8276 16914 8288
rect 18141 8279 18199 8285
rect 18141 8276 18153 8279
rect 16908 8248 18153 8276
rect 16908 8236 16914 8248
rect 18141 8245 18153 8248
rect 18187 8245 18199 8279
rect 18141 8239 18199 8245
rect 368 8186 18860 8208
rect 368 8134 3478 8186
rect 3530 8134 3542 8186
rect 3594 8134 3606 8186
rect 3658 8134 3670 8186
rect 3722 8134 3734 8186
rect 3786 8134 6578 8186
rect 6630 8134 6642 8186
rect 6694 8134 6706 8186
rect 6758 8134 6770 8186
rect 6822 8134 6834 8186
rect 6886 8134 9678 8186
rect 9730 8134 9742 8186
rect 9794 8134 9806 8186
rect 9858 8134 9870 8186
rect 9922 8134 9934 8186
rect 9986 8134 12778 8186
rect 12830 8134 12842 8186
rect 12894 8134 12906 8186
rect 12958 8134 12970 8186
rect 13022 8134 13034 8186
rect 13086 8134 15878 8186
rect 15930 8134 15942 8186
rect 15994 8134 16006 8186
rect 16058 8134 16070 8186
rect 16122 8134 16134 8186
rect 16186 8134 18860 8186
rect 368 8112 18860 8134
rect 3050 8032 3056 8084
rect 3108 8072 3114 8084
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 3108 8044 4077 8072
rect 3108 8032 3114 8044
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 4890 8072 4896 8084
rect 4851 8044 4896 8072
rect 4065 8035 4123 8041
rect 4890 8032 4896 8044
rect 4948 8032 4954 8084
rect 5261 8075 5319 8081
rect 5261 8041 5273 8075
rect 5307 8072 5319 8075
rect 5629 8075 5687 8081
rect 5629 8072 5641 8075
rect 5307 8044 5641 8072
rect 5307 8041 5319 8044
rect 5261 8035 5319 8041
rect 5629 8041 5641 8044
rect 5675 8072 5687 8075
rect 5994 8072 6000 8084
rect 5675 8044 6000 8072
rect 5675 8041 5687 8044
rect 5629 8035 5687 8041
rect 5994 8032 6000 8044
rect 6052 8032 6058 8084
rect 6362 8032 6368 8084
rect 6420 8072 6426 8084
rect 6420 8044 7972 8072
rect 6420 8032 6426 8044
rect 2777 8007 2835 8013
rect 2777 7973 2789 8007
rect 2823 8004 2835 8007
rect 6273 8007 6331 8013
rect 2823 7976 5028 8004
rect 2823 7973 2835 7976
rect 2777 7967 2835 7973
rect 3789 7939 3847 7945
rect 3789 7905 3801 7939
rect 3835 7936 3847 7939
rect 4154 7936 4160 7948
rect 3835 7908 4160 7936
rect 3835 7905 3847 7908
rect 3789 7899 3847 7905
rect 4154 7896 4160 7908
rect 4212 7896 4218 7948
rect 4706 7936 4712 7948
rect 4356 7908 4712 7936
rect 1486 7828 1492 7880
rect 1544 7868 1550 7880
rect 2041 7871 2099 7877
rect 2041 7868 2053 7871
rect 1544 7840 2053 7868
rect 1544 7828 1550 7840
rect 2041 7837 2053 7840
rect 2087 7837 2099 7871
rect 2222 7868 2228 7880
rect 2183 7840 2228 7868
rect 2041 7831 2099 7837
rect 2056 7800 2084 7831
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 2590 7868 2596 7880
rect 2551 7840 2596 7868
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 3142 7868 3148 7880
rect 2823 7840 3148 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 3326 7828 3332 7880
rect 3384 7868 3390 7880
rect 3697 7871 3755 7877
rect 3697 7868 3709 7871
rect 3384 7840 3709 7868
rect 3384 7828 3390 7840
rect 3697 7837 3709 7840
rect 3743 7868 3755 7871
rect 4356 7868 4384 7908
rect 4706 7896 4712 7908
rect 4764 7896 4770 7948
rect 5000 7945 5028 7976
rect 5460 7976 5856 8004
rect 5460 7945 5488 7976
rect 4985 7939 5043 7945
rect 4985 7905 4997 7939
rect 5031 7905 5043 7939
rect 4985 7899 5043 7905
rect 5077 7939 5135 7945
rect 5077 7905 5089 7939
rect 5123 7936 5135 7939
rect 5445 7939 5503 7945
rect 5445 7936 5457 7939
rect 5123 7908 5457 7936
rect 5123 7905 5135 7908
rect 5077 7899 5135 7905
rect 5445 7905 5457 7908
rect 5491 7905 5503 7939
rect 5828 7936 5856 7976
rect 6273 7973 6285 8007
rect 6319 8004 6331 8007
rect 6822 8004 6828 8016
rect 6319 7976 6828 8004
rect 6319 7973 6331 7976
rect 6273 7967 6331 7973
rect 6822 7964 6828 7976
rect 6880 7964 6886 8016
rect 7944 8004 7972 8044
rect 9490 8032 9496 8084
rect 9548 8072 9554 8084
rect 10962 8072 10968 8084
rect 9548 8044 10968 8072
rect 9548 8032 9554 8044
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 18506 8072 18512 8084
rect 11072 8044 18512 8072
rect 9766 8004 9772 8016
rect 7944 7976 9772 8004
rect 9766 7964 9772 7976
rect 9824 8004 9830 8016
rect 10410 8004 10416 8016
rect 9824 7976 10416 8004
rect 9824 7964 9830 7976
rect 10410 7964 10416 7976
rect 10468 7964 10474 8016
rect 5445 7899 5503 7905
rect 5552 7908 5764 7936
rect 5828 7908 7052 7936
rect 3743 7840 4384 7868
rect 4433 7871 4491 7877
rect 3743 7837 3755 7840
rect 3697 7831 3755 7837
rect 4433 7837 4445 7871
rect 4479 7868 4491 7871
rect 4798 7868 4804 7880
rect 4479 7840 4804 7868
rect 4479 7837 4491 7840
rect 4433 7831 4491 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 2682 7800 2688 7812
rect 2056 7772 2688 7800
rect 2682 7760 2688 7772
rect 2740 7760 2746 7812
rect 4338 7760 4344 7812
rect 4396 7800 4402 7812
rect 4525 7803 4583 7809
rect 4525 7800 4537 7803
rect 4396 7772 4537 7800
rect 4396 7760 4402 7772
rect 4525 7769 4537 7772
rect 4571 7800 4583 7803
rect 5092 7800 5120 7899
rect 5353 7871 5411 7877
rect 5353 7837 5365 7871
rect 5399 7868 5411 7871
rect 5552 7868 5580 7908
rect 5736 7877 5764 7908
rect 5399 7840 5580 7868
rect 5721 7871 5779 7877
rect 5399 7837 5411 7840
rect 5353 7831 5411 7837
rect 5721 7837 5733 7871
rect 5767 7868 5779 7871
rect 6362 7868 6368 7880
rect 5767 7840 6368 7868
rect 5767 7837 5779 7840
rect 5721 7831 5779 7837
rect 6362 7828 6368 7840
rect 6420 7828 6426 7880
rect 6822 7868 6828 7880
rect 6783 7840 6828 7868
rect 6822 7828 6828 7840
rect 6880 7828 6886 7880
rect 7024 7868 7052 7908
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7193 7939 7251 7945
rect 7193 7936 7205 7939
rect 7156 7908 7205 7936
rect 7156 7896 7162 7908
rect 7193 7905 7205 7908
rect 7239 7905 7251 7939
rect 9582 7936 9588 7948
rect 7193 7899 7251 7905
rect 7300 7908 9588 7936
rect 7300 7868 7328 7908
rect 9582 7896 9588 7908
rect 9640 7896 9646 7948
rect 11072 7880 11100 8044
rect 18506 8032 18512 8044
rect 18564 8032 18570 8084
rect 14090 7964 14096 8016
rect 14148 8004 14154 8016
rect 14277 8007 14335 8013
rect 14277 8004 14289 8007
rect 14148 7976 14289 8004
rect 14148 7964 14154 7976
rect 14277 7973 14289 7976
rect 14323 8004 14335 8007
rect 14323 7976 16252 8004
rect 14323 7973 14335 7976
rect 14277 7967 14335 7973
rect 11146 7896 11152 7948
rect 11204 7936 11210 7948
rect 11241 7939 11299 7945
rect 11241 7936 11253 7939
rect 11204 7908 11253 7936
rect 11204 7896 11210 7908
rect 11241 7905 11253 7908
rect 11287 7936 11299 7939
rect 13446 7936 13452 7948
rect 11287 7908 13452 7936
rect 11287 7905 11299 7908
rect 11241 7899 11299 7905
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 14734 7936 14740 7948
rect 14695 7908 14740 7936
rect 14734 7896 14740 7908
rect 14792 7896 14798 7948
rect 14918 7896 14924 7948
rect 14976 7936 14982 7948
rect 16224 7945 16252 7976
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 14976 7908 15669 7936
rect 14976 7896 14982 7908
rect 15657 7905 15669 7908
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 16209 7939 16267 7945
rect 16209 7905 16221 7939
rect 16255 7936 16267 7939
rect 17034 7936 17040 7948
rect 16255 7908 17040 7936
rect 16255 7905 16267 7908
rect 16209 7899 16267 7905
rect 17034 7896 17040 7908
rect 17092 7896 17098 7948
rect 11054 7868 11060 7880
rect 7024 7840 7328 7868
rect 10967 7840 11060 7868
rect 11054 7828 11060 7840
rect 11112 7828 11118 7880
rect 11606 7868 11612 7880
rect 11567 7840 11612 7868
rect 11606 7828 11612 7840
rect 11664 7828 11670 7880
rect 12802 7828 12808 7880
rect 12860 7868 12866 7880
rect 13035 7871 13093 7877
rect 13035 7868 13047 7871
rect 12860 7840 13047 7868
rect 12860 7828 12866 7840
rect 13035 7837 13047 7840
rect 13081 7868 13093 7871
rect 13633 7871 13691 7877
rect 13633 7868 13645 7871
rect 13081 7840 13645 7868
rect 13081 7837 13093 7840
rect 13035 7831 13093 7837
rect 13633 7837 13645 7840
rect 13679 7837 13691 7871
rect 13998 7868 14004 7880
rect 13959 7840 14004 7868
rect 13633 7831 13691 7837
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 14182 7868 14188 7880
rect 14143 7840 14188 7868
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 14829 7871 14887 7877
rect 14829 7837 14841 7871
rect 14875 7837 14887 7871
rect 14829 7831 14887 7837
rect 4571 7772 5120 7800
rect 5445 7803 5503 7809
rect 4571 7769 4583 7772
rect 4525 7763 4583 7769
rect 5445 7769 5457 7803
rect 5491 7800 5503 7803
rect 5902 7800 5908 7812
rect 5491 7772 5908 7800
rect 5491 7769 5503 7772
rect 5445 7763 5503 7769
rect 5902 7760 5908 7772
rect 5960 7760 5966 7812
rect 6454 7800 6460 7812
rect 6415 7772 6460 7800
rect 6454 7760 6460 7772
rect 6512 7760 6518 7812
rect 6641 7803 6699 7809
rect 6641 7769 6653 7803
rect 6687 7769 6699 7803
rect 6641 7763 6699 7769
rect 2225 7735 2283 7741
rect 2225 7701 2237 7735
rect 2271 7732 2283 7735
rect 2406 7732 2412 7744
rect 2271 7704 2412 7732
rect 2271 7701 2283 7704
rect 2225 7695 2283 7701
rect 2406 7692 2412 7704
rect 2464 7692 2470 7744
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 5997 7735 6055 7741
rect 5997 7732 6009 7735
rect 5592 7704 6009 7732
rect 5592 7692 5598 7704
rect 5997 7701 6009 7704
rect 6043 7701 6055 7735
rect 6656 7732 6684 7763
rect 8202 7760 8208 7812
rect 8260 7760 8266 7812
rect 8312 7772 9812 7800
rect 8312 7732 8340 7772
rect 6656 7704 8340 7732
rect 5997 7695 6055 7701
rect 8478 7692 8484 7744
rect 8536 7732 8542 7744
rect 8619 7735 8677 7741
rect 8619 7732 8631 7735
rect 8536 7704 8631 7732
rect 8536 7692 8542 7704
rect 8619 7701 8631 7704
rect 8665 7732 8677 7735
rect 9122 7732 9128 7744
rect 8665 7704 9128 7732
rect 8665 7701 8677 7704
rect 8619 7695 8677 7701
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 9784 7741 9812 7772
rect 12342 7760 12348 7812
rect 12400 7760 12406 7812
rect 13265 7803 13323 7809
rect 13265 7800 13277 7803
rect 12820 7772 13277 7800
rect 9769 7735 9827 7741
rect 9769 7701 9781 7735
rect 9815 7732 9827 7735
rect 12820 7732 12848 7772
rect 13265 7769 13277 7772
rect 13311 7769 13323 7803
rect 13446 7800 13452 7812
rect 13407 7772 13452 7800
rect 13265 7763 13323 7769
rect 13446 7760 13452 7772
rect 13504 7760 13510 7812
rect 14844 7800 14872 7831
rect 15378 7828 15384 7880
rect 15436 7868 15442 7880
rect 16025 7871 16083 7877
rect 16025 7868 16037 7871
rect 15436 7840 16037 7868
rect 15436 7828 15442 7840
rect 16025 7837 16037 7840
rect 16071 7837 16083 7871
rect 16025 7831 16083 7837
rect 15565 7803 15623 7809
rect 14844 7772 15148 7800
rect 13722 7732 13728 7744
rect 9815 7704 12848 7732
rect 13683 7704 13728 7732
rect 9815 7701 9827 7704
rect 9769 7695 9827 7701
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 15120 7741 15148 7772
rect 15565 7769 15577 7803
rect 15611 7800 15623 7803
rect 16390 7800 16396 7812
rect 15611 7772 16396 7800
rect 15611 7769 15623 7772
rect 15565 7763 15623 7769
rect 16390 7760 16396 7772
rect 16448 7760 16454 7812
rect 16485 7803 16543 7809
rect 16485 7769 16497 7803
rect 16531 7769 16543 7803
rect 16485 7763 16543 7769
rect 15105 7735 15163 7741
rect 15105 7701 15117 7735
rect 15151 7701 15163 7735
rect 15105 7695 15163 7701
rect 15194 7692 15200 7744
rect 15252 7732 15258 7744
rect 15473 7735 15531 7741
rect 15473 7732 15485 7735
rect 15252 7704 15485 7732
rect 15252 7692 15258 7704
rect 15473 7701 15485 7704
rect 15519 7701 15531 7735
rect 15473 7695 15531 7701
rect 16114 7692 16120 7744
rect 16172 7732 16178 7744
rect 16500 7732 16528 7763
rect 17126 7760 17132 7812
rect 17184 7760 17190 7812
rect 17862 7760 17868 7812
rect 17920 7800 17926 7812
rect 18233 7803 18291 7809
rect 18233 7800 18245 7803
rect 17920 7772 18245 7800
rect 17920 7760 17926 7772
rect 18233 7769 18245 7772
rect 18279 7769 18291 7803
rect 18233 7763 18291 7769
rect 16172 7704 16528 7732
rect 16172 7692 16178 7704
rect 368 7642 18860 7664
rect 368 7590 5028 7642
rect 5080 7590 5092 7642
rect 5144 7590 5156 7642
rect 5208 7590 5220 7642
rect 5272 7590 5284 7642
rect 5336 7590 8128 7642
rect 8180 7590 8192 7642
rect 8244 7590 8256 7642
rect 8308 7590 8320 7642
rect 8372 7590 8384 7642
rect 8436 7590 11228 7642
rect 11280 7590 11292 7642
rect 11344 7590 11356 7642
rect 11408 7590 11420 7642
rect 11472 7590 11484 7642
rect 11536 7590 14328 7642
rect 14380 7590 14392 7642
rect 14444 7590 14456 7642
rect 14508 7590 14520 7642
rect 14572 7590 14584 7642
rect 14636 7590 17428 7642
rect 17480 7590 17492 7642
rect 17544 7590 17556 7642
rect 17608 7590 17620 7642
rect 17672 7590 17684 7642
rect 17736 7590 18860 7642
rect 368 7568 18860 7590
rect 2222 7488 2228 7540
rect 2280 7528 2286 7540
rect 2593 7531 2651 7537
rect 2593 7528 2605 7531
rect 2280 7500 2605 7528
rect 2280 7488 2286 7500
rect 2593 7497 2605 7500
rect 2639 7497 2651 7531
rect 2593 7491 2651 7497
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 2961 7531 3019 7537
rect 2961 7528 2973 7531
rect 2740 7500 2973 7528
rect 2740 7488 2746 7500
rect 2961 7497 2973 7500
rect 3007 7497 3019 7531
rect 2961 7491 3019 7497
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 4212 7500 6132 7528
rect 4212 7488 4218 7500
rect 2406 7420 2412 7472
rect 2464 7460 2470 7472
rect 6104 7460 6132 7500
rect 6178 7488 6184 7540
rect 6236 7528 6242 7540
rect 6549 7531 6607 7537
rect 6549 7528 6561 7531
rect 6236 7500 6561 7528
rect 6236 7488 6242 7500
rect 6549 7497 6561 7500
rect 6595 7497 6607 7531
rect 6549 7491 6607 7497
rect 6822 7488 6828 7540
rect 6880 7528 6886 7540
rect 7745 7531 7803 7537
rect 7745 7528 7757 7531
rect 6880 7500 7757 7528
rect 6880 7488 6886 7500
rect 7745 7497 7757 7500
rect 7791 7497 7803 7531
rect 7745 7491 7803 7497
rect 8754 7488 8760 7540
rect 8812 7528 8818 7540
rect 8849 7531 8907 7537
rect 8849 7528 8861 7531
rect 8812 7500 8861 7528
rect 8812 7488 8818 7500
rect 8849 7497 8861 7500
rect 8895 7528 8907 7531
rect 9490 7528 9496 7540
rect 8895 7500 9496 7528
rect 8895 7497 8907 7500
rect 8849 7491 8907 7497
rect 9490 7488 9496 7500
rect 9548 7488 9554 7540
rect 9861 7531 9919 7537
rect 9861 7497 9873 7531
rect 9907 7528 9919 7531
rect 10042 7528 10048 7540
rect 9907 7500 10048 7528
rect 9907 7497 9919 7500
rect 9861 7491 9919 7497
rect 10042 7488 10048 7500
rect 10100 7488 10106 7540
rect 10873 7531 10931 7537
rect 10873 7497 10885 7531
rect 10919 7497 10931 7531
rect 10873 7491 10931 7497
rect 11425 7531 11483 7537
rect 11425 7497 11437 7531
rect 11471 7528 11483 7531
rect 11606 7528 11612 7540
rect 11471 7500 11612 7528
rect 11471 7497 11483 7500
rect 11425 7491 11483 7497
rect 7285 7463 7343 7469
rect 7285 7460 7297 7463
rect 2464 7432 4936 7460
rect 2464 7420 2470 7432
rect 658 7392 664 7404
rect 619 7364 664 7392
rect 658 7352 664 7364
rect 716 7352 722 7404
rect 2038 7352 2044 7404
rect 2096 7352 2102 7404
rect 2501 7395 2559 7401
rect 2501 7392 2513 7395
rect 2424 7364 2513 7392
rect 937 7327 995 7333
rect 937 7293 949 7327
rect 983 7324 995 7327
rect 1302 7324 1308 7336
rect 983 7296 1308 7324
rect 983 7293 995 7296
rect 937 7287 995 7293
rect 1302 7284 1308 7296
rect 1360 7284 1366 7336
rect 1946 7148 1952 7200
rect 2004 7188 2010 7200
rect 2424 7197 2452 7364
rect 2501 7361 2513 7364
rect 2547 7392 2559 7395
rect 2590 7392 2596 7404
rect 2547 7364 2596 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2590 7352 2596 7364
rect 2648 7352 2654 7404
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7392 3111 7395
rect 3142 7392 3148 7404
rect 3099 7364 3148 7392
rect 3099 7361 3111 7364
rect 3053 7355 3111 7361
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7392 3295 7395
rect 4062 7392 4068 7404
rect 3283 7364 4068 7392
rect 3283 7361 3295 7364
rect 3237 7355 3295 7361
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 4908 7401 4936 7432
rect 5092 7432 5948 7460
rect 6104 7432 7297 7460
rect 5092 7401 5120 7432
rect 5920 7404 5948 7432
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7361 4951 7395
rect 4893 7355 4951 7361
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7361 5135 7395
rect 5626 7392 5632 7404
rect 5587 7364 5632 7392
rect 5077 7355 5135 7361
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 5902 7352 5908 7404
rect 5960 7392 5966 7404
rect 7024 7401 7052 7432
rect 7285 7429 7297 7432
rect 7331 7429 7343 7463
rect 10060 7460 10088 7488
rect 10060 7432 10272 7460
rect 7285 7423 7343 7429
rect 6825 7395 6883 7401
rect 6825 7392 6837 7395
rect 5960 7364 6837 7392
rect 5960 7352 5966 7364
rect 6825 7361 6837 7364
rect 6871 7361 6883 7395
rect 6825 7355 6883 7361
rect 7009 7395 7067 7401
rect 7009 7361 7021 7395
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7361 7895 7395
rect 8754 7392 8760 7404
rect 8715 7364 8760 7392
rect 7837 7355 7895 7361
rect 3789 7327 3847 7333
rect 3789 7293 3801 7327
rect 3835 7324 3847 7327
rect 3970 7324 3976 7336
rect 3835 7296 3976 7324
rect 3835 7293 3847 7296
rect 3789 7287 3847 7293
rect 3970 7284 3976 7296
rect 4028 7284 4034 7336
rect 4706 7284 4712 7336
rect 4764 7324 4770 7336
rect 5718 7324 5724 7336
rect 4764 7296 5724 7324
rect 4764 7284 4770 7296
rect 5718 7284 5724 7296
rect 5776 7284 5782 7336
rect 5813 7327 5871 7333
rect 5813 7293 5825 7327
rect 5859 7324 5871 7327
rect 6089 7327 6147 7333
rect 6089 7324 6101 7327
rect 5859 7296 6101 7324
rect 5859 7293 5871 7296
rect 5813 7287 5871 7293
rect 6089 7293 6101 7296
rect 6135 7293 6147 7327
rect 6089 7287 6147 7293
rect 2958 7216 2964 7268
rect 3016 7256 3022 7268
rect 3513 7259 3571 7265
rect 3513 7256 3525 7259
rect 3016 7228 3525 7256
rect 3016 7216 3022 7228
rect 3513 7225 3525 7228
rect 3559 7256 3571 7259
rect 3878 7256 3884 7268
rect 3559 7228 3884 7256
rect 3559 7225 3571 7228
rect 3513 7219 3571 7225
rect 3878 7216 3884 7228
rect 3936 7216 3942 7268
rect 4893 7259 4951 7265
rect 4893 7225 4905 7259
rect 4939 7256 4951 7259
rect 5828 7256 5856 7287
rect 6454 7284 6460 7336
rect 6512 7324 6518 7336
rect 7852 7324 7880 7355
rect 8754 7352 8760 7364
rect 8812 7352 8818 7404
rect 9306 7392 9312 7404
rect 8864 7364 9312 7392
rect 6512 7296 7880 7324
rect 6512 7284 6518 7296
rect 7926 7284 7932 7336
rect 7984 7324 7990 7336
rect 8864 7324 8892 7364
rect 9306 7352 9312 7364
rect 9364 7392 9370 7404
rect 9493 7395 9551 7401
rect 9493 7392 9505 7395
rect 9364 7364 9505 7392
rect 9364 7352 9370 7364
rect 9493 7361 9505 7364
rect 9539 7361 9551 7395
rect 9493 7355 9551 7361
rect 9582 7352 9588 7404
rect 9640 7392 9646 7404
rect 9677 7395 9735 7401
rect 9677 7392 9689 7395
rect 9640 7364 9689 7392
rect 9640 7352 9646 7364
rect 9677 7361 9689 7364
rect 9723 7361 9735 7395
rect 9677 7355 9735 7361
rect 10042 7352 10048 7404
rect 10100 7390 10106 7404
rect 10244 7401 10272 7432
rect 10410 7420 10416 7472
rect 10468 7460 10474 7472
rect 10888 7460 10916 7491
rect 11606 7488 11612 7500
rect 11664 7488 11670 7540
rect 11698 7488 11704 7540
rect 11756 7488 11762 7540
rect 11882 7528 11888 7540
rect 11843 7500 11888 7528
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 13173 7531 13231 7537
rect 13173 7497 13185 7531
rect 13219 7528 13231 7531
rect 14182 7528 14188 7540
rect 13219 7500 14188 7528
rect 13219 7497 13231 7500
rect 13173 7491 13231 7497
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 14553 7531 14611 7537
rect 14553 7497 14565 7531
rect 14599 7528 14611 7531
rect 14734 7528 14740 7540
rect 14599 7500 14740 7528
rect 14599 7497 14611 7500
rect 14553 7491 14611 7497
rect 11149 7463 11207 7469
rect 11149 7460 11161 7463
rect 10468 7432 10824 7460
rect 10888 7432 11161 7460
rect 10468 7420 10474 7432
rect 10137 7395 10195 7401
rect 10137 7390 10149 7395
rect 10100 7362 10149 7390
rect 10100 7352 10106 7362
rect 10137 7361 10149 7362
rect 10183 7361 10195 7395
rect 10137 7355 10195 7361
rect 10229 7395 10287 7401
rect 10229 7361 10241 7395
rect 10275 7361 10287 7395
rect 10229 7355 10287 7361
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7361 10379 7395
rect 10594 7392 10600 7404
rect 10555 7364 10600 7392
rect 10321 7355 10379 7361
rect 7984 7296 8892 7324
rect 9033 7327 9091 7333
rect 7984 7284 7990 7296
rect 9033 7293 9045 7327
rect 9079 7324 9091 7327
rect 9214 7324 9220 7336
rect 9079 7296 9220 7324
rect 9079 7293 9091 7296
rect 9033 7287 9091 7293
rect 9214 7284 9220 7296
rect 9272 7284 9278 7336
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7324 9459 7327
rect 9766 7324 9772 7336
rect 9447 7296 9772 7324
rect 9447 7293 9459 7296
rect 9401 7287 9459 7293
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 4939 7228 5856 7256
rect 7469 7259 7527 7265
rect 4939 7225 4951 7228
rect 4893 7219 4951 7225
rect 7469 7225 7481 7259
rect 7515 7256 7527 7259
rect 7558 7256 7564 7268
rect 7515 7228 7564 7256
rect 7515 7225 7527 7228
rect 7469 7219 7527 7225
rect 7558 7216 7564 7228
rect 7616 7256 7622 7268
rect 10336 7256 10364 7355
rect 10594 7352 10600 7364
rect 10652 7352 10658 7404
rect 10796 7401 10824 7432
rect 11149 7429 11161 7432
rect 11195 7429 11207 7463
rect 11149 7423 11207 7429
rect 10781 7395 10839 7401
rect 10781 7361 10793 7395
rect 10827 7392 10839 7395
rect 10870 7392 10876 7404
rect 10827 7364 10876 7392
rect 10827 7361 10839 7364
rect 10781 7355 10839 7361
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 11330 7392 11336 7404
rect 11291 7364 11336 7392
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 11716 7401 11744 7488
rect 11977 7463 12035 7469
rect 11977 7429 11989 7463
rect 12023 7460 12035 7463
rect 12066 7460 12072 7472
rect 12023 7432 12072 7460
rect 12023 7429 12035 7432
rect 11977 7423 12035 7429
rect 12066 7420 12072 7432
rect 12124 7420 12130 7472
rect 14568 7460 14596 7491
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 14918 7528 14924 7540
rect 14879 7500 14924 7528
rect 14918 7488 14924 7500
rect 14976 7488 14982 7540
rect 15289 7531 15347 7537
rect 15289 7497 15301 7531
rect 15335 7528 15347 7531
rect 16114 7528 16120 7540
rect 15335 7500 16120 7528
rect 15335 7497 15347 7500
rect 15289 7491 15347 7497
rect 16114 7488 16120 7500
rect 16172 7488 16178 7540
rect 15102 7460 15108 7472
rect 14200 7432 14596 7460
rect 14844 7432 15108 7460
rect 11425 7395 11483 7401
rect 11425 7361 11437 7395
rect 11471 7361 11483 7395
rect 11425 7355 11483 7361
rect 11701 7395 11759 7401
rect 11701 7361 11713 7395
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 10505 7327 10563 7333
rect 10505 7293 10517 7327
rect 10551 7324 10563 7327
rect 11440 7324 11468 7355
rect 11790 7352 11796 7404
rect 11848 7392 11854 7404
rect 12802 7392 12808 7404
rect 11848 7364 11893 7392
rect 12763 7364 12808 7392
rect 11848 7352 11854 7364
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 14200 7401 14228 7432
rect 14093 7395 14151 7401
rect 14093 7361 14105 7395
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 14185 7395 14243 7401
rect 14185 7361 14197 7395
rect 14231 7361 14243 7395
rect 14185 7355 14243 7361
rect 12710 7324 12716 7336
rect 10551 7296 11468 7324
rect 12671 7296 12716 7324
rect 10551 7293 10563 7296
rect 10505 7287 10563 7293
rect 12710 7284 12716 7296
rect 12768 7284 12774 7336
rect 14108 7324 14136 7355
rect 14274 7352 14280 7404
rect 14332 7392 14338 7404
rect 14369 7395 14427 7401
rect 14369 7392 14381 7395
rect 14332 7364 14381 7392
rect 14332 7352 14338 7364
rect 14369 7361 14381 7364
rect 14415 7361 14427 7395
rect 14369 7355 14427 7361
rect 14458 7352 14464 7404
rect 14516 7392 14522 7404
rect 14844 7401 14872 7432
rect 15102 7420 15108 7432
rect 15160 7420 15166 7472
rect 15378 7420 15384 7472
rect 15436 7460 15442 7472
rect 15436 7432 15594 7460
rect 15436 7420 15442 7432
rect 14829 7395 14887 7401
rect 14516 7364 14561 7392
rect 14516 7352 14522 7364
rect 14829 7361 14841 7395
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 14918 7352 14924 7404
rect 14976 7392 14982 7404
rect 15013 7395 15071 7401
rect 15013 7392 15025 7395
rect 14976 7364 15025 7392
rect 14976 7352 14982 7364
rect 15013 7361 15025 7364
rect 15059 7361 15071 7395
rect 15013 7355 15071 7361
rect 15120 7324 15148 7420
rect 17034 7352 17040 7404
rect 17092 7392 17098 7404
rect 17092 7364 17137 7392
rect 17092 7352 17098 7364
rect 17310 7352 17316 7404
rect 17368 7392 17374 7404
rect 17405 7395 17463 7401
rect 17405 7392 17417 7395
rect 17368 7364 17417 7392
rect 17368 7352 17374 7364
rect 17405 7361 17417 7364
rect 17451 7361 17463 7395
rect 17405 7355 17463 7361
rect 16666 7324 16672 7336
rect 14108 7296 14872 7324
rect 15120 7296 16672 7324
rect 14844 7268 14872 7296
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 16761 7327 16819 7333
rect 16761 7293 16773 7327
rect 16807 7324 16819 7327
rect 18322 7324 18328 7336
rect 16807 7296 18328 7324
rect 16807 7293 16819 7296
rect 16761 7287 16819 7293
rect 18322 7284 18328 7296
rect 18380 7284 18386 7336
rect 11057 7259 11115 7265
rect 11057 7256 11069 7259
rect 7616 7228 8524 7256
rect 10336 7228 11069 7256
rect 7616 7216 7622 7228
rect 2409 7191 2467 7197
rect 2409 7188 2421 7191
rect 2004 7160 2421 7188
rect 2004 7148 2010 7160
rect 2409 7157 2421 7160
rect 2455 7157 2467 7191
rect 2409 7151 2467 7157
rect 3234 7148 3240 7200
rect 3292 7188 3298 7200
rect 3329 7191 3387 7197
rect 3329 7188 3341 7191
rect 3292 7160 3341 7188
rect 3292 7148 3298 7160
rect 3329 7157 3341 7160
rect 3375 7157 3387 7191
rect 5258 7188 5264 7200
rect 5219 7160 5264 7188
rect 3329 7151 3387 7157
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 5626 7148 5632 7200
rect 5684 7188 5690 7200
rect 7009 7191 7067 7197
rect 7009 7188 7021 7191
rect 5684 7160 7021 7188
rect 5684 7148 5690 7160
rect 7009 7157 7021 7160
rect 7055 7188 7067 7191
rect 8018 7188 8024 7200
rect 7055 7160 8024 7188
rect 7055 7157 7067 7160
rect 7009 7151 7067 7157
rect 8018 7148 8024 7160
rect 8076 7148 8082 7200
rect 8386 7188 8392 7200
rect 8347 7160 8392 7188
rect 8386 7148 8392 7160
rect 8444 7148 8450 7200
rect 8496 7188 8524 7228
rect 11057 7225 11069 7228
rect 11103 7256 11115 7259
rect 13722 7256 13728 7268
rect 11103 7228 13728 7256
rect 11103 7225 11115 7228
rect 11057 7219 11115 7225
rect 13722 7216 13728 7228
rect 13780 7216 13786 7268
rect 14826 7216 14832 7268
rect 14884 7216 14890 7268
rect 11330 7188 11336 7200
rect 8496 7160 11336 7188
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11609 7191 11667 7197
rect 11609 7157 11621 7191
rect 11655 7188 11667 7191
rect 12250 7188 12256 7200
rect 11655 7160 12256 7188
rect 11655 7157 11667 7160
rect 11609 7151 11667 7157
rect 12250 7148 12256 7160
rect 12308 7148 12314 7200
rect 14090 7188 14096 7200
rect 14051 7160 14096 7188
rect 14090 7148 14096 7160
rect 14148 7148 14154 7200
rect 14366 7148 14372 7200
rect 14424 7188 14430 7200
rect 15105 7191 15163 7197
rect 15105 7188 15117 7191
rect 14424 7160 15117 7188
rect 14424 7148 14430 7160
rect 15105 7157 15117 7160
rect 15151 7188 15163 7191
rect 15378 7188 15384 7200
rect 15151 7160 15384 7188
rect 15151 7157 15163 7160
rect 15105 7151 15163 7157
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 17218 7188 17224 7200
rect 17179 7160 17224 7188
rect 17218 7148 17224 7160
rect 17276 7148 17282 7200
rect 368 7098 18860 7120
rect 368 7046 3478 7098
rect 3530 7046 3542 7098
rect 3594 7046 3606 7098
rect 3658 7046 3670 7098
rect 3722 7046 3734 7098
rect 3786 7046 6578 7098
rect 6630 7046 6642 7098
rect 6694 7046 6706 7098
rect 6758 7046 6770 7098
rect 6822 7046 6834 7098
rect 6886 7046 9678 7098
rect 9730 7046 9742 7098
rect 9794 7046 9806 7098
rect 9858 7046 9870 7098
rect 9922 7046 9934 7098
rect 9986 7046 12778 7098
rect 12830 7046 12842 7098
rect 12894 7046 12906 7098
rect 12958 7046 12970 7098
rect 13022 7046 13034 7098
rect 13086 7046 15878 7098
rect 15930 7046 15942 7098
rect 15994 7046 16006 7098
rect 16058 7046 16070 7098
rect 16122 7046 16134 7098
rect 16186 7046 18860 7098
rect 368 7024 18860 7046
rect 2406 6984 2412 6996
rect 2367 6956 2412 6984
rect 2406 6944 2412 6956
rect 2464 6944 2470 6996
rect 5718 6944 5724 6996
rect 5776 6984 5782 6996
rect 6270 6984 6276 6996
rect 5776 6956 6276 6984
rect 5776 6944 5782 6956
rect 6270 6944 6276 6956
rect 6328 6944 6334 6996
rect 8754 6944 8760 6996
rect 8812 6984 8818 6996
rect 9033 6987 9091 6993
rect 9033 6984 9045 6987
rect 8812 6956 9045 6984
rect 8812 6944 8818 6956
rect 9033 6953 9045 6956
rect 9079 6953 9091 6987
rect 9033 6947 9091 6953
rect 9122 6944 9128 6996
rect 9180 6984 9186 6996
rect 9180 6956 9628 6984
rect 9180 6944 9186 6956
rect 1397 6919 1455 6925
rect 1397 6885 1409 6919
rect 1443 6916 1455 6919
rect 2869 6919 2927 6925
rect 1443 6888 2176 6916
rect 1443 6885 1455 6888
rect 1397 6879 1455 6885
rect 1213 6851 1271 6857
rect 1213 6817 1225 6851
rect 1259 6848 1271 6851
rect 2148 6848 2176 6888
rect 2869 6885 2881 6919
rect 2915 6916 2927 6919
rect 3050 6916 3056 6928
rect 2915 6888 3056 6916
rect 2915 6885 2927 6888
rect 2869 6879 2927 6885
rect 3050 6876 3056 6888
rect 3108 6876 3114 6928
rect 9600 6916 9628 6956
rect 10612 6956 10916 6984
rect 10410 6916 10416 6928
rect 6840 6888 7144 6916
rect 9600 6888 10416 6916
rect 3234 6848 3240 6860
rect 1259 6820 2084 6848
rect 2148 6820 3240 6848
rect 1259 6817 1271 6820
rect 1213 6811 1271 6817
rect 934 6780 940 6792
rect 895 6752 940 6780
rect 934 6740 940 6752
rect 992 6740 998 6792
rect 1486 6780 1492 6792
rect 1447 6752 1492 6780
rect 1486 6740 1492 6752
rect 1544 6740 1550 6792
rect 1946 6780 1952 6792
rect 1907 6752 1952 6780
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 2056 6789 2084 6820
rect 3234 6808 3240 6820
rect 3292 6808 3298 6860
rect 5353 6851 5411 6857
rect 3988 6820 4494 6848
rect 3988 6792 4016 6820
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6780 2099 6783
rect 2498 6780 2504 6792
rect 2087 6752 2360 6780
rect 2459 6752 2504 6780
rect 2087 6749 2099 6752
rect 2041 6743 2099 6749
rect 1302 6672 1308 6724
rect 1360 6712 1366 6724
rect 1360 6684 2268 6712
rect 1360 6672 1366 6684
rect 845 6647 903 6653
rect 845 6644 857 6647
rect 308 6616 857 6644
rect 308 6304 336 6616
rect 845 6613 857 6616
rect 891 6613 903 6647
rect 845 6607 903 6613
rect 1026 6604 1032 6656
rect 1084 6644 1090 6656
rect 2240 6653 2268 6684
rect 1213 6647 1271 6653
rect 1213 6644 1225 6647
rect 1084 6616 1225 6644
rect 1084 6604 1090 6616
rect 1213 6613 1225 6616
rect 1259 6613 1271 6647
rect 1213 6607 1271 6613
rect 2225 6647 2283 6653
rect 2225 6613 2237 6647
rect 2271 6613 2283 6647
rect 2332 6644 2360 6752
rect 2498 6740 2504 6752
rect 2556 6740 2562 6792
rect 2958 6780 2964 6792
rect 2919 6752 2964 6780
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6749 3387 6783
rect 3329 6743 3387 6749
rect 3344 6712 3372 6743
rect 3418 6740 3424 6792
rect 3476 6780 3482 6792
rect 3513 6783 3571 6789
rect 3513 6780 3525 6783
rect 3476 6752 3525 6780
rect 3476 6740 3482 6752
rect 3513 6749 3525 6752
rect 3559 6749 3571 6783
rect 3513 6743 3571 6749
rect 3602 6740 3608 6792
rect 3660 6780 3666 6792
rect 3660 6752 3705 6780
rect 3660 6740 3666 6752
rect 3786 6740 3792 6792
rect 3844 6780 3850 6792
rect 3970 6780 3976 6792
rect 3844 6752 3976 6780
rect 3844 6740 3850 6752
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 4466 6789 4494 6820
rect 5353 6817 5365 6851
rect 5399 6848 5411 6851
rect 5626 6848 5632 6860
rect 5399 6820 5632 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 5810 6808 5816 6860
rect 5868 6848 5874 6860
rect 6733 6851 6791 6857
rect 5868 6820 6684 6848
rect 5868 6808 5874 6820
rect 4249 6783 4307 6789
rect 4249 6780 4261 6783
rect 4212 6752 4261 6780
rect 4212 6740 4218 6752
rect 4249 6749 4261 6752
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 4433 6783 4494 6789
rect 4433 6749 4445 6783
rect 4479 6754 4494 6783
rect 4893 6783 4951 6789
rect 4479 6749 4491 6754
rect 4433 6743 4491 6749
rect 4893 6749 4905 6783
rect 4939 6780 4951 6783
rect 5258 6780 5264 6792
rect 4939 6752 5264 6780
rect 4939 6749 4951 6752
rect 4893 6743 4951 6749
rect 3697 6715 3755 6721
rect 3697 6712 3709 6715
rect 2746 6684 3280 6712
rect 3344 6684 3709 6712
rect 2746 6644 2774 6684
rect 3252 6653 3280 6684
rect 3697 6681 3709 6684
rect 3743 6681 3755 6715
rect 3697 6675 3755 6681
rect 3878 6672 3884 6724
rect 3936 6712 3942 6724
rect 4356 6712 4384 6743
rect 4908 6712 4936 6743
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 5445 6783 5503 6789
rect 5445 6749 5457 6783
rect 5491 6780 5503 6783
rect 5902 6780 5908 6792
rect 5491 6752 5908 6780
rect 5491 6749 5503 6752
rect 5445 6743 5503 6749
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 6656 6789 6684 6820
rect 6733 6817 6745 6851
rect 6779 6848 6791 6851
rect 6840 6848 6868 6888
rect 7006 6848 7012 6860
rect 6779 6820 6868 6848
rect 6967 6820 7012 6848
rect 6779 6817 6791 6820
rect 6733 6811 6791 6817
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 7116 6848 7144 6888
rect 10410 6876 10416 6888
rect 10468 6876 10474 6928
rect 7834 6848 7840 6860
rect 7116 6820 7840 6848
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6848 8171 6851
rect 8386 6848 8392 6860
rect 8159 6820 8392 6848
rect 8159 6817 8171 6820
rect 8113 6811 8171 6817
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 8478 6808 8484 6860
rect 8536 6848 8542 6860
rect 9585 6851 9643 6857
rect 9585 6848 9597 6851
rect 8536 6820 9597 6848
rect 8536 6808 8542 6820
rect 9585 6817 9597 6820
rect 9631 6848 9643 6851
rect 10612 6848 10640 6956
rect 10686 6876 10692 6928
rect 10744 6876 10750 6928
rect 10888 6925 10916 6956
rect 11054 6944 11060 6996
rect 11112 6984 11118 6996
rect 11241 6987 11299 6993
rect 11241 6984 11253 6987
rect 11112 6956 11253 6984
rect 11112 6944 11118 6956
rect 11241 6953 11253 6956
rect 11287 6953 11299 6987
rect 11241 6947 11299 6953
rect 13446 6944 13452 6996
rect 13504 6984 13510 6996
rect 16390 6984 16396 6996
rect 13504 6956 16396 6984
rect 13504 6944 13510 6956
rect 10873 6919 10931 6925
rect 10873 6885 10885 6919
rect 10919 6916 10931 6919
rect 12986 6916 12992 6928
rect 10919 6888 12992 6916
rect 10919 6885 10931 6888
rect 10873 6879 10931 6885
rect 12986 6876 12992 6888
rect 13044 6876 13050 6928
rect 9631 6820 10640 6848
rect 9631 6817 9643 6820
rect 9585 6811 9643 6817
rect 10702 6799 10730 6876
rect 13648 6857 13676 6956
rect 16390 6944 16396 6956
rect 16448 6944 16454 6996
rect 15194 6876 15200 6928
rect 15252 6916 15258 6928
rect 15427 6919 15485 6925
rect 15427 6916 15439 6919
rect 15252 6888 15439 6916
rect 15252 6876 15258 6888
rect 15427 6885 15439 6888
rect 15473 6885 15485 6919
rect 15427 6879 15485 6885
rect 13633 6851 13691 6857
rect 13633 6817 13645 6851
rect 13679 6817 13691 6851
rect 13633 6811 13691 6817
rect 13906 6808 13912 6860
rect 13964 6848 13970 6860
rect 14458 6848 14464 6860
rect 13964 6820 14464 6848
rect 13964 6808 13970 6820
rect 14458 6808 14464 6820
rect 14516 6848 14522 6860
rect 15010 6848 15016 6860
rect 14516 6820 15016 6848
rect 14516 6808 14522 6820
rect 15010 6808 15016 6820
rect 15068 6808 15074 6860
rect 16298 6848 16304 6860
rect 15856 6820 16304 6848
rect 10687 6793 10745 6799
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6780 6699 6783
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 6687 6752 7113 6780
rect 6687 6749 6699 6752
rect 6641 6743 6699 6749
rect 7101 6749 7113 6752
rect 7147 6749 7159 6783
rect 7653 6783 7711 6789
rect 7653 6780 7665 6783
rect 7101 6743 7159 6749
rect 7208 6752 7665 6780
rect 3936 6684 4200 6712
rect 4356 6684 4936 6712
rect 3936 6672 3942 6684
rect 2332 6616 2774 6644
rect 3237 6647 3295 6653
rect 2225 6607 2283 6613
rect 3237 6613 3249 6647
rect 3283 6613 3295 6647
rect 3237 6607 3295 6613
rect 3510 6604 3516 6656
rect 3568 6644 3574 6656
rect 4065 6647 4123 6653
rect 4065 6644 4077 6647
rect 3568 6616 4077 6644
rect 3568 6604 3574 6616
rect 4065 6613 4077 6616
rect 4111 6613 4123 6647
rect 4172 6644 4200 6684
rect 5534 6672 5540 6724
rect 5592 6712 5598 6724
rect 7208 6712 7236 6752
rect 7653 6749 7665 6752
rect 7699 6749 7711 6783
rect 7653 6743 7711 6749
rect 7374 6712 7380 6724
rect 5592 6684 7236 6712
rect 7335 6684 7380 6712
rect 5592 6672 5598 6684
rect 7374 6672 7380 6684
rect 7432 6672 7438 6724
rect 7558 6712 7564 6724
rect 7519 6684 7564 6712
rect 7558 6672 7564 6684
rect 7616 6672 7622 6724
rect 7668 6712 7696 6743
rect 8018 6740 8024 6792
rect 8076 6780 8082 6792
rect 8205 6783 8263 6789
rect 8205 6780 8217 6783
rect 8076 6752 8217 6780
rect 8076 6740 8082 6752
rect 8205 6749 8217 6752
rect 8251 6749 8263 6783
rect 10226 6780 10232 6792
rect 8205 6743 8263 6749
rect 8864 6752 10232 6780
rect 8864 6712 8892 6752
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 10687 6759 10699 6793
rect 10733 6759 10745 6793
rect 10687 6753 10745 6759
rect 10781 6785 10839 6791
rect 10781 6751 10793 6785
rect 10827 6780 10839 6785
rect 10870 6780 10876 6792
rect 10827 6752 10876 6780
rect 10827 6751 10839 6752
rect 10781 6745 10839 6751
rect 10870 6740 10876 6752
rect 10928 6740 10934 6792
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 12253 6783 12311 6789
rect 12253 6780 12265 6783
rect 11112 6752 12265 6780
rect 11112 6740 11118 6752
rect 12253 6749 12265 6752
rect 12299 6780 12311 6783
rect 12618 6780 12624 6792
rect 12299 6752 12624 6780
rect 12299 6749 12311 6752
rect 12253 6743 12311 6749
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 13998 6780 14004 6792
rect 13959 6752 14004 6780
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 15856 6789 15884 6820
rect 16298 6808 16304 6820
rect 16356 6808 16362 6860
rect 16761 6851 16819 6857
rect 16761 6817 16773 6851
rect 16807 6848 16819 6851
rect 17218 6848 17224 6860
rect 16807 6820 17224 6848
rect 16807 6817 16819 6820
rect 16761 6811 16819 6817
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 17770 6808 17776 6860
rect 17828 6848 17834 6860
rect 18187 6851 18245 6857
rect 18187 6848 18199 6851
rect 17828 6820 18199 6848
rect 17828 6808 17834 6820
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6780 16267 6783
rect 16255 6752 16344 6780
rect 16255 6749 16267 6752
rect 16209 6743 16267 6749
rect 7668 6684 8892 6712
rect 8938 6672 8944 6724
rect 8996 6712 9002 6724
rect 10410 6712 10416 6724
rect 8996 6684 10416 6712
rect 8996 6672 9002 6684
rect 10410 6672 10416 6684
rect 10468 6672 10474 6724
rect 10577 6715 10635 6721
rect 10577 6681 10589 6715
rect 10623 6712 10635 6715
rect 11330 6712 11336 6724
rect 10623 6684 11336 6712
rect 10623 6681 10635 6684
rect 10577 6675 10635 6681
rect 11330 6672 11336 6684
rect 11388 6672 11394 6724
rect 14366 6672 14372 6724
rect 14424 6672 14430 6724
rect 4709 6647 4767 6653
rect 4709 6644 4721 6647
rect 4172 6616 4721 6644
rect 4065 6607 4123 6613
rect 4709 6613 4721 6616
rect 4755 6613 4767 6647
rect 4709 6607 4767 6613
rect 4798 6604 4804 6656
rect 4856 6644 4862 6656
rect 5169 6647 5227 6653
rect 5169 6644 5181 6647
rect 4856 6616 5181 6644
rect 4856 6604 4862 6616
rect 5169 6613 5181 6616
rect 5215 6613 5227 6647
rect 5169 6607 5227 6613
rect 5718 6604 5724 6656
rect 5776 6644 5782 6656
rect 5813 6647 5871 6653
rect 5813 6644 5825 6647
rect 5776 6616 5825 6644
rect 5776 6604 5782 6616
rect 5813 6613 5825 6616
rect 5859 6613 5871 6647
rect 5813 6607 5871 6613
rect 7193 6647 7251 6653
rect 7193 6613 7205 6647
rect 7239 6644 7251 6647
rect 7466 6644 7472 6656
rect 7239 6616 7472 6644
rect 7239 6613 7251 6616
rect 7193 6607 7251 6613
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 7653 6647 7711 6653
rect 7653 6613 7665 6647
rect 7699 6644 7711 6647
rect 7745 6647 7803 6653
rect 7745 6644 7757 6647
rect 7699 6616 7757 6644
rect 7699 6613 7711 6616
rect 7653 6607 7711 6613
rect 7745 6613 7757 6616
rect 7791 6613 7803 6647
rect 7745 6607 7803 6613
rect 8389 6647 8447 6653
rect 8389 6613 8401 6647
rect 8435 6644 8447 6647
rect 8570 6644 8576 6656
rect 8435 6616 8576 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 9398 6644 9404 6656
rect 9359 6616 9404 6644
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 9490 6604 9496 6656
rect 9548 6644 9554 6656
rect 10689 6647 10747 6653
rect 9548 6616 9593 6644
rect 9548 6604 9554 6616
rect 10689 6613 10701 6647
rect 10735 6644 10747 6647
rect 10778 6644 10784 6656
rect 10735 6616 10784 6644
rect 10735 6613 10747 6616
rect 10689 6607 10747 6613
rect 10778 6604 10784 6616
rect 10836 6604 10842 6656
rect 12253 6647 12311 6653
rect 12253 6613 12265 6647
rect 12299 6644 12311 6647
rect 12802 6644 12808 6656
rect 12299 6616 12808 6644
rect 12299 6613 12311 6616
rect 12253 6607 12311 6613
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 13354 6644 13360 6656
rect 13315 6616 13360 6644
rect 13354 6604 13360 6616
rect 13412 6644 13418 6656
rect 14384 6644 14412 6672
rect 15746 6644 15752 6656
rect 13412 6616 14412 6644
rect 15707 6616 15752 6644
rect 13412 6604 13418 6616
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 16206 6644 16212 6656
rect 16167 6616 16212 6644
rect 16206 6604 16212 6616
rect 16264 6604 16270 6656
rect 16316 6644 16344 6752
rect 16390 6740 16396 6792
rect 16448 6780 16454 6792
rect 16448 6752 16493 6780
rect 16448 6740 16454 6752
rect 17126 6672 17132 6724
rect 17184 6672 17190 6724
rect 16666 6644 16672 6656
rect 16316 6616 16672 6644
rect 16666 6604 16672 6616
rect 16724 6644 16730 6656
rect 17880 6644 17908 6820
rect 18187 6817 18199 6820
rect 18233 6817 18245 6851
rect 18187 6811 18245 6817
rect 16724 6616 17908 6644
rect 16724 6604 16730 6616
rect 368 6554 18860 6576
rect 368 6502 5028 6554
rect 5080 6502 5092 6554
rect 5144 6502 5156 6554
rect 5208 6502 5220 6554
rect 5272 6502 5284 6554
rect 5336 6502 8128 6554
rect 8180 6502 8192 6554
rect 8244 6502 8256 6554
rect 8308 6502 8320 6554
rect 8372 6502 8384 6554
rect 8436 6502 11228 6554
rect 11280 6502 11292 6554
rect 11344 6502 11356 6554
rect 11408 6502 11420 6554
rect 11472 6502 11484 6554
rect 11536 6502 14328 6554
rect 14380 6502 14392 6554
rect 14444 6502 14456 6554
rect 14508 6502 14520 6554
rect 14572 6502 14584 6554
rect 14636 6502 17428 6554
rect 17480 6502 17492 6554
rect 17544 6502 17556 6554
rect 17608 6502 17620 6554
rect 17672 6502 17684 6554
rect 17736 6502 18860 6554
rect 368 6480 18860 6502
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 3510 6440 3516 6452
rect 2556 6412 3516 6440
rect 2556 6400 2562 6412
rect 3510 6400 3516 6412
rect 3568 6400 3574 6452
rect 5718 6440 5724 6452
rect 5679 6412 5724 6440
rect 5718 6400 5724 6412
rect 5776 6400 5782 6452
rect 5902 6440 5908 6452
rect 5863 6412 5908 6440
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 6273 6443 6331 6449
rect 6273 6409 6285 6443
rect 6319 6440 6331 6443
rect 6733 6443 6791 6449
rect 6733 6440 6745 6443
rect 6319 6412 6745 6440
rect 6319 6409 6331 6412
rect 6273 6403 6331 6409
rect 6733 6409 6745 6412
rect 6779 6409 6791 6443
rect 6733 6403 6791 6409
rect 7006 6400 7012 6452
rect 7064 6440 7070 6452
rect 7101 6443 7159 6449
rect 7101 6440 7113 6443
rect 7064 6412 7113 6440
rect 7064 6400 7070 6412
rect 7101 6409 7113 6412
rect 7147 6409 7159 6443
rect 7558 6440 7564 6452
rect 7101 6403 7159 6409
rect 7208 6412 7564 6440
rect 2038 6332 2044 6384
rect 2096 6372 2102 6384
rect 2096 6344 2728 6372
rect 2096 6332 2102 6344
rect 661 6307 719 6313
rect 661 6304 673 6307
rect 308 6276 673 6304
rect 661 6273 673 6276
rect 707 6273 719 6307
rect 1026 6304 1032 6316
rect 987 6276 1032 6304
rect 661 6267 719 6273
rect 1026 6264 1032 6276
rect 1084 6264 1090 6316
rect 2700 6245 2728 6344
rect 3050 6332 3056 6384
rect 3108 6372 3114 6384
rect 5629 6375 5687 6381
rect 3108 6344 3188 6372
rect 3108 6332 3114 6344
rect 3160 6313 3188 6344
rect 5629 6341 5641 6375
rect 5675 6372 5687 6375
rect 7208 6372 7236 6412
rect 7558 6400 7564 6412
rect 7616 6400 7622 6452
rect 8849 6443 8907 6449
rect 8849 6409 8861 6443
rect 8895 6440 8907 6443
rect 10042 6440 10048 6452
rect 8895 6412 10048 6440
rect 8895 6409 8907 6412
rect 8849 6403 8907 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10689 6443 10747 6449
rect 10689 6409 10701 6443
rect 10735 6440 10747 6443
rect 10778 6440 10784 6452
rect 10735 6412 10784 6440
rect 10735 6409 10747 6412
rect 10689 6403 10747 6409
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 11793 6443 11851 6449
rect 11793 6409 11805 6443
rect 11839 6440 11851 6443
rect 12437 6443 12495 6449
rect 12437 6440 12449 6443
rect 11839 6412 12449 6440
rect 11839 6409 11851 6412
rect 11793 6403 11851 6409
rect 12437 6409 12449 6412
rect 12483 6409 12495 6443
rect 12802 6440 12808 6452
rect 12763 6412 12808 6440
rect 12437 6403 12495 6409
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 12897 6443 12955 6449
rect 12897 6409 12909 6443
rect 12943 6440 12955 6443
rect 13814 6440 13820 6452
rect 12943 6412 13820 6440
rect 12943 6409 12955 6412
rect 12897 6403 12955 6409
rect 8478 6372 8484 6384
rect 5675 6344 7236 6372
rect 7300 6344 8484 6372
rect 5675 6341 5687 6344
rect 5629 6335 5687 6341
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6273 3203 6307
rect 5534 6304 5540 6316
rect 5495 6276 5540 6304
rect 3145 6267 3203 6273
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 5810 6304 5816 6316
rect 5771 6276 5816 6304
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 5994 6264 6000 6316
rect 6052 6304 6058 6316
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 6052 6276 6377 6304
rect 6052 6264 6058 6276
rect 6365 6273 6377 6276
rect 6411 6304 6423 6307
rect 6411 6276 7236 6304
rect 6411 6273 6423 6276
rect 6365 6267 6423 6273
rect 2685 6239 2743 6245
rect 2685 6205 2697 6239
rect 2731 6236 2743 6239
rect 2774 6236 2780 6248
rect 2731 6208 2780 6236
rect 2731 6205 2743 6208
rect 2685 6199 2743 6205
rect 2774 6196 2780 6208
rect 2832 6196 2838 6248
rect 3050 6236 3056 6248
rect 3011 6208 3056 6236
rect 3050 6196 3056 6208
rect 3108 6196 3114 6248
rect 6270 6196 6276 6248
rect 6328 6236 6334 6248
rect 7208 6245 7236 6276
rect 7300 6245 7328 6344
rect 8478 6332 8484 6344
rect 8536 6332 8542 6384
rect 8757 6375 8815 6381
rect 8757 6341 8769 6375
rect 8803 6372 8815 6375
rect 9125 6375 9183 6381
rect 9125 6372 9137 6375
rect 8803 6344 9137 6372
rect 8803 6341 8815 6344
rect 8757 6335 8815 6341
rect 9125 6341 9137 6344
rect 9171 6341 9183 6375
rect 9125 6335 9183 6341
rect 9582 6332 9588 6384
rect 9640 6372 9646 6384
rect 9640 6344 11284 6372
rect 9640 6332 9646 6344
rect 7466 6264 7472 6316
rect 7524 6304 7530 6316
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 7524 6276 8677 6304
rect 7524 6264 7530 6276
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 8938 6304 8944 6316
rect 8899 6276 8944 6304
rect 8665 6267 8723 6273
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 9033 6307 9091 6313
rect 9033 6273 9045 6307
rect 9079 6273 9091 6307
rect 11146 6304 11152 6316
rect 9033 6267 9091 6273
rect 9140 6276 11152 6304
rect 6549 6239 6607 6245
rect 6549 6236 6561 6239
rect 6328 6208 6561 6236
rect 6328 6196 6334 6208
rect 6549 6205 6561 6208
rect 6595 6205 6607 6239
rect 6549 6199 6607 6205
rect 7193 6239 7251 6245
rect 7193 6205 7205 6239
rect 7239 6205 7251 6239
rect 7193 6199 7251 6205
rect 7285 6239 7343 6245
rect 7285 6205 7297 6239
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 2455 6171 2513 6177
rect 2455 6137 2467 6171
rect 2501 6168 2513 6171
rect 3142 6168 3148 6180
rect 2501 6140 3148 6168
rect 2501 6137 2513 6140
rect 2455 6131 2513 6137
rect 3142 6128 3148 6140
rect 3200 6168 3206 6180
rect 3602 6168 3608 6180
rect 3200 6140 3608 6168
rect 3200 6128 3206 6140
rect 3602 6128 3608 6140
rect 3660 6128 3666 6180
rect 2866 6100 2872 6112
rect 2827 6072 2872 6100
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 4157 6103 4215 6109
rect 4157 6100 4169 6103
rect 4120 6072 4169 6100
rect 4120 6060 4126 6072
rect 4157 6069 4169 6072
rect 4203 6069 4215 6103
rect 6564 6100 6592 6199
rect 7208 6168 7236 6199
rect 7374 6196 7380 6248
rect 7432 6236 7438 6248
rect 8478 6236 8484 6248
rect 7432 6208 8484 6236
rect 7432 6196 7438 6208
rect 8478 6196 8484 6208
rect 8536 6236 8542 6248
rect 9048 6236 9076 6267
rect 8536 6208 9076 6236
rect 8536 6196 8542 6208
rect 7926 6168 7932 6180
rect 7208 6140 7932 6168
rect 7926 6128 7932 6140
rect 7984 6128 7990 6180
rect 8018 6128 8024 6180
rect 8076 6168 8082 6180
rect 9140 6168 9168 6276
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 11256 6304 11284 6344
rect 11885 6310 11943 6313
rect 11885 6307 12020 6310
rect 11885 6304 11897 6307
rect 11256 6276 11897 6304
rect 11885 6273 11897 6276
rect 11931 6304 12020 6307
rect 11931 6282 12434 6304
rect 11931 6273 11943 6282
rect 11992 6276 12434 6282
rect 11885 6267 11943 6273
rect 11054 6236 11060 6248
rect 11015 6208 11060 6236
rect 11054 6196 11060 6208
rect 11112 6196 11118 6248
rect 12069 6239 12127 6245
rect 12069 6236 12081 6239
rect 11164 6208 12081 6236
rect 8076 6140 9168 6168
rect 8076 6128 8082 6140
rect 9214 6128 9220 6180
rect 9272 6168 9278 6180
rect 11164 6168 11192 6208
rect 12069 6205 12081 6208
rect 12115 6236 12127 6239
rect 12158 6236 12164 6248
rect 12115 6208 12164 6236
rect 12115 6205 12127 6208
rect 12069 6199 12127 6205
rect 12158 6196 12164 6208
rect 12216 6196 12222 6248
rect 9272 6140 11192 6168
rect 11333 6171 11391 6177
rect 9272 6128 9278 6140
rect 11333 6137 11345 6171
rect 11379 6168 11391 6171
rect 11514 6168 11520 6180
rect 11379 6140 11520 6168
rect 11379 6137 11391 6140
rect 11333 6131 11391 6137
rect 11514 6128 11520 6140
rect 11572 6128 11578 6180
rect 12406 6168 12434 6276
rect 12986 6236 12992 6248
rect 12947 6208 12992 6236
rect 12986 6196 12992 6208
rect 13044 6196 13050 6248
rect 13096 6168 13124 6412
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 13998 6440 14004 6452
rect 13959 6412 14004 6440
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 14553 6443 14611 6449
rect 14553 6409 14565 6443
rect 14599 6440 14611 6443
rect 14826 6440 14832 6452
rect 14599 6412 14832 6440
rect 14599 6409 14611 6412
rect 14553 6403 14611 6409
rect 14826 6400 14832 6412
rect 14884 6440 14890 6452
rect 14884 6412 15332 6440
rect 14884 6400 14890 6412
rect 14182 6332 14188 6384
rect 14240 6372 14246 6384
rect 14921 6375 14979 6381
rect 14921 6372 14933 6375
rect 14240 6344 14933 6372
rect 14240 6332 14246 6344
rect 13909 6307 13967 6313
rect 13909 6273 13921 6307
rect 13955 6273 13967 6307
rect 14090 6304 14096 6316
rect 14051 6276 14096 6304
rect 13909 6267 13967 6273
rect 13924 6236 13952 6267
rect 14090 6264 14096 6276
rect 14148 6264 14154 6316
rect 14384 6313 14412 6344
rect 14921 6341 14933 6344
rect 14967 6341 14979 6375
rect 15304 6372 15332 6412
rect 16206 6400 16212 6452
rect 16264 6440 16270 6452
rect 16577 6443 16635 6449
rect 16577 6440 16589 6443
rect 16264 6412 16589 6440
rect 16264 6400 16270 6412
rect 16577 6409 16589 6412
rect 16623 6409 16635 6443
rect 16577 6403 16635 6409
rect 16669 6443 16727 6449
rect 16669 6409 16681 6443
rect 16715 6440 16727 6443
rect 16850 6440 16856 6452
rect 16715 6412 16856 6440
rect 16715 6409 16727 6412
rect 16669 6403 16727 6409
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 17037 6443 17095 6449
rect 17037 6409 17049 6443
rect 17083 6440 17095 6443
rect 17589 6443 17647 6449
rect 17589 6440 17601 6443
rect 17083 6412 17601 6440
rect 17083 6409 17095 6412
rect 17037 6403 17095 6409
rect 17589 6409 17601 6412
rect 17635 6409 17647 6443
rect 17589 6403 17647 6409
rect 17681 6443 17739 6449
rect 17681 6409 17693 6443
rect 17727 6440 17739 6443
rect 17770 6440 17776 6452
rect 17727 6412 17776 6440
rect 17727 6409 17739 6412
rect 17681 6403 17739 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 18322 6440 18328 6452
rect 18283 6412 18328 6440
rect 18322 6400 18328 6412
rect 18380 6400 18386 6452
rect 16298 6372 16304 6384
rect 15304 6344 16304 6372
rect 14921 6335 14979 6341
rect 16298 6332 16304 6344
rect 16356 6332 16362 6384
rect 14369 6307 14427 6313
rect 14369 6273 14381 6307
rect 14415 6273 14427 6307
rect 14369 6267 14427 6273
rect 14645 6307 14703 6313
rect 14645 6273 14657 6307
rect 14691 6304 14703 6307
rect 14734 6304 14740 6316
rect 14691 6276 14740 6304
rect 14691 6273 14703 6276
rect 14645 6267 14703 6273
rect 14734 6264 14740 6276
rect 14792 6264 14798 6316
rect 15013 6307 15071 6313
rect 15013 6273 15025 6307
rect 15059 6304 15071 6307
rect 15194 6304 15200 6316
rect 15059 6276 15200 6304
rect 15059 6273 15071 6276
rect 15013 6267 15071 6273
rect 15194 6264 15200 6276
rect 15252 6264 15258 6316
rect 15565 6307 15623 6313
rect 15565 6304 15577 6307
rect 15304 6276 15577 6304
rect 14185 6239 14243 6245
rect 14185 6236 14197 6239
rect 13924 6208 14197 6236
rect 14185 6205 14197 6208
rect 14231 6205 14243 6239
rect 14185 6199 14243 6205
rect 14918 6196 14924 6248
rect 14976 6236 14982 6248
rect 15304 6236 15332 6276
rect 15565 6273 15577 6276
rect 15611 6273 15623 6307
rect 15565 6267 15623 6273
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6304 18291 6307
rect 18506 6304 18512 6316
rect 18279 6276 18512 6304
rect 18279 6273 18291 6276
rect 18233 6267 18291 6273
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 14976 6208 15332 6236
rect 14976 6196 14982 6208
rect 15470 6196 15476 6248
rect 15528 6236 15534 6248
rect 15657 6239 15715 6245
rect 15657 6236 15669 6239
rect 15528 6208 15669 6236
rect 15528 6196 15534 6208
rect 15657 6205 15669 6208
rect 15703 6205 15715 6239
rect 15657 6199 15715 6205
rect 15746 6196 15752 6248
rect 15804 6236 15810 6248
rect 16393 6239 16451 6245
rect 16393 6236 16405 6239
rect 15804 6208 16405 6236
rect 15804 6196 15810 6208
rect 16393 6205 16405 6208
rect 16439 6205 16451 6239
rect 17862 6236 17868 6248
rect 17823 6208 17868 6236
rect 16393 6199 16451 6205
rect 17862 6196 17868 6208
rect 17920 6196 17926 6248
rect 12406 6140 13124 6168
rect 14458 6128 14464 6180
rect 14516 6168 14522 6180
rect 15197 6171 15255 6177
rect 15197 6168 15209 6171
rect 14516 6140 15209 6168
rect 14516 6128 14522 6140
rect 15197 6137 15209 6140
rect 15243 6137 15255 6171
rect 15197 6131 15255 6137
rect 17221 6171 17279 6177
rect 17221 6137 17233 6171
rect 17267 6168 17279 6171
rect 17310 6168 17316 6180
rect 17267 6140 17316 6168
rect 17267 6137 17279 6140
rect 17221 6131 17279 6137
rect 17310 6128 17316 6140
rect 17368 6128 17374 6180
rect 9232 6100 9260 6128
rect 6564 6072 9260 6100
rect 4157 6063 4215 6069
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 11425 6103 11483 6109
rect 11425 6100 11437 6103
rect 11112 6072 11437 6100
rect 11112 6060 11118 6072
rect 11425 6069 11437 6072
rect 11471 6069 11483 6103
rect 11425 6063 11483 6069
rect 15746 6060 15752 6112
rect 15804 6100 15810 6112
rect 16117 6103 16175 6109
rect 16117 6100 16129 6103
rect 15804 6072 16129 6100
rect 15804 6060 15810 6072
rect 16117 6069 16129 6072
rect 16163 6069 16175 6103
rect 16117 6063 16175 6069
rect 368 6010 18860 6032
rect 368 5958 3478 6010
rect 3530 5958 3542 6010
rect 3594 5958 3606 6010
rect 3658 5958 3670 6010
rect 3722 5958 3734 6010
rect 3786 5958 6578 6010
rect 6630 5958 6642 6010
rect 6694 5958 6706 6010
rect 6758 5958 6770 6010
rect 6822 5958 6834 6010
rect 6886 5958 9678 6010
rect 9730 5958 9742 6010
rect 9794 5958 9806 6010
rect 9858 5958 9870 6010
rect 9922 5958 9934 6010
rect 9986 5958 12778 6010
rect 12830 5958 12842 6010
rect 12894 5958 12906 6010
rect 12958 5958 12970 6010
rect 13022 5958 13034 6010
rect 13086 5958 15878 6010
rect 15930 5958 15942 6010
rect 15994 5958 16006 6010
rect 16058 5958 16070 6010
rect 16122 5958 16134 6010
rect 16186 5958 18860 6010
rect 368 5936 18860 5958
rect 2304 5899 2362 5905
rect 2304 5865 2316 5899
rect 2350 5896 2362 5899
rect 2866 5896 2872 5908
rect 2350 5868 2872 5896
rect 2350 5865 2362 5868
rect 2304 5859 2362 5865
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 3050 5856 3056 5908
rect 3108 5896 3114 5908
rect 3789 5899 3847 5905
rect 3789 5896 3801 5899
rect 3108 5868 3801 5896
rect 3108 5856 3114 5868
rect 3789 5865 3801 5868
rect 3835 5896 3847 5899
rect 3878 5896 3884 5908
rect 3835 5868 3884 5896
rect 3835 5865 3847 5868
rect 3789 5859 3847 5865
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 5626 5856 5632 5908
rect 5684 5896 5690 5908
rect 6549 5899 6607 5905
rect 6549 5896 6561 5899
rect 5684 5868 6561 5896
rect 5684 5856 5690 5868
rect 6549 5865 6561 5868
rect 6595 5896 6607 5899
rect 7190 5896 7196 5908
rect 6595 5868 7196 5896
rect 6595 5865 6607 5868
rect 6549 5859 6607 5865
rect 7190 5856 7196 5868
rect 7248 5896 7254 5908
rect 7742 5896 7748 5908
rect 7248 5868 7748 5896
rect 7248 5856 7254 5868
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 10781 5899 10839 5905
rect 10781 5865 10793 5899
rect 10827 5896 10839 5899
rect 15654 5896 15660 5908
rect 10827 5868 15660 5896
rect 10827 5865 10839 5868
rect 10781 5859 10839 5865
rect 5810 5788 5816 5840
rect 5868 5828 5874 5840
rect 5997 5831 6055 5837
rect 5997 5828 6009 5831
rect 5868 5800 6009 5828
rect 5868 5788 5874 5800
rect 5997 5797 6009 5800
rect 6043 5797 6055 5831
rect 5997 5791 6055 5797
rect 6871 5831 6929 5837
rect 6871 5797 6883 5831
rect 6917 5828 6929 5831
rect 7374 5828 7380 5840
rect 6917 5800 7380 5828
rect 6917 5797 6929 5800
rect 6871 5791 6929 5797
rect 7374 5788 7380 5800
rect 7432 5788 7438 5840
rect 934 5720 940 5772
rect 992 5760 998 5772
rect 2041 5763 2099 5769
rect 2041 5760 2053 5763
rect 992 5732 2053 5760
rect 992 5720 998 5732
rect 2041 5729 2053 5732
rect 2087 5760 2099 5763
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 2087 5732 4261 5760
rect 2087 5729 2099 5732
rect 2041 5723 2099 5729
rect 4249 5729 4261 5732
rect 4295 5760 4307 5763
rect 6454 5760 6460 5772
rect 4295 5732 6460 5760
rect 4295 5729 4307 5732
rect 4249 5723 4307 5729
rect 6454 5720 6460 5732
rect 6512 5720 6518 5772
rect 8849 5763 8907 5769
rect 8849 5760 8861 5763
rect 6656 5732 8861 5760
rect 2774 5584 2780 5636
rect 2832 5584 2838 5636
rect 4525 5627 4583 5633
rect 2792 5556 2820 5584
rect 3528 5556 3556 5610
rect 4525 5593 4537 5627
rect 4571 5624 4583 5627
rect 4798 5624 4804 5636
rect 4571 5596 4804 5624
rect 4571 5593 4583 5596
rect 4525 5587 4583 5593
rect 4798 5584 4804 5596
rect 4856 5584 4862 5636
rect 6472 5624 6500 5720
rect 6656 5701 6684 5732
rect 8849 5729 8861 5732
rect 8895 5760 8907 5763
rect 9674 5760 9680 5772
rect 8895 5732 9680 5760
rect 8895 5729 8907 5732
rect 8849 5723 8907 5729
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5661 6699 5695
rect 6641 5655 6699 5661
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5692 8355 5695
rect 8570 5692 8576 5704
rect 8343 5664 8576 5692
rect 8343 5661 8355 5664
rect 8297 5655 8355 5661
rect 8570 5652 8576 5664
rect 8628 5652 8634 5704
rect 8665 5695 8723 5701
rect 8665 5661 8677 5695
rect 8711 5661 8723 5695
rect 8665 5655 8723 5661
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5692 10655 5695
rect 10796 5692 10824 5859
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 17862 5896 17868 5908
rect 16316 5868 17868 5896
rect 12618 5788 12624 5840
rect 12676 5828 12682 5840
rect 12989 5831 13047 5837
rect 12989 5828 13001 5831
rect 12676 5800 13001 5828
rect 12676 5788 12682 5800
rect 12989 5797 13001 5800
rect 13035 5797 13047 5831
rect 15470 5828 15476 5840
rect 15431 5800 15476 5828
rect 12989 5791 13047 5797
rect 15470 5788 15476 5800
rect 15528 5788 15534 5840
rect 16316 5837 16344 5868
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 15565 5831 15623 5837
rect 15565 5797 15577 5831
rect 15611 5828 15623 5831
rect 16301 5831 16359 5837
rect 16301 5828 16313 5831
rect 15611 5800 16313 5828
rect 15611 5797 15623 5800
rect 15565 5791 15623 5797
rect 16301 5797 16313 5800
rect 16347 5797 16359 5831
rect 16301 5791 16359 5797
rect 16390 5788 16396 5840
rect 16448 5828 16454 5840
rect 16448 5800 16528 5828
rect 16448 5788 16454 5800
rect 11241 5763 11299 5769
rect 11241 5729 11253 5763
rect 11287 5760 11299 5763
rect 13446 5760 13452 5772
rect 11287 5732 13452 5760
rect 11287 5729 11299 5732
rect 11241 5723 11299 5729
rect 13446 5720 13452 5732
rect 13504 5720 13510 5772
rect 14737 5763 14795 5769
rect 14737 5729 14749 5763
rect 14783 5760 14795 5763
rect 14826 5760 14832 5772
rect 14783 5732 14832 5760
rect 14783 5729 14795 5732
rect 14737 5723 14795 5729
rect 14826 5720 14832 5732
rect 14884 5720 14890 5772
rect 16500 5769 16528 5800
rect 15197 5763 15255 5769
rect 15197 5729 15209 5763
rect 15243 5760 15255 5763
rect 16492 5763 16550 5769
rect 15243 5732 16436 5760
rect 15243 5729 15255 5732
rect 15197 5723 15255 5729
rect 10643 5664 10824 5692
rect 13817 5695 13875 5701
rect 10643 5661 10655 5664
rect 10597 5655 10655 5661
rect 13817 5661 13829 5695
rect 13863 5692 13875 5695
rect 14458 5692 14464 5704
rect 13863 5664 14136 5692
rect 14419 5664 14464 5692
rect 13863 5661 13875 5664
rect 13817 5655 13875 5661
rect 4062 5556 4068 5568
rect 2792 5528 4068 5556
rect 4062 5516 4068 5528
rect 4120 5556 4126 5568
rect 4157 5559 4215 5565
rect 4157 5556 4169 5559
rect 4120 5528 4169 5556
rect 4120 5516 4126 5528
rect 4157 5525 4169 5528
rect 4203 5556 4215 5559
rect 5534 5556 5540 5568
rect 4203 5528 5540 5556
rect 4203 5525 4215 5528
rect 4157 5519 4215 5525
rect 5534 5516 5540 5528
rect 5592 5556 5598 5568
rect 5736 5556 5764 5610
rect 6472 5596 7236 5624
rect 6273 5559 6331 5565
rect 6273 5556 6285 5559
rect 5592 5528 6285 5556
rect 5592 5516 5598 5528
rect 6273 5525 6285 5528
rect 6319 5556 6331 5559
rect 7006 5556 7012 5568
rect 6319 5528 7012 5556
rect 6319 5525 6331 5528
rect 6273 5519 6331 5525
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 7208 5556 7236 5596
rect 7926 5584 7932 5636
rect 7984 5584 7990 5636
rect 8680 5556 8708 5655
rect 11514 5624 11520 5636
rect 11475 5596 11520 5624
rect 11514 5584 11520 5596
rect 11572 5584 11578 5636
rect 12250 5584 12256 5636
rect 12308 5584 12314 5636
rect 7208 5528 8708 5556
rect 10410 5516 10416 5568
rect 10468 5556 10474 5568
rect 10965 5559 11023 5565
rect 10965 5556 10977 5559
rect 10468 5528 10977 5556
rect 10468 5516 10474 5528
rect 10965 5525 10977 5528
rect 11011 5525 11023 5559
rect 10965 5519 11023 5525
rect 13170 5516 13176 5568
rect 13228 5556 13234 5568
rect 14108 5565 14136 5664
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 16408 5701 16436 5732
rect 16492 5729 16504 5763
rect 16538 5729 16550 5763
rect 16492 5723 16550 5729
rect 15105 5695 15163 5701
rect 15105 5692 15117 5695
rect 15028 5664 15117 5692
rect 14553 5627 14611 5633
rect 14553 5593 14565 5627
rect 14599 5624 14611 5627
rect 14734 5624 14740 5636
rect 14599 5596 14740 5624
rect 14599 5593 14611 5596
rect 14553 5587 14611 5593
rect 14734 5584 14740 5596
rect 14792 5624 14798 5636
rect 15028 5624 15056 5664
rect 15105 5661 15117 5664
rect 15151 5661 15163 5695
rect 15105 5655 15163 5661
rect 16393 5695 16451 5701
rect 16393 5661 16405 5695
rect 16439 5661 16451 5695
rect 16393 5655 16451 5661
rect 16117 5627 16175 5633
rect 16117 5624 16129 5627
rect 14792 5596 16129 5624
rect 14792 5584 14798 5596
rect 16117 5593 16129 5596
rect 16163 5624 16175 5627
rect 16206 5624 16212 5636
rect 16163 5596 16212 5624
rect 16163 5593 16175 5596
rect 16117 5587 16175 5593
rect 16206 5584 16212 5596
rect 16264 5584 16270 5636
rect 16408 5624 16436 5655
rect 16758 5624 16764 5636
rect 16408 5596 16620 5624
rect 16719 5596 16764 5624
rect 16592 5568 16620 5596
rect 16758 5584 16764 5596
rect 16816 5584 16822 5636
rect 16850 5584 16856 5636
rect 16908 5624 16914 5636
rect 17218 5624 17224 5636
rect 16908 5596 17224 5624
rect 16908 5584 16914 5596
rect 17218 5584 17224 5596
rect 17276 5584 17282 5636
rect 13633 5559 13691 5565
rect 13633 5556 13645 5559
rect 13228 5528 13645 5556
rect 13228 5516 13234 5528
rect 13633 5525 13645 5528
rect 13679 5525 13691 5559
rect 13633 5519 13691 5525
rect 14093 5559 14151 5565
rect 14093 5525 14105 5559
rect 14139 5525 14151 5559
rect 14093 5519 14151 5525
rect 14826 5516 14832 5568
rect 14884 5556 14890 5568
rect 15565 5559 15623 5565
rect 15565 5556 15577 5559
rect 14884 5528 15577 5556
rect 14884 5516 14890 5528
rect 15565 5525 15577 5528
rect 15611 5525 15623 5559
rect 15746 5556 15752 5568
rect 15707 5528 15752 5556
rect 15565 5519 15623 5525
rect 15746 5516 15752 5528
rect 15804 5516 15810 5568
rect 15838 5516 15844 5568
rect 15896 5556 15902 5568
rect 16393 5559 16451 5565
rect 16393 5556 16405 5559
rect 15896 5528 16405 5556
rect 15896 5516 15902 5528
rect 16393 5525 16405 5528
rect 16439 5525 16451 5559
rect 16393 5519 16451 5525
rect 16574 5516 16580 5568
rect 16632 5516 16638 5568
rect 16666 5516 16672 5568
rect 16724 5556 16730 5568
rect 18233 5559 18291 5565
rect 18233 5556 18245 5559
rect 16724 5528 18245 5556
rect 16724 5516 16730 5528
rect 18233 5525 18245 5528
rect 18279 5525 18291 5559
rect 18233 5519 18291 5525
rect 368 5466 18860 5488
rect 368 5414 5028 5466
rect 5080 5414 5092 5466
rect 5144 5414 5156 5466
rect 5208 5414 5220 5466
rect 5272 5414 5284 5466
rect 5336 5414 8128 5466
rect 8180 5414 8192 5466
rect 8244 5414 8256 5466
rect 8308 5414 8320 5466
rect 8372 5414 8384 5466
rect 8436 5414 11228 5466
rect 11280 5414 11292 5466
rect 11344 5414 11356 5466
rect 11408 5414 11420 5466
rect 11472 5414 11484 5466
rect 11536 5414 14328 5466
rect 14380 5414 14392 5466
rect 14444 5414 14456 5466
rect 14508 5414 14520 5466
rect 14572 5414 14584 5466
rect 14636 5414 17428 5466
rect 17480 5414 17492 5466
rect 17544 5414 17556 5466
rect 17608 5414 17620 5466
rect 17672 5414 17684 5466
rect 17736 5414 18860 5466
rect 368 5392 18860 5414
rect 4062 5352 4068 5364
rect 4023 5324 4068 5352
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 5534 5352 5540 5364
rect 5495 5324 5540 5352
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 7834 5312 7840 5364
rect 7892 5352 7898 5364
rect 8665 5355 8723 5361
rect 8665 5352 8677 5355
rect 7892 5324 8677 5352
rect 7892 5312 7898 5324
rect 8665 5321 8677 5324
rect 8711 5321 8723 5355
rect 9398 5352 9404 5364
rect 9359 5324 9404 5352
rect 8665 5315 8723 5321
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 10686 5352 10692 5364
rect 10152 5324 10692 5352
rect 7012 5296 7064 5302
rect 10152 5296 10180 5324
rect 10686 5312 10692 5324
rect 10744 5352 10750 5364
rect 13354 5352 13360 5364
rect 10744 5324 11836 5352
rect 10744 5312 10750 5324
rect 7190 5284 7196 5296
rect 7064 5256 7196 5284
rect 7190 5244 7196 5256
rect 7248 5284 7254 5296
rect 7926 5284 7932 5296
rect 7248 5256 7932 5284
rect 7248 5244 7254 5256
rect 7926 5244 7932 5256
rect 7984 5244 7990 5296
rect 9674 5284 9680 5296
rect 8588 5256 9076 5284
rect 9635 5256 9680 5284
rect 7012 5238 7064 5244
rect 5626 5216 5632 5228
rect 5587 5188 5632 5216
rect 5626 5176 5632 5188
rect 5684 5176 5690 5228
rect 8478 5176 8484 5228
rect 8536 5216 8542 5228
rect 8588 5225 8616 5256
rect 9048 5225 9076 5256
rect 9674 5244 9680 5256
rect 9732 5244 9738 5296
rect 9861 5287 9919 5293
rect 9861 5253 9873 5287
rect 9907 5284 9919 5287
rect 10134 5284 10140 5296
rect 9907 5256 10140 5284
rect 9907 5253 9919 5256
rect 9861 5247 9919 5253
rect 10134 5244 10140 5256
rect 10192 5244 10198 5296
rect 8573 5219 8631 5225
rect 8573 5216 8585 5219
rect 8536 5188 8585 5216
rect 8536 5176 8542 5188
rect 8573 5185 8585 5188
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 9033 5219 9091 5225
rect 9033 5185 9045 5219
rect 9079 5185 9091 5219
rect 9033 5179 9091 5185
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 5997 5151 6055 5157
rect 5997 5148 6009 5151
rect 5960 5120 6009 5148
rect 5960 5108 5966 5120
rect 5997 5117 6009 5120
rect 6043 5117 6055 5151
rect 8772 5148 8800 5179
rect 10410 5176 10416 5228
rect 10468 5176 10474 5228
rect 11808 5225 11836 5324
rect 12728 5324 13360 5352
rect 12250 5244 12256 5296
rect 12308 5284 12314 5296
rect 12728 5293 12756 5324
rect 13354 5312 13360 5324
rect 13412 5352 13418 5364
rect 14645 5355 14703 5361
rect 13412 5324 13676 5352
rect 13412 5312 13418 5324
rect 12713 5287 12771 5293
rect 12713 5284 12725 5287
rect 12308 5256 12725 5284
rect 12308 5244 12314 5256
rect 12713 5253 12725 5256
rect 12759 5253 12771 5287
rect 13446 5284 13452 5296
rect 12713 5247 12771 5253
rect 12912 5256 13452 5284
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5216 11851 5219
rect 12618 5216 12624 5228
rect 11839 5188 12624 5216
rect 11839 5185 11851 5188
rect 11793 5179 11851 5185
rect 12618 5176 12624 5188
rect 12676 5176 12682 5228
rect 12912 5225 12940 5256
rect 13446 5244 13452 5256
rect 13504 5244 13510 5296
rect 13648 5270 13676 5324
rect 14645 5321 14657 5355
rect 14691 5352 14703 5355
rect 14734 5352 14740 5364
rect 14691 5324 14740 5352
rect 14691 5321 14703 5324
rect 14645 5315 14703 5321
rect 14734 5312 14740 5324
rect 14792 5312 14798 5364
rect 16298 5352 16304 5364
rect 16259 5324 16304 5352
rect 16298 5312 16304 5324
rect 16356 5312 16362 5364
rect 16574 5312 16580 5364
rect 16632 5352 16638 5364
rect 16632 5324 17080 5352
rect 16632 5312 16638 5324
rect 15764 5256 16712 5284
rect 15764 5225 15792 5256
rect 16684 5228 16712 5256
rect 12897 5219 12955 5225
rect 12897 5185 12909 5219
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 15749 5219 15807 5225
rect 15749 5185 15761 5219
rect 15795 5185 15807 5219
rect 16206 5216 16212 5228
rect 16167 5188 16212 5216
rect 15749 5179 15807 5185
rect 16206 5176 16212 5188
rect 16264 5176 16270 5228
rect 16666 5216 16672 5228
rect 16627 5188 16672 5216
rect 16666 5176 16672 5188
rect 16724 5176 16730 5228
rect 17052 5225 17080 5324
rect 17037 5219 17095 5225
rect 17037 5185 17049 5219
rect 17083 5185 17095 5219
rect 17037 5179 17095 5185
rect 18233 5219 18291 5225
rect 18233 5185 18245 5219
rect 18279 5216 18291 5219
rect 18506 5216 18512 5228
rect 18279 5188 18512 5216
rect 18279 5185 18291 5188
rect 18233 5179 18291 5185
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 8938 5148 8944 5160
rect 8772 5120 8944 5148
rect 5997 5111 6055 5117
rect 8938 5108 8944 5120
rect 8996 5108 9002 5160
rect 10045 5151 10103 5157
rect 10045 5117 10057 5151
rect 10091 5148 10103 5151
rect 10318 5148 10324 5160
rect 10091 5120 10324 5148
rect 10091 5117 10103 5120
rect 10045 5111 10103 5117
rect 10318 5108 10324 5120
rect 10376 5108 10382 5160
rect 11517 5151 11575 5157
rect 11517 5117 11529 5151
rect 11563 5148 11575 5151
rect 13170 5148 13176 5160
rect 11563 5120 12434 5148
rect 13131 5120 13176 5148
rect 11563 5117 11575 5120
rect 11517 5111 11575 5117
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 7377 5015 7435 5021
rect 7377 5012 7389 5015
rect 6972 4984 7389 5012
rect 6972 4972 6978 4984
rect 7377 4981 7389 4984
rect 7423 4981 7435 5015
rect 12406 5012 12434 5120
rect 13170 5108 13176 5120
rect 13228 5108 13234 5160
rect 15838 5148 15844 5160
rect 15799 5120 15844 5148
rect 15838 5108 15844 5120
rect 15896 5108 15902 5160
rect 16117 5151 16175 5157
rect 16117 5117 16129 5151
rect 16163 5148 16175 5151
rect 16758 5148 16764 5160
rect 16163 5120 16764 5148
rect 16163 5117 16175 5120
rect 16117 5111 16175 5117
rect 16758 5108 16764 5120
rect 16816 5108 16822 5160
rect 18138 5012 18144 5024
rect 12406 4984 18144 5012
rect 7377 4975 7435 4981
rect 18138 4972 18144 4984
rect 18196 4972 18202 5024
rect 18322 5012 18328 5024
rect 18283 4984 18328 5012
rect 18322 4972 18328 4984
rect 18380 4972 18386 5024
rect 368 4922 18860 4944
rect 368 4870 3478 4922
rect 3530 4870 3542 4922
rect 3594 4870 3606 4922
rect 3658 4870 3670 4922
rect 3722 4870 3734 4922
rect 3786 4870 6578 4922
rect 6630 4870 6642 4922
rect 6694 4870 6706 4922
rect 6758 4870 6770 4922
rect 6822 4870 6834 4922
rect 6886 4870 9678 4922
rect 9730 4870 9742 4922
rect 9794 4870 9806 4922
rect 9858 4870 9870 4922
rect 9922 4870 9934 4922
rect 9986 4870 12778 4922
rect 12830 4870 12842 4922
rect 12894 4870 12906 4922
rect 12958 4870 12970 4922
rect 13022 4870 13034 4922
rect 13086 4870 15878 4922
rect 15930 4870 15942 4922
rect 15994 4870 16006 4922
rect 16058 4870 16070 4922
rect 16122 4870 16134 4922
rect 16186 4870 18860 4922
rect 368 4848 18860 4870
rect 4893 4811 4951 4817
rect 4893 4808 4905 4811
rect 1228 4780 4905 4808
rect 934 4672 940 4684
rect 895 4644 940 4672
rect 934 4632 940 4644
rect 992 4632 998 4684
rect 1228 4681 1256 4780
rect 4893 4777 4905 4780
rect 4939 4777 4951 4811
rect 5902 4808 5908 4820
rect 5863 4780 5908 4808
rect 4893 4771 4951 4777
rect 5902 4768 5908 4780
rect 5960 4768 5966 4820
rect 7926 4808 7932 4820
rect 7839 4780 7932 4808
rect 7926 4768 7932 4780
rect 7984 4808 7990 4820
rect 9398 4808 9404 4820
rect 7984 4780 9404 4808
rect 7984 4768 7990 4780
rect 9398 4768 9404 4780
rect 9456 4808 9462 4820
rect 12731 4811 12789 4817
rect 9456 4780 9674 4808
rect 9456 4768 9462 4780
rect 3881 4743 3939 4749
rect 3881 4709 3893 4743
rect 3927 4740 3939 4743
rect 4062 4740 4068 4752
rect 3927 4712 4068 4740
rect 3927 4709 3939 4712
rect 3881 4703 3939 4709
rect 4062 4700 4068 4712
rect 4120 4700 4126 4752
rect 5626 4740 5632 4752
rect 4448 4712 5632 4740
rect 1213 4675 1271 4681
rect 1213 4641 1225 4675
rect 1259 4641 1271 4675
rect 2130 4672 2136 4684
rect 2043 4644 2136 4672
rect 1213 4635 1271 4641
rect 2130 4632 2136 4644
rect 2188 4672 2194 4684
rect 4448 4672 4476 4712
rect 5626 4700 5632 4712
rect 5684 4700 5690 4752
rect 6457 4743 6515 4749
rect 6457 4709 6469 4743
rect 6503 4709 6515 4743
rect 6457 4703 6515 4709
rect 2188 4644 4476 4672
rect 4709 4675 4767 4681
rect 2188 4632 2194 4644
rect 4709 4641 4721 4675
rect 4755 4672 4767 4675
rect 4755 4644 5212 4672
rect 4755 4641 4767 4644
rect 4709 4635 4767 4641
rect 1302 4604 1308 4616
rect 1263 4576 1308 4604
rect 1302 4564 1308 4576
rect 1360 4564 1366 4616
rect 4062 4564 4068 4616
rect 4120 4604 4126 4616
rect 4525 4607 4583 4613
rect 4525 4604 4537 4607
rect 4120 4576 4537 4604
rect 4120 4564 4126 4576
rect 4525 4573 4537 4576
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4573 4951 4607
rect 4893 4567 4951 4573
rect 2409 4539 2467 4545
rect 2409 4505 2421 4539
rect 2455 4505 2467 4539
rect 3878 4536 3884 4548
rect 3634 4508 3884 4536
rect 2409 4499 2467 4505
rect 2424 4468 2452 4499
rect 3878 4496 3884 4508
rect 3936 4496 3942 4548
rect 2774 4468 2780 4480
rect 2424 4440 2780 4468
rect 2774 4428 2780 4440
rect 2832 4428 2838 4480
rect 3970 4428 3976 4480
rect 4028 4468 4034 4480
rect 4065 4471 4123 4477
rect 4065 4468 4077 4471
rect 4028 4440 4077 4468
rect 4028 4428 4034 4440
rect 4065 4437 4077 4440
rect 4111 4437 4123 4471
rect 4430 4468 4436 4480
rect 4391 4440 4436 4468
rect 4065 4431 4123 4437
rect 4430 4428 4436 4440
rect 4488 4428 4494 4480
rect 4798 4428 4804 4480
rect 4856 4468 4862 4480
rect 4908 4468 4936 4567
rect 4982 4564 4988 4616
rect 5040 4604 5046 4616
rect 5040 4576 5085 4604
rect 5040 4564 5046 4576
rect 5184 4545 5212 4644
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4604 6147 4607
rect 6472 4604 6500 4703
rect 6914 4672 6920 4684
rect 6875 4644 6920 4672
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 7101 4675 7159 4681
rect 7101 4641 7113 4675
rect 7147 4672 7159 4675
rect 7926 4672 7932 4684
rect 7147 4644 7932 4672
rect 7147 4641 7159 4644
rect 7101 4635 7159 4641
rect 7116 4604 7144 4635
rect 7926 4632 7932 4644
rect 7984 4632 7990 4684
rect 9646 4672 9674 4780
rect 12731 4777 12743 4811
rect 12777 4808 12789 4811
rect 18322 4808 18328 4820
rect 12777 4780 18328 4808
rect 12777 4777 12789 4780
rect 12731 4771 12789 4777
rect 18322 4768 18328 4780
rect 18380 4768 18386 4820
rect 9953 4675 10011 4681
rect 9953 4672 9965 4675
rect 9646 4644 9965 4672
rect 9953 4641 9965 4644
rect 9999 4672 10011 4675
rect 10410 4672 10416 4684
rect 9999 4644 10416 4672
rect 9999 4641 10011 4644
rect 9953 4635 10011 4641
rect 10410 4632 10416 4644
rect 10468 4672 10474 4684
rect 11057 4675 11115 4681
rect 11057 4672 11069 4675
rect 10468 4644 11069 4672
rect 10468 4632 10474 4644
rect 11057 4641 11069 4644
rect 11103 4672 11115 4675
rect 12250 4672 12256 4684
rect 11103 4644 12256 4672
rect 11103 4641 11115 4644
rect 11057 4635 11115 4641
rect 12250 4632 12256 4644
rect 12308 4632 12314 4684
rect 12618 4632 12624 4684
rect 12676 4672 12682 4684
rect 14090 4672 14096 4684
rect 12676 4644 14096 4672
rect 12676 4632 12682 4644
rect 14090 4632 14096 4644
rect 14148 4632 14154 4684
rect 6135 4576 6500 4604
rect 6564 4576 7144 4604
rect 12989 4607 13047 4613
rect 6135 4573 6147 4576
rect 6089 4567 6147 4573
rect 5169 4539 5227 4545
rect 5169 4505 5181 4539
rect 5215 4536 5227 4539
rect 6564 4536 6592 4576
rect 12989 4573 13001 4607
rect 13035 4604 13047 4607
rect 13262 4604 13268 4616
rect 13035 4576 13268 4604
rect 13035 4573 13047 4576
rect 12989 4567 13047 4573
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 13354 4564 13360 4616
rect 13412 4604 13418 4616
rect 13909 4607 13967 4613
rect 13909 4604 13921 4607
rect 13412 4576 13921 4604
rect 13412 4564 13418 4576
rect 13909 4573 13921 4576
rect 13955 4573 13967 4607
rect 13909 4567 13967 4573
rect 17865 4607 17923 4613
rect 17865 4573 17877 4607
rect 17911 4604 17923 4607
rect 17954 4604 17960 4616
rect 17911 4576 17960 4604
rect 17911 4573 17923 4576
rect 17865 4567 17923 4573
rect 17954 4564 17960 4576
rect 18012 4564 18018 4616
rect 18230 4604 18236 4616
rect 18191 4576 18236 4604
rect 18230 4564 18236 4576
rect 18288 4564 18294 4616
rect 5215 4508 6592 4536
rect 6825 4539 6883 4545
rect 5215 4505 5227 4508
rect 5169 4499 5227 4505
rect 6825 4505 6837 4539
rect 6871 4536 6883 4539
rect 7098 4536 7104 4548
rect 6871 4508 7104 4536
rect 6871 4505 6883 4508
rect 6825 4499 6883 4505
rect 7098 4496 7104 4508
rect 7156 4496 7162 4548
rect 12250 4496 12256 4548
rect 12308 4496 12314 4548
rect 13446 4496 13452 4548
rect 13504 4536 13510 4548
rect 13725 4539 13783 4545
rect 13725 4536 13737 4539
rect 13504 4508 13737 4536
rect 13504 4496 13510 4508
rect 13725 4505 13737 4508
rect 13771 4505 13783 4539
rect 13725 4499 13783 4505
rect 14182 4496 14188 4548
rect 14240 4536 14246 4548
rect 14338 4539 14396 4545
rect 14338 4536 14350 4539
rect 14240 4508 14350 4536
rect 14240 4496 14246 4508
rect 14338 4505 14350 4508
rect 14384 4505 14396 4539
rect 14338 4499 14396 4505
rect 15746 4496 15752 4548
rect 15804 4536 15810 4548
rect 16850 4536 16856 4548
rect 15804 4508 16856 4536
rect 15804 4496 15810 4508
rect 16224 4480 16252 4508
rect 16850 4496 16856 4508
rect 16908 4496 16914 4548
rect 6914 4468 6920 4480
rect 4856 4440 6920 4468
rect 4856 4428 4862 4440
rect 6914 4428 6920 4440
rect 6972 4428 6978 4480
rect 11241 4471 11299 4477
rect 11241 4437 11253 4471
rect 11287 4468 11299 4471
rect 12710 4468 12716 4480
rect 11287 4440 12716 4468
rect 11287 4437 11299 4440
rect 11241 4431 11299 4437
rect 12710 4428 12716 4440
rect 12768 4428 12774 4480
rect 15470 4468 15476 4480
rect 15431 4440 15476 4468
rect 15470 4428 15476 4440
rect 15528 4428 15534 4480
rect 16206 4468 16212 4480
rect 16167 4440 16212 4468
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 16439 4471 16497 4477
rect 16439 4437 16451 4471
rect 16485 4468 16497 4471
rect 17862 4468 17868 4480
rect 16485 4440 17868 4468
rect 16485 4437 16497 4440
rect 16439 4431 16497 4437
rect 17862 4428 17868 4440
rect 17920 4428 17926 4480
rect 368 4378 18860 4400
rect 368 4326 5028 4378
rect 5080 4326 5092 4378
rect 5144 4326 5156 4378
rect 5208 4326 5220 4378
rect 5272 4326 5284 4378
rect 5336 4326 8128 4378
rect 8180 4326 8192 4378
rect 8244 4326 8256 4378
rect 8308 4326 8320 4378
rect 8372 4326 8384 4378
rect 8436 4326 11228 4378
rect 11280 4326 11292 4378
rect 11344 4326 11356 4378
rect 11408 4326 11420 4378
rect 11472 4326 11484 4378
rect 11536 4326 14328 4378
rect 14380 4326 14392 4378
rect 14444 4326 14456 4378
rect 14508 4326 14520 4378
rect 14572 4326 14584 4378
rect 14636 4326 17428 4378
rect 17480 4326 17492 4378
rect 17544 4326 17556 4378
rect 17608 4326 17620 4378
rect 17672 4326 17684 4378
rect 17736 4326 18860 4378
rect 368 4304 18860 4326
rect 2774 4224 2780 4276
rect 2832 4264 2838 4276
rect 2961 4267 3019 4273
rect 2961 4264 2973 4267
rect 2832 4236 2973 4264
rect 2832 4224 2838 4236
rect 2961 4233 2973 4236
rect 3007 4233 3019 4267
rect 2961 4227 3019 4233
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 5537 4267 5595 4273
rect 5537 4264 5549 4267
rect 4488 4236 5549 4264
rect 4488 4224 4494 4236
rect 5537 4233 5549 4236
rect 5583 4233 5595 4267
rect 7098 4264 7104 4276
rect 7059 4236 7104 4264
rect 5537 4227 5595 4233
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 10686 4264 10692 4276
rect 7208 4236 10548 4264
rect 10647 4236 10692 4264
rect 934 4196 940 4208
rect 895 4168 940 4196
rect 934 4156 940 4168
rect 992 4156 998 4208
rect 3970 4196 3976 4208
rect 3160 4168 3976 4196
rect 2774 4128 2780 4140
rect 2070 4100 2780 4128
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 3160 4137 3188 4168
rect 3970 4156 3976 4168
rect 4028 4156 4034 4208
rect 6733 4199 6791 4205
rect 6733 4165 6745 4199
rect 6779 4196 6791 4199
rect 7208 4196 7236 4236
rect 6779 4168 7236 4196
rect 6779 4165 6791 4168
rect 6733 4159 6791 4165
rect 9398 4156 9404 4208
rect 9456 4156 9462 4208
rect 10520 4196 10548 4236
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 14182 4264 14188 4276
rect 11072 4236 14188 4264
rect 11072 4196 11100 4236
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 17954 4224 17960 4276
rect 18012 4264 18018 4276
rect 18325 4267 18383 4273
rect 18325 4264 18337 4267
rect 18012 4236 18337 4264
rect 18012 4224 18018 4236
rect 18325 4233 18337 4236
rect 18371 4233 18383 4267
rect 18325 4227 18383 4233
rect 10520 4168 11100 4196
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4097 3939 4131
rect 4062 4128 4068 4140
rect 4023 4100 4068 4128
rect 3881 4091 3939 4097
rect 201 4063 259 4069
rect 201 4029 213 4063
rect 247 4060 259 4063
rect 661 4063 719 4069
rect 661 4060 673 4063
rect 247 4032 673 4060
rect 247 4029 259 4032
rect 201 4023 259 4029
rect 661 4029 673 4032
rect 707 4029 719 4063
rect 661 4023 719 4029
rect 1302 4020 1308 4072
rect 1360 4060 1366 4072
rect 2409 4063 2467 4069
rect 2409 4060 2421 4063
rect 1360 4032 2421 4060
rect 1360 4020 1366 4032
rect 2409 4029 2421 4032
rect 2455 4060 2467 4063
rect 3896 4060 3924 4091
rect 4062 4088 4068 4100
rect 4120 4128 4126 4140
rect 4709 4131 4767 4137
rect 4709 4128 4721 4131
rect 4120 4100 4721 4128
rect 4120 4088 4126 4100
rect 4709 4097 4721 4100
rect 4755 4128 4767 4131
rect 4890 4128 4896 4140
rect 4755 4100 4896 4128
rect 4755 4097 4767 4100
rect 4709 4091 4767 4097
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5905 4131 5963 4137
rect 5905 4097 5917 4131
rect 5951 4128 5963 4131
rect 6086 4128 6092 4140
rect 5951 4100 6092 4128
rect 5951 4097 5963 4100
rect 5905 4091 5963 4097
rect 6086 4088 6092 4100
rect 6144 4088 6150 4140
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 7285 4131 7343 4137
rect 7285 4128 7297 4131
rect 6972 4100 7297 4128
rect 6972 4088 6978 4100
rect 7285 4097 7297 4100
rect 7331 4097 7343 4131
rect 7742 4128 7748 4140
rect 7703 4100 7748 4128
rect 7285 4091 7343 4097
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 8021 4131 8079 4137
rect 8021 4097 8033 4131
rect 8067 4128 8079 4131
rect 8067 4100 8524 4128
rect 8067 4097 8079 4100
rect 8021 4091 8079 4097
rect 4798 4060 4804 4072
rect 2455 4032 3924 4060
rect 4759 4032 4804 4060
rect 2455 4029 2467 4032
rect 2409 4023 2467 4029
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 5997 4063 6055 4069
rect 5997 4060 6009 4063
rect 5092 4032 6009 4060
rect 5092 4001 5120 4032
rect 5997 4029 6009 4032
rect 6043 4029 6055 4063
rect 5997 4023 6055 4029
rect 6181 4063 6239 4069
rect 6181 4029 6193 4063
rect 6227 4060 6239 4063
rect 6454 4060 6460 4072
rect 6227 4032 6460 4060
rect 6227 4029 6239 4032
rect 6181 4023 6239 4029
rect 6454 4020 6460 4032
rect 6512 4020 6518 4072
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4060 6699 4063
rect 7193 4063 7251 4069
rect 7193 4060 7205 4063
rect 6687 4032 7205 4060
rect 6687 4029 6699 4032
rect 6641 4023 6699 4029
rect 7193 4029 7205 4032
rect 7239 4029 7251 4063
rect 7193 4023 7251 4029
rect 8202 4020 8208 4072
rect 8260 4060 8266 4072
rect 8389 4063 8447 4069
rect 8389 4060 8401 4063
rect 8260 4032 8401 4060
rect 8260 4020 8266 4032
rect 8389 4029 8401 4032
rect 8435 4029 8447 4063
rect 8496 4060 8524 4100
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 11072 4137 11100 4168
rect 12250 4156 12256 4208
rect 12308 4196 12314 4208
rect 12308 4168 13202 4196
rect 12308 4156 12314 4168
rect 10597 4131 10655 4137
rect 10597 4128 10609 4131
rect 10100 4100 10609 4128
rect 10100 4088 10106 4100
rect 10597 4097 10609 4100
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 11057 4131 11115 4137
rect 11057 4097 11069 4131
rect 11103 4097 11115 4131
rect 11238 4128 11244 4140
rect 11199 4100 11244 4128
rect 11057 4091 11115 4097
rect 11238 4088 11244 4100
rect 11296 4088 11302 4140
rect 14200 4128 14228 4224
rect 15470 4128 15476 4140
rect 14200 4100 14964 4128
rect 15431 4100 15476 4128
rect 10686 4060 10692 4072
rect 8496 4032 10692 4060
rect 8389 4023 8447 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 10873 4063 10931 4069
rect 10873 4029 10885 4063
rect 10919 4060 10931 4063
rect 11149 4063 11207 4069
rect 11149 4060 11161 4063
rect 10919 4032 11161 4060
rect 10919 4029 10931 4032
rect 10873 4023 10931 4029
rect 11149 4029 11161 4032
rect 11195 4029 11207 4063
rect 11149 4023 11207 4029
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4029 12495 4063
rect 12710 4060 12716 4072
rect 12671 4032 12716 4060
rect 12437 4023 12495 4029
rect 5077 3995 5135 4001
rect 5077 3961 5089 3995
rect 5123 3961 5135 3995
rect 5077 3955 5135 3961
rect 12452 3936 12480 4023
rect 12710 4020 12716 4032
rect 12768 4020 12774 4072
rect 13354 4020 13360 4072
rect 13412 4060 13418 4072
rect 14461 4063 14519 4069
rect 14461 4060 14473 4063
rect 13412 4032 14473 4060
rect 13412 4020 13418 4032
rect 14461 4029 14473 4032
rect 14507 4029 14519 4063
rect 14461 4023 14519 4029
rect 2593 3927 2651 3933
rect 2593 3893 2605 3927
rect 2639 3924 2651 3927
rect 2774 3924 2780 3936
rect 2639 3896 2780 3924
rect 2639 3893 2651 3896
rect 2593 3887 2651 3893
rect 2774 3884 2780 3896
rect 2832 3884 2838 3936
rect 4065 3927 4123 3933
rect 4065 3893 4077 3927
rect 4111 3924 4123 3927
rect 6362 3924 6368 3936
rect 4111 3896 6368 3924
rect 4111 3893 4123 3896
rect 4065 3887 4123 3893
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 7837 3927 7895 3933
rect 7837 3893 7849 3927
rect 7883 3924 7895 3927
rect 8018 3924 8024 3936
rect 7883 3896 8024 3924
rect 7883 3893 7895 3896
rect 7837 3887 7895 3893
rect 8018 3884 8024 3896
rect 8076 3884 8082 3936
rect 9815 3927 9873 3933
rect 9815 3893 9827 3927
rect 9861 3924 9873 3927
rect 10042 3924 10048 3936
rect 9861 3896 10048 3924
rect 9861 3893 9873 3896
rect 9815 3887 9873 3893
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10226 3924 10232 3936
rect 10187 3896 10232 3924
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 12250 3924 12256 3936
rect 12211 3896 12256 3924
rect 12250 3884 12256 3896
rect 12308 3884 12314 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 13262 3924 13268 3936
rect 12492 3896 13268 3924
rect 12492 3884 12498 3896
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 14936 3924 14964 4100
rect 15470 4088 15476 4100
rect 15528 4088 15534 4140
rect 16025 4131 16083 4137
rect 16025 4097 16037 4131
rect 16071 4128 16083 4131
rect 16390 4128 16396 4140
rect 16071 4100 16396 4128
rect 16071 4097 16083 4100
rect 16025 4091 16083 4097
rect 16390 4088 16396 4100
rect 16448 4088 16454 4140
rect 18233 4131 18291 4137
rect 18233 4097 18245 4131
rect 18279 4128 18291 4131
rect 18506 4128 18512 4140
rect 18279 4100 18512 4128
rect 18279 4097 18291 4100
rect 18233 4091 18291 4097
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 15013 3995 15071 4001
rect 15013 3961 15025 3995
rect 15059 3992 15071 3995
rect 15378 3992 15384 4004
rect 15059 3964 15384 3992
rect 15059 3961 15071 3964
rect 15013 3955 15071 3961
rect 15378 3952 15384 3964
rect 15436 3952 15442 4004
rect 15488 3992 15516 4088
rect 15488 3964 15792 3992
rect 15194 3924 15200 3936
rect 14936 3896 15200 3924
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 15470 3884 15476 3936
rect 15528 3924 15534 3936
rect 15764 3933 15792 3964
rect 15565 3927 15623 3933
rect 15565 3924 15577 3927
rect 15528 3896 15577 3924
rect 15528 3884 15534 3896
rect 15565 3893 15577 3896
rect 15611 3893 15623 3927
rect 15565 3887 15623 3893
rect 15749 3927 15807 3933
rect 15749 3893 15761 3927
rect 15795 3893 15807 3927
rect 15749 3887 15807 3893
rect 368 3834 18860 3856
rect 368 3782 3478 3834
rect 3530 3782 3542 3834
rect 3594 3782 3606 3834
rect 3658 3782 3670 3834
rect 3722 3782 3734 3834
rect 3786 3782 6578 3834
rect 6630 3782 6642 3834
rect 6694 3782 6706 3834
rect 6758 3782 6770 3834
rect 6822 3782 6834 3834
rect 6886 3782 9678 3834
rect 9730 3782 9742 3834
rect 9794 3782 9806 3834
rect 9858 3782 9870 3834
rect 9922 3782 9934 3834
rect 9986 3782 12778 3834
rect 12830 3782 12842 3834
rect 12894 3782 12906 3834
rect 12958 3782 12970 3834
rect 13022 3782 13034 3834
rect 13086 3782 15878 3834
rect 15930 3782 15942 3834
rect 15994 3782 16006 3834
rect 16058 3782 16070 3834
rect 16122 3782 16134 3834
rect 16186 3782 18860 3834
rect 368 3760 18860 3782
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 4433 3723 4491 3729
rect 4433 3720 4445 3723
rect 3936 3692 4445 3720
rect 3936 3680 3942 3692
rect 4433 3689 4445 3692
rect 4479 3689 4491 3723
rect 4433 3683 4491 3689
rect 6454 3680 6460 3732
rect 6512 3720 6518 3732
rect 6549 3723 6607 3729
rect 6549 3720 6561 3723
rect 6512 3692 6561 3720
rect 6512 3680 6518 3692
rect 6549 3689 6561 3692
rect 6595 3689 6607 3723
rect 6549 3683 6607 3689
rect 7558 3680 7564 3732
rect 7616 3720 7622 3732
rect 7926 3720 7932 3732
rect 7616 3692 7932 3720
rect 7616 3680 7622 3692
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 8202 3720 8208 3732
rect 8163 3692 8208 3720
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 13262 3680 13268 3732
rect 13320 3720 13326 3732
rect 16298 3720 16304 3732
rect 13320 3692 16304 3720
rect 13320 3680 13326 3692
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 10226 3652 10232 3664
rect 6472 3624 7788 3652
rect 10187 3624 10232 3652
rect 201 3587 259 3593
rect 201 3553 213 3587
rect 247 3584 259 3587
rect 2130 3584 2136 3596
rect 247 3556 2136 3584
rect 247 3553 259 3556
rect 201 3547 259 3553
rect 952 3525 980 3556
rect 2130 3544 2136 3556
rect 2188 3544 2194 3596
rect 3881 3587 3939 3593
rect 3881 3553 3893 3587
rect 3927 3584 3939 3587
rect 4430 3584 4436 3596
rect 3927 3556 4436 3584
rect 3927 3553 3939 3556
rect 3881 3547 3939 3553
rect 4430 3544 4436 3556
rect 4488 3584 4494 3596
rect 4488 3556 5304 3584
rect 4488 3544 4494 3556
rect 937 3519 995 3525
rect 937 3485 949 3519
rect 983 3485 995 3519
rect 4062 3516 4068 3528
rect 4023 3488 4068 3516
rect 937 3479 995 3485
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 5276 3525 5304 3556
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 5445 3519 5503 3525
rect 5445 3485 5457 3519
rect 5491 3485 5503 3519
rect 5445 3479 5503 3485
rect 2406 3448 2412 3460
rect 2367 3420 2412 3448
rect 2406 3408 2412 3420
rect 2464 3408 2470 3460
rect 3878 3448 3884 3460
rect 3634 3434 3884 3448
rect 3620 3420 3884 3434
rect 845 3383 903 3389
rect 845 3380 857 3383
rect 308 3352 857 3380
rect 308 3040 336 3352
rect 845 3349 857 3352
rect 891 3349 903 3383
rect 845 3343 903 3349
rect 2774 3340 2780 3392
rect 2832 3380 2838 3392
rect 3620 3380 3648 3420
rect 3878 3408 3884 3420
rect 3936 3408 3942 3460
rect 4706 3408 4712 3460
rect 4764 3448 4770 3460
rect 5460 3448 5488 3479
rect 6362 3476 6368 3528
rect 6420 3516 6426 3528
rect 6472 3525 6500 3624
rect 6932 3556 7686 3584
rect 6932 3528 6960 3556
rect 6457 3519 6515 3525
rect 6457 3516 6469 3519
rect 6420 3488 6469 3516
rect 6420 3476 6426 3488
rect 6457 3485 6469 3488
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3516 6699 3519
rect 6914 3516 6920 3528
rect 6687 3488 6920 3516
rect 6687 3485 6699 3488
rect 6641 3479 6699 3485
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7549 3525 7555 3528
rect 7525 3519 7555 3525
rect 7525 3485 7537 3519
rect 7525 3479 7555 3485
rect 7549 3476 7555 3479
rect 7607 3476 7613 3528
rect 7658 3525 7686 3556
rect 7760 3535 7788 3624
rect 10226 3612 10232 3624
rect 10284 3612 10290 3664
rect 12713 3655 12771 3661
rect 12713 3621 12725 3655
rect 12759 3621 12771 3655
rect 12713 3615 12771 3621
rect 13173 3655 13231 3661
rect 13173 3621 13185 3655
rect 13219 3652 13231 3655
rect 13725 3655 13783 3661
rect 13725 3652 13737 3655
rect 13219 3624 13737 3652
rect 13219 3621 13231 3624
rect 13173 3615 13231 3621
rect 13725 3621 13737 3624
rect 13771 3621 13783 3655
rect 13725 3615 13783 3621
rect 7929 3587 7987 3593
rect 7929 3553 7941 3587
rect 7975 3584 7987 3587
rect 8389 3587 8447 3593
rect 8389 3584 8401 3587
rect 7975 3556 8401 3584
rect 7975 3553 7987 3556
rect 7929 3547 7987 3553
rect 8389 3553 8401 3556
rect 8435 3553 8447 3587
rect 10042 3584 10048 3596
rect 8389 3547 8447 3553
rect 8496 3556 10048 3584
rect 7745 3529 7803 3535
rect 7643 3519 7701 3525
rect 7643 3485 7655 3519
rect 7689 3485 7701 3519
rect 7745 3495 7757 3529
rect 7791 3495 7803 3529
rect 8496 3525 8524 3556
rect 10042 3544 10048 3556
rect 10100 3544 10106 3596
rect 10686 3544 10692 3596
rect 10744 3584 10750 3596
rect 11333 3587 11391 3593
rect 11333 3584 11345 3587
rect 10744 3556 11345 3584
rect 10744 3544 10750 3556
rect 11333 3553 11345 3556
rect 11379 3553 11391 3587
rect 12728 3584 12756 3615
rect 13357 3587 13415 3593
rect 12728 3556 13032 3584
rect 11333 3547 11391 3553
rect 7745 3489 7803 3495
rect 8481 3519 8539 3525
rect 7643 3479 7701 3485
rect 8481 3485 8493 3519
rect 8527 3485 8539 3519
rect 8846 3516 8852 3528
rect 8807 3488 8852 3516
rect 8481 3479 8539 3485
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 10502 3516 10508 3528
rect 9999 3488 10508 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 4764 3420 5488 3448
rect 4764 3408 4770 3420
rect 7926 3408 7932 3460
rect 7984 3448 7990 3460
rect 9968 3448 9996 3479
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 11589 3519 11647 3525
rect 11589 3516 11601 3519
rect 11296 3488 11601 3516
rect 11296 3476 11302 3488
rect 11589 3485 11601 3488
rect 11635 3516 11647 3519
rect 12066 3516 12072 3528
rect 11635 3488 12072 3516
rect 11635 3485 11647 3488
rect 11589 3479 11647 3485
rect 12066 3476 12072 3488
rect 12124 3516 12130 3528
rect 13004 3525 13032 3556
rect 13357 3553 13369 3587
rect 13403 3584 13415 3587
rect 13909 3587 13967 3593
rect 13909 3584 13921 3587
rect 13403 3556 13676 3584
rect 13403 3553 13415 3556
rect 13357 3547 13415 3553
rect 12897 3519 12955 3525
rect 12124 3488 12434 3516
rect 12124 3476 12130 3488
rect 10594 3448 10600 3460
rect 7984 3420 9996 3448
rect 10244 3420 10600 3448
rect 7984 3408 7990 3420
rect 2832 3352 3648 3380
rect 4249 3383 4307 3389
rect 2832 3340 2838 3352
rect 4249 3349 4261 3383
rect 4295 3380 4307 3383
rect 4338 3380 4344 3392
rect 4295 3352 4344 3380
rect 4295 3349 4307 3352
rect 4249 3343 4307 3349
rect 4338 3340 4344 3352
rect 4396 3340 4402 3392
rect 5353 3383 5411 3389
rect 5353 3349 5365 3383
rect 5399 3380 5411 3383
rect 5810 3380 5816 3392
rect 5399 3352 5816 3380
rect 5399 3349 5411 3352
rect 5353 3343 5411 3349
rect 5810 3340 5816 3352
rect 5868 3340 5874 3392
rect 9309 3383 9367 3389
rect 9309 3349 9321 3383
rect 9355 3380 9367 3383
rect 10244 3380 10272 3420
rect 10594 3408 10600 3420
rect 10652 3408 10658 3460
rect 12406 3448 12434 3488
rect 12897 3485 12909 3519
rect 12943 3485 12955 3519
rect 12897 3479 12955 3485
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3516 13047 3519
rect 13265 3519 13323 3525
rect 13265 3516 13277 3519
rect 13035 3488 13277 3516
rect 13035 3485 13047 3488
rect 12989 3479 13047 3485
rect 13265 3485 13277 3488
rect 13311 3485 13323 3519
rect 13446 3516 13452 3528
rect 13407 3488 13452 3516
rect 13265 3479 13323 3485
rect 12912 3448 12940 3479
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 13648 3525 13676 3556
rect 13740 3556 13921 3584
rect 13740 3528 13768 3556
rect 13909 3553 13921 3556
rect 13955 3553 13967 3587
rect 13909 3547 13967 3553
rect 14090 3544 14096 3596
rect 14148 3584 14154 3596
rect 14185 3587 14243 3593
rect 14185 3584 14197 3587
rect 14148 3556 14197 3584
rect 14148 3544 14154 3556
rect 14185 3553 14197 3556
rect 14231 3553 14243 3587
rect 14185 3547 14243 3553
rect 16298 3544 16304 3596
rect 16356 3584 16362 3596
rect 18230 3584 18236 3596
rect 16356 3556 18236 3584
rect 16356 3544 16362 3556
rect 18230 3544 18236 3556
rect 18288 3544 18294 3596
rect 13633 3519 13691 3525
rect 13633 3485 13645 3519
rect 13679 3485 13691 3519
rect 13633 3479 13691 3485
rect 13722 3476 13728 3528
rect 13780 3476 13786 3528
rect 15194 3476 15200 3528
rect 15252 3516 15258 3528
rect 16482 3516 16488 3528
rect 15252 3488 16488 3516
rect 15252 3476 15258 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 17862 3516 17868 3528
rect 17823 3488 17868 3516
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 13464 3448 13492 3476
rect 12406 3420 13492 3448
rect 14452 3451 14510 3457
rect 14452 3417 14464 3451
rect 14498 3448 14510 3451
rect 15286 3448 15292 3460
rect 14498 3420 15292 3448
rect 14498 3417 14510 3420
rect 14452 3411 14510 3417
rect 15286 3408 15292 3420
rect 15344 3408 15350 3460
rect 16206 3448 16212 3460
rect 15764 3420 16212 3448
rect 15764 3392 15792 3420
rect 16206 3408 16212 3420
rect 16264 3448 16270 3460
rect 16264 3420 16882 3448
rect 16264 3408 16270 3420
rect 10410 3380 10416 3392
rect 9355 3352 10272 3380
rect 10371 3352 10416 3380
rect 9355 3349 9367 3352
rect 9309 3343 9367 3349
rect 10410 3340 10416 3352
rect 10468 3340 10474 3392
rect 13909 3383 13967 3389
rect 13909 3349 13921 3383
rect 13955 3380 13967 3383
rect 15194 3380 15200 3392
rect 13955 3352 15200 3380
rect 13955 3349 13967 3352
rect 13909 3343 13967 3349
rect 15194 3340 15200 3352
rect 15252 3340 15258 3392
rect 15565 3383 15623 3389
rect 15565 3349 15577 3383
rect 15611 3380 15623 3383
rect 15654 3380 15660 3392
rect 15611 3352 15660 3380
rect 15611 3349 15623 3352
rect 15565 3343 15623 3349
rect 15654 3340 15660 3352
rect 15712 3340 15718 3392
rect 15746 3340 15752 3392
rect 15804 3380 15810 3392
rect 16114 3380 16120 3392
rect 15804 3352 15849 3380
rect 16075 3352 16120 3380
rect 15804 3340 15810 3352
rect 16114 3340 16120 3352
rect 16172 3380 16178 3392
rect 16390 3380 16396 3392
rect 16172 3352 16396 3380
rect 16172 3340 16178 3352
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 368 3290 18860 3312
rect 368 3238 5028 3290
rect 5080 3238 5092 3290
rect 5144 3238 5156 3290
rect 5208 3238 5220 3290
rect 5272 3238 5284 3290
rect 5336 3238 8128 3290
rect 8180 3238 8192 3290
rect 8244 3238 8256 3290
rect 8308 3238 8320 3290
rect 8372 3238 8384 3290
rect 8436 3238 11228 3290
rect 11280 3238 11292 3290
rect 11344 3238 11356 3290
rect 11408 3238 11420 3290
rect 11472 3238 11484 3290
rect 11536 3238 14328 3290
rect 14380 3238 14392 3290
rect 14444 3238 14456 3290
rect 14508 3238 14520 3290
rect 14572 3238 14584 3290
rect 14636 3238 17428 3290
rect 17480 3238 17492 3290
rect 17544 3238 17556 3290
rect 17608 3238 17620 3290
rect 17672 3238 17684 3290
rect 17736 3238 18860 3290
rect 368 3216 18860 3238
rect 2406 3136 2412 3188
rect 2464 3176 2470 3188
rect 3421 3179 3479 3185
rect 3421 3176 3433 3179
rect 2464 3148 3433 3176
rect 2464 3136 2470 3148
rect 3421 3145 3433 3148
rect 3467 3145 3479 3179
rect 3421 3139 3479 3145
rect 6825 3179 6883 3185
rect 6825 3145 6837 3179
rect 6871 3176 6883 3179
rect 7190 3176 7196 3188
rect 6871 3148 7196 3176
rect 6871 3145 6883 3148
rect 6825 3139 6883 3145
rect 7190 3136 7196 3148
rect 7248 3136 7254 3188
rect 10226 3176 10232 3188
rect 7484 3148 10232 3176
rect 2774 3108 2780 3120
rect 2070 3080 2780 3108
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 4062 3108 4068 3120
rect 3620 3080 4068 3108
rect 661 3043 719 3049
rect 661 3040 673 3043
rect 308 3012 673 3040
rect 661 3009 673 3012
rect 707 3009 719 3043
rect 661 3003 719 3009
rect 3050 3000 3056 3052
rect 3108 3040 3114 3052
rect 3145 3043 3203 3049
rect 3145 3040 3157 3043
rect 3108 3012 3157 3040
rect 3108 3000 3114 3012
rect 3145 3009 3157 3012
rect 3191 3009 3203 3043
rect 3145 3003 3203 3009
rect 3326 3000 3332 3052
rect 3384 3040 3390 3052
rect 3620 3049 3648 3080
rect 4062 3068 4068 3080
rect 4120 3068 4126 3120
rect 4338 3108 4344 3120
rect 4299 3080 4344 3108
rect 4338 3068 4344 3080
rect 4396 3068 4402 3120
rect 5718 3068 5724 3120
rect 5776 3108 5782 3120
rect 7374 3108 7380 3120
rect 5776 3080 7380 3108
rect 5776 3068 5782 3080
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 3384 3012 3617 3040
rect 3384 3000 3390 3012
rect 3605 3009 3617 3012
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3009 3755 3043
rect 3970 3040 3976 3052
rect 3931 3012 3976 3040
rect 3697 3003 3755 3009
rect 1029 2975 1087 2981
rect 1029 2941 1041 2975
rect 1075 2972 1087 2975
rect 3712 2972 3740 3003
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 4430 3040 4436 3052
rect 4080 3012 4436 3040
rect 4080 2972 4108 3012
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 4706 3040 4712 3052
rect 4667 3012 4712 3040
rect 4706 3000 4712 3012
rect 4764 3000 4770 3052
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3040 5135 3043
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 5123 3012 5273 3040
rect 5123 3009 5135 3012
rect 5077 3003 5135 3009
rect 5261 3009 5273 3012
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 5445 3043 5503 3049
rect 5445 3009 5457 3043
rect 5491 3009 5503 3043
rect 5810 3040 5816 3052
rect 5771 3012 5816 3040
rect 5445 3003 5503 3009
rect 1075 2944 2544 2972
rect 3712 2944 4108 2972
rect 4157 2975 4215 2981
rect 1075 2941 1087 2944
rect 1029 2935 1087 2941
rect 2516 2904 2544 2944
rect 4157 2941 4169 2975
rect 4203 2941 4215 2975
rect 4157 2935 4215 2941
rect 4525 2975 4583 2981
rect 4525 2941 4537 2975
rect 4571 2972 4583 2975
rect 5460 2972 5488 3003
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 5920 3049 5948 3080
rect 7374 3068 7380 3080
rect 7432 3068 7438 3120
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3009 5963 3043
rect 5905 3003 5963 3009
rect 6086 3000 6092 3052
rect 6144 3040 6150 3052
rect 6181 3043 6239 3049
rect 6181 3040 6193 3043
rect 6144 3012 6193 3040
rect 6144 3000 6150 3012
rect 6181 3009 6193 3012
rect 6227 3040 6239 3043
rect 7190 3040 7196 3052
rect 6227 3012 7196 3040
rect 6227 3009 6239 3012
rect 6181 3003 6239 3009
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 7484 3040 7512 3148
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 10502 3136 10508 3188
rect 10560 3176 10566 3188
rect 13081 3179 13139 3185
rect 10560 3148 12434 3176
rect 10560 3136 10566 3148
rect 9214 3108 9220 3120
rect 9062 3080 9220 3108
rect 9214 3068 9220 3080
rect 9272 3068 9278 3120
rect 10321 3111 10379 3117
rect 10321 3077 10333 3111
rect 10367 3108 10379 3111
rect 12406 3108 12434 3148
rect 13081 3145 13093 3179
rect 13127 3176 13139 3179
rect 13170 3176 13176 3188
rect 13127 3148 13176 3176
rect 13127 3145 13139 3148
rect 13081 3139 13139 3145
rect 13170 3136 13176 3148
rect 13228 3176 13234 3188
rect 13722 3176 13728 3188
rect 13228 3148 13728 3176
rect 13228 3136 13234 3148
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 15286 3176 15292 3188
rect 13832 3148 15292 3176
rect 13832 3108 13860 3148
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 15381 3179 15439 3185
rect 15381 3145 15393 3179
rect 15427 3145 15439 3179
rect 16482 3176 16488 3188
rect 16443 3148 16488 3176
rect 15381 3139 15439 3145
rect 15396 3108 15424 3139
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 10367 3080 11192 3108
rect 12406 3080 13860 3108
rect 15304 3080 15424 3108
rect 10367 3077 10379 3080
rect 10321 3071 10379 3077
rect 11164 3052 11192 3080
rect 7300 3012 7512 3040
rect 7653 3043 7711 3049
rect 7300 2972 7328 3012
rect 7653 3009 7665 3043
rect 7699 3040 7711 3043
rect 7926 3040 7932 3052
rect 7699 3012 7932 3040
rect 7699 3009 7711 3012
rect 7653 3003 7711 3009
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 9447 3043 9505 3049
rect 9447 3009 9459 3043
rect 9493 3040 9505 3043
rect 9769 3043 9827 3049
rect 9769 3040 9781 3043
rect 9493 3012 9781 3040
rect 9493 3009 9505 3012
rect 9447 3003 9505 3009
rect 9769 3009 9781 3012
rect 9815 3040 9827 3043
rect 10042 3040 10048 3052
rect 9815 3012 10048 3040
rect 9815 3009 9827 3012
rect 9769 3003 9827 3009
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 10137 3043 10195 3049
rect 10137 3009 10149 3043
rect 10183 3040 10195 3043
rect 10226 3040 10232 3052
rect 10183 3012 10232 3040
rect 10183 3009 10195 3012
rect 10137 3003 10195 3009
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 10410 3040 10416 3052
rect 10371 3012 10416 3040
rect 10410 3000 10416 3012
rect 10468 3000 10474 3052
rect 10778 3040 10784 3052
rect 10739 3012 10784 3040
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 11146 3040 11152 3052
rect 11107 3012 11152 3040
rect 11146 3000 11152 3012
rect 11204 3000 11210 3052
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 13280 3049 13308 3080
rect 12713 3043 12771 3049
rect 12713 3040 12725 3043
rect 11848 3012 12725 3040
rect 11848 3000 11854 3012
rect 12713 3009 12725 3012
rect 12759 3009 12771 3043
rect 12713 3003 12771 3009
rect 13265 3043 13323 3049
rect 13265 3009 13277 3043
rect 13311 3009 13323 3043
rect 13265 3003 13323 3009
rect 13446 3000 13452 3052
rect 13504 3040 13510 3052
rect 13541 3043 13599 3049
rect 13541 3040 13553 3043
rect 13504 3012 13553 3040
rect 13504 3000 13510 3012
rect 13541 3009 13553 3012
rect 13587 3009 13599 3043
rect 13541 3003 13599 3009
rect 13998 3000 14004 3052
rect 14056 3040 14062 3052
rect 15013 3043 15071 3049
rect 15013 3040 15025 3043
rect 14056 3012 15025 3040
rect 14056 3000 14062 3012
rect 15013 3009 15025 3012
rect 15059 3009 15071 3043
rect 15194 3040 15200 3052
rect 15155 3012 15200 3040
rect 15013 3003 15071 3009
rect 15194 3000 15200 3012
rect 15252 3000 15258 3052
rect 15304 3049 15332 3080
rect 15470 3068 15476 3120
rect 15528 3108 15534 3120
rect 15654 3108 15660 3120
rect 15528 3080 15573 3108
rect 15615 3080 15660 3108
rect 15528 3068 15534 3080
rect 15654 3068 15660 3080
rect 15712 3068 15718 3120
rect 15289 3043 15347 3049
rect 15289 3009 15301 3043
rect 15335 3009 15347 3043
rect 15289 3003 15347 3009
rect 15378 3000 15384 3052
rect 15436 3040 15442 3052
rect 16393 3043 16451 3049
rect 15436 3012 15481 3040
rect 15436 3000 15442 3012
rect 16393 3009 16405 3043
rect 16439 3009 16451 3043
rect 16393 3003 16451 3009
rect 7466 2972 7472 2984
rect 4571 2944 5488 2972
rect 6104 2944 7328 2972
rect 7427 2944 7472 2972
rect 4571 2941 4583 2944
rect 4525 2935 4583 2941
rect 3510 2904 3516 2916
rect 2516 2876 3516 2904
rect 3510 2864 3516 2876
rect 3568 2864 3574 2916
rect 3694 2864 3700 2916
rect 3752 2904 3758 2916
rect 3973 2907 4031 2913
rect 3973 2904 3985 2907
rect 3752 2876 3985 2904
rect 3752 2864 3758 2876
rect 3973 2873 3985 2876
rect 4019 2873 4031 2907
rect 4172 2904 4200 2935
rect 6104 2913 6132 2944
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 8021 2975 8079 2981
rect 8021 2972 8033 2975
rect 7576 2944 8033 2972
rect 4801 2907 4859 2913
rect 4801 2904 4813 2907
rect 4172 2876 4813 2904
rect 3973 2867 4031 2873
rect 4801 2873 4813 2876
rect 4847 2904 4859 2907
rect 5077 2907 5135 2913
rect 5077 2904 5089 2907
rect 4847 2876 5089 2904
rect 4847 2873 4859 2876
rect 4801 2867 4859 2873
rect 5077 2873 5089 2876
rect 5123 2873 5135 2907
rect 5077 2867 5135 2873
rect 5353 2907 5411 2913
rect 5353 2873 5365 2907
rect 5399 2904 5411 2907
rect 6089 2907 6147 2913
rect 5399 2876 5948 2904
rect 5399 2873 5411 2876
rect 5353 2867 5411 2873
rect 2498 2845 2504 2848
rect 2455 2839 2504 2845
rect 2455 2805 2467 2839
rect 2501 2805 2504 2839
rect 2455 2799 2504 2805
rect 2498 2796 2504 2799
rect 2556 2796 2562 2848
rect 2685 2839 2743 2845
rect 2685 2805 2697 2839
rect 2731 2836 2743 2839
rect 2774 2836 2780 2848
rect 2731 2808 2780 2836
rect 2731 2805 2743 2808
rect 2685 2799 2743 2805
rect 2774 2796 2780 2808
rect 2832 2796 2838 2848
rect 3237 2839 3295 2845
rect 3237 2805 3249 2839
rect 3283 2836 3295 2839
rect 5368 2836 5396 2867
rect 5810 2836 5816 2848
rect 3283 2808 5396 2836
rect 5771 2808 5816 2836
rect 3283 2805 3295 2808
rect 3237 2799 3295 2805
rect 5810 2796 5816 2808
rect 5868 2796 5874 2848
rect 5920 2836 5948 2876
rect 6089 2873 6101 2907
rect 6135 2873 6147 2907
rect 7098 2904 7104 2916
rect 6089 2867 6147 2873
rect 6194 2876 7104 2904
rect 6194 2836 6222 2876
rect 7098 2864 7104 2876
rect 7156 2864 7162 2916
rect 7282 2864 7288 2916
rect 7340 2904 7346 2916
rect 7576 2904 7604 2944
rect 8021 2941 8033 2944
rect 8067 2941 8079 2975
rect 8021 2935 8079 2941
rect 8570 2932 8576 2984
rect 8628 2972 8634 2984
rect 9677 2975 9735 2981
rect 9677 2972 9689 2975
rect 8628 2944 9689 2972
rect 8628 2932 8634 2944
rect 9677 2941 9689 2944
rect 9723 2941 9735 2975
rect 9677 2935 9735 2941
rect 10873 2975 10931 2981
rect 10873 2941 10885 2975
rect 10919 2972 10931 2975
rect 12434 2972 12440 2984
rect 10919 2944 12440 2972
rect 10919 2941 10931 2944
rect 10873 2935 10931 2941
rect 12434 2932 12440 2944
rect 12492 2932 12498 2984
rect 16114 2972 16120 2984
rect 14108 2944 16120 2972
rect 7340 2876 7604 2904
rect 7340 2864 7346 2876
rect 11054 2864 11060 2916
rect 11112 2904 11118 2916
rect 11112 2876 13400 2904
rect 11112 2864 11118 2876
rect 5920 2808 6222 2836
rect 7009 2839 7067 2845
rect 7009 2805 7021 2839
rect 7055 2836 7067 2839
rect 7650 2836 7656 2848
rect 7055 2808 7656 2836
rect 7055 2805 7067 2808
rect 7009 2799 7067 2805
rect 7650 2796 7656 2808
rect 7708 2796 7714 2848
rect 12618 2796 12624 2848
rect 12676 2836 12682 2848
rect 12805 2839 12863 2845
rect 12805 2836 12817 2839
rect 12676 2808 12817 2836
rect 12676 2796 12682 2808
rect 12805 2805 12817 2808
rect 12851 2805 12863 2839
rect 13372 2836 13400 2876
rect 13449 2839 13507 2845
rect 13449 2836 13461 2839
rect 13372 2808 13461 2836
rect 12805 2799 12863 2805
rect 13449 2805 13461 2808
rect 13495 2836 13507 2839
rect 14108 2836 14136 2944
rect 16114 2932 16120 2944
rect 16172 2972 16178 2984
rect 16408 2972 16436 3003
rect 16172 2944 16436 2972
rect 16172 2932 16178 2944
rect 13495 2808 14136 2836
rect 13495 2805 13507 2808
rect 13449 2799 13507 2805
rect 14182 2796 14188 2848
rect 14240 2836 14246 2848
rect 14829 2839 14887 2845
rect 14829 2836 14841 2839
rect 14240 2808 14841 2836
rect 14240 2796 14246 2808
rect 14829 2805 14841 2808
rect 14875 2805 14887 2839
rect 14829 2799 14887 2805
rect 368 2746 18860 2768
rect 368 2694 3478 2746
rect 3530 2694 3542 2746
rect 3594 2694 3606 2746
rect 3658 2694 3670 2746
rect 3722 2694 3734 2746
rect 3786 2694 6578 2746
rect 6630 2694 6642 2746
rect 6694 2694 6706 2746
rect 6758 2694 6770 2746
rect 6822 2694 6834 2746
rect 6886 2694 9678 2746
rect 9730 2694 9742 2746
rect 9794 2694 9806 2746
rect 9858 2694 9870 2746
rect 9922 2694 9934 2746
rect 9986 2694 12778 2746
rect 12830 2694 12842 2746
rect 12894 2694 12906 2746
rect 12958 2694 12970 2746
rect 13022 2694 13034 2746
rect 13086 2694 15878 2746
rect 15930 2694 15942 2746
rect 15994 2694 16006 2746
rect 16058 2694 16070 2746
rect 16122 2694 16134 2746
rect 16186 2694 18860 2746
rect 368 2672 18860 2694
rect 1489 2635 1547 2641
rect 1489 2601 1501 2635
rect 1535 2632 1547 2635
rect 3970 2632 3976 2644
rect 1535 2604 3976 2632
rect 1535 2601 1547 2604
rect 1489 2595 1547 2601
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 4893 2635 4951 2641
rect 4893 2632 4905 2635
rect 4632 2604 4905 2632
rect 1397 2567 1455 2573
rect 1397 2533 1409 2567
rect 1443 2564 1455 2567
rect 3142 2564 3148 2576
rect 1443 2536 3148 2564
rect 1443 2533 1455 2536
rect 1397 2527 1455 2533
rect 3142 2524 3148 2536
rect 3200 2564 3206 2576
rect 3200 2536 4200 2564
rect 3200 2524 3206 2536
rect 658 2456 664 2508
rect 716 2496 722 2508
rect 1029 2499 1087 2505
rect 1029 2496 1041 2499
rect 716 2468 1041 2496
rect 716 2456 722 2468
rect 1029 2465 1041 2468
rect 1075 2496 1087 2499
rect 1857 2499 1915 2505
rect 1857 2496 1869 2499
rect 1075 2468 1869 2496
rect 1075 2465 1087 2468
rect 1029 2459 1087 2465
rect 1857 2465 1869 2468
rect 1903 2496 1915 2499
rect 2682 2496 2688 2508
rect 1903 2468 2688 2496
rect 1903 2465 1915 2468
rect 1857 2459 1915 2465
rect 2682 2456 2688 2468
rect 2740 2456 2746 2508
rect 3326 2496 3332 2508
rect 3287 2468 3332 2496
rect 3326 2456 3332 2468
rect 3384 2456 3390 2508
rect 4172 2505 4200 2536
rect 4157 2499 4215 2505
rect 4157 2465 4169 2499
rect 4203 2465 4215 2499
rect 4157 2459 4215 2465
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2428 2007 2431
rect 2593 2431 2651 2437
rect 2593 2428 2605 2431
rect 1995 2400 2605 2428
rect 1995 2397 2007 2400
rect 1949 2391 2007 2397
rect 2593 2397 2605 2400
rect 2639 2428 2651 2431
rect 2958 2428 2964 2440
rect 2639 2400 2964 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 3234 2428 3240 2440
rect 3195 2400 3240 2428
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 3878 2428 3884 2440
rect 3839 2400 3884 2428
rect 3878 2388 3884 2400
rect 3936 2428 3942 2440
rect 4632 2428 4660 2604
rect 4893 2601 4905 2604
rect 4939 2601 4951 2635
rect 11287 2635 11345 2641
rect 11287 2632 11299 2635
rect 4893 2595 4951 2601
rect 6472 2604 7972 2632
rect 5902 2564 5908 2576
rect 4724 2536 5908 2564
rect 4724 2437 4752 2536
rect 5902 2524 5908 2536
rect 5960 2524 5966 2576
rect 4893 2499 4951 2505
rect 4893 2465 4905 2499
rect 4939 2496 4951 2499
rect 5537 2499 5595 2505
rect 5537 2496 5549 2499
rect 4939 2468 5549 2496
rect 4939 2465 4951 2468
rect 4893 2459 4951 2465
rect 5537 2465 5549 2468
rect 5583 2496 5595 2499
rect 6472 2496 6500 2604
rect 6641 2567 6699 2573
rect 6641 2533 6653 2567
rect 6687 2533 6699 2567
rect 6914 2564 6920 2576
rect 6875 2536 6920 2564
rect 6641 2527 6699 2533
rect 5583 2468 6500 2496
rect 6656 2496 6684 2527
rect 6914 2524 6920 2536
rect 6972 2524 6978 2576
rect 7282 2524 7288 2576
rect 7340 2564 7346 2576
rect 7340 2536 7385 2564
rect 7340 2524 7346 2536
rect 6656 2468 7236 2496
rect 5583 2465 5595 2468
rect 5537 2459 5595 2465
rect 3936 2400 4660 2428
rect 4709 2431 4767 2437
rect 3936 2388 3942 2400
rect 4709 2397 4721 2431
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 5353 2431 5411 2437
rect 5353 2397 5365 2431
rect 5399 2428 5411 2431
rect 5442 2428 5448 2440
rect 5399 2400 5448 2428
rect 5399 2397 5411 2400
rect 5353 2391 5411 2397
rect 2317 2363 2375 2369
rect 2317 2329 2329 2363
rect 2363 2360 2375 2363
rect 3050 2360 3056 2372
rect 2363 2332 3056 2360
rect 2363 2329 2375 2332
rect 2317 2323 2375 2329
rect 3050 2320 3056 2332
rect 3108 2320 3114 2372
rect 3602 2320 3608 2372
rect 3660 2360 3666 2372
rect 4724 2360 4752 2391
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 5810 2428 5816 2440
rect 5771 2400 5816 2428
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 5994 2428 6000 2440
rect 5955 2400 6000 2428
rect 5994 2388 6000 2400
rect 6052 2388 6058 2440
rect 6454 2428 6460 2440
rect 6415 2400 6460 2428
rect 6454 2388 6460 2400
rect 6512 2388 6518 2440
rect 6575 2431 6633 2437
rect 6575 2428 6587 2431
rect 6564 2397 6587 2428
rect 6621 2397 6633 2431
rect 7006 2428 7012 2440
rect 6967 2400 7012 2428
rect 6564 2391 6633 2397
rect 5718 2360 5724 2372
rect 3660 2332 4752 2360
rect 5460 2332 5724 2360
rect 3660 2320 3666 2332
rect 1670 2292 1676 2304
rect 1631 2264 1676 2292
rect 1670 2252 1676 2264
rect 1728 2252 1734 2304
rect 2038 2252 2044 2304
rect 2096 2292 2102 2304
rect 2774 2292 2780 2304
rect 2096 2264 2780 2292
rect 2096 2252 2102 2264
rect 2774 2252 2780 2264
rect 2832 2292 2838 2304
rect 3970 2292 3976 2304
rect 2832 2264 3976 2292
rect 2832 2252 2838 2264
rect 3970 2252 3976 2264
rect 4028 2252 4034 2304
rect 4890 2252 4896 2304
rect 4948 2292 4954 2304
rect 5460 2301 5488 2332
rect 5718 2320 5724 2332
rect 5776 2320 5782 2372
rect 5828 2360 5856 2388
rect 6564 2360 6592 2391
rect 7006 2388 7012 2400
rect 7064 2388 7070 2440
rect 7208 2437 7236 2468
rect 7944 2440 7972 2604
rect 9876 2604 11299 2632
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2496 8171 2499
rect 8846 2496 8852 2508
rect 8159 2468 8852 2496
rect 8159 2465 8171 2468
rect 8113 2459 8171 2465
rect 8846 2456 8852 2468
rect 8904 2456 8910 2508
rect 7193 2431 7251 2437
rect 7193 2397 7205 2431
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 7282 2388 7288 2440
rect 7340 2428 7346 2440
rect 7340 2400 7385 2428
rect 7340 2388 7346 2400
rect 7466 2388 7472 2440
rect 7524 2428 7530 2440
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7524 2400 7849 2428
rect 7524 2388 7530 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 7377 2363 7435 2369
rect 7377 2360 7389 2363
rect 5828 2332 6592 2360
rect 6656 2332 7389 2360
rect 4985 2295 5043 2301
rect 4985 2292 4997 2295
rect 4948 2264 4997 2292
rect 4948 2252 4954 2264
rect 4985 2261 4997 2264
rect 5031 2261 5043 2295
rect 4985 2255 5043 2261
rect 5445 2295 5503 2301
rect 5445 2261 5457 2295
rect 5491 2261 5503 2295
rect 5445 2255 5503 2261
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 5813 2295 5871 2301
rect 5813 2292 5825 2295
rect 5592 2264 5825 2292
rect 5592 2252 5598 2264
rect 5813 2261 5825 2264
rect 5859 2261 5871 2295
rect 5813 2255 5871 2261
rect 5902 2252 5908 2304
rect 5960 2292 5966 2304
rect 6656 2292 6684 2332
rect 7377 2329 7389 2332
rect 7423 2329 7435 2363
rect 7852 2360 7880 2391
rect 7926 2388 7932 2440
rect 7984 2428 7990 2440
rect 9876 2437 9904 2604
rect 11287 2601 11299 2604
rect 11333 2632 11345 2635
rect 11790 2632 11796 2644
rect 11333 2604 11796 2632
rect 11333 2601 11345 2604
rect 11287 2595 11345 2601
rect 11790 2592 11796 2604
rect 11848 2592 11854 2644
rect 12250 2632 12256 2644
rect 11992 2604 12256 2632
rect 10229 2567 10287 2573
rect 10229 2533 10241 2567
rect 10275 2564 10287 2567
rect 10778 2564 10784 2576
rect 10275 2536 10784 2564
rect 10275 2533 10287 2536
rect 10229 2527 10287 2533
rect 10778 2524 10784 2536
rect 10836 2524 10842 2576
rect 11698 2524 11704 2576
rect 11756 2564 11762 2576
rect 11992 2564 12020 2604
rect 12250 2592 12256 2604
rect 12308 2632 12314 2644
rect 13446 2632 13452 2644
rect 12308 2604 13452 2632
rect 12308 2592 12314 2604
rect 13446 2592 13452 2604
rect 13504 2632 13510 2644
rect 13633 2635 13691 2641
rect 13633 2632 13645 2635
rect 13504 2604 13645 2632
rect 13504 2592 13510 2604
rect 13633 2601 13645 2604
rect 13679 2632 13691 2635
rect 14550 2632 14556 2644
rect 13679 2604 14556 2632
rect 13679 2601 13691 2604
rect 13633 2595 13691 2601
rect 14550 2592 14556 2604
rect 14608 2632 14614 2644
rect 15102 2632 15108 2644
rect 14608 2604 15108 2632
rect 14608 2592 14614 2604
rect 15102 2592 15108 2604
rect 15160 2632 15166 2644
rect 15746 2632 15752 2644
rect 15160 2604 15752 2632
rect 15160 2592 15166 2604
rect 15746 2592 15752 2604
rect 15804 2632 15810 2644
rect 16025 2635 16083 2641
rect 16025 2632 16037 2635
rect 15804 2604 16037 2632
rect 15804 2592 15810 2604
rect 16025 2601 16037 2604
rect 16071 2601 16083 2635
rect 16025 2595 16083 2601
rect 11756 2536 12020 2564
rect 11756 2524 11762 2536
rect 13078 2524 13084 2576
rect 13136 2564 13142 2576
rect 13173 2567 13231 2573
rect 13173 2564 13185 2567
rect 13136 2536 13185 2564
rect 13136 2524 13142 2536
rect 13173 2533 13185 2536
rect 13219 2533 13231 2567
rect 16040 2564 16068 2595
rect 16040 2536 16896 2564
rect 13173 2527 13231 2533
rect 9953 2499 10011 2505
rect 9953 2465 9965 2499
rect 9999 2496 10011 2499
rect 10042 2496 10048 2508
rect 9999 2468 10048 2496
rect 9999 2465 10011 2468
rect 9953 2459 10011 2465
rect 10042 2456 10048 2468
rect 10100 2456 10106 2508
rect 11054 2496 11060 2508
rect 11015 2468 11060 2496
rect 11054 2456 11060 2468
rect 11112 2456 11118 2508
rect 14093 2499 14151 2505
rect 13096 2468 13860 2496
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7984 2400 8033 2428
rect 7984 2388 7990 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 9033 2431 9091 2437
rect 9033 2397 9045 2431
rect 9079 2397 9091 2431
rect 9033 2391 9091 2397
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2397 9643 2431
rect 9585 2391 9643 2397
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 12713 2431 12771 2437
rect 12713 2397 12725 2431
rect 12759 2428 12771 2431
rect 12986 2428 12992 2440
rect 12759 2400 12992 2428
rect 12759 2397 12771 2400
rect 12713 2391 12771 2397
rect 8849 2363 8907 2369
rect 8849 2360 8861 2363
rect 7852 2332 8861 2360
rect 7377 2323 7435 2329
rect 8849 2329 8861 2332
rect 8895 2329 8907 2363
rect 8849 2323 8907 2329
rect 5960 2264 6684 2292
rect 5960 2252 5966 2264
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 9048 2292 9076 2391
rect 9600 2360 9628 2391
rect 12986 2388 12992 2400
rect 13044 2388 13050 2440
rect 13096 2437 13124 2468
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 13189 2431 13247 2437
rect 13189 2397 13201 2431
rect 13235 2428 13247 2431
rect 13354 2428 13360 2440
rect 13235 2400 13360 2428
rect 13235 2397 13247 2400
rect 13189 2391 13247 2397
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 13832 2437 13860 2468
rect 14093 2465 14105 2499
rect 14139 2496 14151 2499
rect 14182 2496 14188 2508
rect 14139 2468 14188 2496
rect 14139 2465 14151 2468
rect 14093 2459 14151 2465
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 15286 2456 15292 2508
rect 15344 2496 15350 2508
rect 16209 2499 16267 2505
rect 16209 2496 16221 2499
rect 15344 2468 16221 2496
rect 15344 2456 15350 2468
rect 16209 2465 16221 2468
rect 16255 2465 16267 2499
rect 16209 2459 16267 2465
rect 13817 2431 13875 2437
rect 13817 2397 13829 2431
rect 13863 2397 13875 2431
rect 16868 2414 16896 2536
rect 18230 2496 18236 2508
rect 18191 2468 18236 2496
rect 18230 2456 18236 2468
rect 18288 2456 18294 2508
rect 13817 2391 13875 2397
rect 10226 2360 10232 2372
rect 9600 2332 10232 2360
rect 10226 2320 10232 2332
rect 10284 2320 10290 2372
rect 11698 2320 11704 2372
rect 11756 2320 11762 2372
rect 13265 2363 13323 2369
rect 13265 2329 13277 2363
rect 13311 2329 13323 2363
rect 13265 2323 13323 2329
rect 13449 2363 13507 2369
rect 13449 2329 13461 2363
rect 13495 2360 13507 2363
rect 13538 2360 13544 2372
rect 13495 2332 13544 2360
rect 13495 2329 13507 2332
rect 13449 2323 13507 2329
rect 7156 2264 9076 2292
rect 7156 2252 7162 2264
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10597 2295 10655 2301
rect 10597 2292 10609 2295
rect 10376 2264 10609 2292
rect 10376 2252 10382 2264
rect 10597 2261 10609 2264
rect 10643 2261 10655 2295
rect 10597 2255 10655 2261
rect 12434 2252 12440 2304
rect 12492 2292 12498 2304
rect 13280 2292 13308 2323
rect 13538 2320 13544 2332
rect 13596 2320 13602 2372
rect 13832 2360 13860 2391
rect 14090 2360 14096 2372
rect 13832 2332 14096 2360
rect 14090 2320 14096 2332
rect 14148 2320 14154 2372
rect 14550 2320 14556 2372
rect 14608 2320 14614 2372
rect 15838 2360 15844 2372
rect 15799 2332 15844 2360
rect 15838 2320 15844 2332
rect 15896 2320 15902 2372
rect 17954 2360 17960 2372
rect 17915 2332 17960 2360
rect 17954 2320 17960 2332
rect 18012 2320 18018 2372
rect 14734 2292 14740 2304
rect 12492 2264 14740 2292
rect 12492 2252 12498 2264
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 368 2202 18860 2224
rect 368 2150 5028 2202
rect 5080 2150 5092 2202
rect 5144 2150 5156 2202
rect 5208 2150 5220 2202
rect 5272 2150 5284 2202
rect 5336 2150 8128 2202
rect 8180 2150 8192 2202
rect 8244 2150 8256 2202
rect 8308 2150 8320 2202
rect 8372 2150 8384 2202
rect 8436 2150 11228 2202
rect 11280 2150 11292 2202
rect 11344 2150 11356 2202
rect 11408 2150 11420 2202
rect 11472 2150 11484 2202
rect 11536 2150 14328 2202
rect 14380 2150 14392 2202
rect 14444 2150 14456 2202
rect 14508 2150 14520 2202
rect 14572 2150 14584 2202
rect 14636 2150 17428 2202
rect 17480 2150 17492 2202
rect 17544 2150 17556 2202
rect 17608 2150 17620 2202
rect 17672 2150 17684 2202
rect 17736 2150 18860 2202
rect 368 2128 18860 2150
rect 658 2088 664 2100
rect 619 2060 664 2088
rect 658 2048 664 2060
rect 716 2048 722 2100
rect 2593 2091 2651 2097
rect 2593 2057 2605 2091
rect 2639 2088 2651 2091
rect 2958 2088 2964 2100
rect 2639 2060 2774 2088
rect 2919 2060 2964 2088
rect 2639 2057 2651 2060
rect 2593 2051 2651 2057
rect 2038 2020 2044 2032
rect 1702 1992 2044 2020
rect 2038 1980 2044 1992
rect 2096 1980 2102 2032
rect 2130 1980 2136 2032
rect 2188 2020 2194 2032
rect 2746 2020 2774 2060
rect 2958 2048 2964 2060
rect 3016 2048 3022 2100
rect 3602 2088 3608 2100
rect 3528 2060 3608 2088
rect 3234 2020 3240 2032
rect 2188 1992 2452 2020
rect 2746 1992 3240 2020
rect 2188 1980 2194 1992
rect 2424 1961 2452 1992
rect 3234 1980 3240 1992
rect 3292 1980 3298 2032
rect 2409 1955 2467 1961
rect 2409 1921 2421 1955
rect 2455 1921 2467 1955
rect 2409 1915 2467 1921
rect 2498 1912 2504 1964
rect 2556 1952 2562 1964
rect 2556 1924 2601 1952
rect 2556 1912 2562 1924
rect 2682 1912 2688 1964
rect 2740 1952 2746 1964
rect 3053 1955 3111 1961
rect 2740 1924 2833 1952
rect 2740 1912 2746 1924
rect 3053 1921 3065 1955
rect 3099 1952 3111 1955
rect 3142 1952 3148 1964
rect 3099 1924 3148 1952
rect 3099 1921 3111 1924
rect 3053 1915 3111 1921
rect 3142 1912 3148 1924
rect 3200 1912 3206 1964
rect 3528 1961 3556 2060
rect 3602 2048 3608 2060
rect 3660 2048 3666 2100
rect 7282 2048 7288 2100
rect 7340 2088 7346 2100
rect 7653 2091 7711 2097
rect 7653 2088 7665 2091
rect 7340 2060 7665 2088
rect 7340 2048 7346 2060
rect 7653 2057 7665 2060
rect 7699 2057 7711 2091
rect 8478 2088 8484 2100
rect 7653 2051 7711 2057
rect 7760 2060 8484 2088
rect 5626 2020 5632 2032
rect 4264 1992 5632 2020
rect 3421 1955 3479 1961
rect 3421 1921 3433 1955
rect 3467 1921 3479 1955
rect 3421 1915 3479 1921
rect 3513 1955 3571 1961
rect 3513 1921 3525 1955
rect 3559 1921 3571 1955
rect 3513 1915 3571 1921
rect 1670 1844 1676 1896
rect 1728 1884 1734 1896
rect 2133 1887 2191 1893
rect 2133 1884 2145 1887
rect 1728 1856 2145 1884
rect 1728 1844 1734 1856
rect 2133 1853 2145 1856
rect 2179 1853 2191 1887
rect 2700 1884 2728 1912
rect 3436 1884 3464 1915
rect 3602 1912 3608 1964
rect 3660 1952 3666 1964
rect 3660 1924 3705 1952
rect 3660 1912 3666 1924
rect 3878 1912 3884 1964
rect 3936 1952 3942 1964
rect 4264 1961 4292 1992
rect 5626 1980 5632 1992
rect 5684 1980 5690 2032
rect 6914 1980 6920 2032
rect 6972 2020 6978 2032
rect 7760 2029 7788 2060
rect 8478 2048 8484 2060
rect 8536 2048 8542 2100
rect 10318 2048 10324 2100
rect 10376 2048 10382 2100
rect 12805 2091 12863 2097
rect 12805 2057 12817 2091
rect 12851 2088 12863 2091
rect 13354 2088 13360 2100
rect 12851 2060 13360 2088
rect 12851 2057 12863 2060
rect 12805 2051 12863 2057
rect 13354 2048 13360 2060
rect 13412 2048 13418 2100
rect 13538 2088 13544 2100
rect 13499 2060 13544 2088
rect 13538 2048 13544 2060
rect 13596 2048 13602 2100
rect 13630 2048 13636 2100
rect 13688 2088 13694 2100
rect 15562 2088 15568 2100
rect 13688 2060 15568 2088
rect 13688 2048 13694 2060
rect 7745 2023 7803 2029
rect 7745 2020 7757 2023
rect 6972 1992 7757 2020
rect 6972 1980 6978 1992
rect 7745 1989 7757 1992
rect 7791 1989 7803 2023
rect 8573 2023 8631 2029
rect 7745 1983 7803 1989
rect 8220 1992 8524 2020
rect 4157 1955 4215 1961
rect 4157 1952 4169 1955
rect 3936 1924 4169 1952
rect 3936 1912 3942 1924
rect 4157 1921 4169 1924
rect 4203 1921 4215 1955
rect 4157 1915 4215 1921
rect 4249 1955 4307 1961
rect 4249 1921 4261 1955
rect 4295 1921 4307 1955
rect 4249 1915 4307 1921
rect 4890 1912 4896 1964
rect 4948 1952 4954 1964
rect 5261 1955 5319 1961
rect 5261 1952 5273 1955
rect 4948 1924 5273 1952
rect 4948 1912 4954 1924
rect 5261 1921 5273 1924
rect 5307 1921 5319 1955
rect 5261 1915 5319 1921
rect 5445 1955 5503 1961
rect 5445 1921 5457 1955
rect 5491 1952 5503 1955
rect 5534 1952 5540 1964
rect 5491 1924 5540 1952
rect 5491 1921 5503 1924
rect 5445 1915 5503 1921
rect 5534 1912 5540 1924
rect 5592 1912 5598 1964
rect 5994 1952 6000 1964
rect 5736 1924 6000 1952
rect 4065 1887 4123 1893
rect 4065 1884 4077 1887
rect 2700 1856 3372 1884
rect 3436 1856 4077 1884
rect 2133 1847 2191 1853
rect 3050 1776 3056 1828
rect 3108 1816 3114 1828
rect 3237 1819 3295 1825
rect 3237 1816 3249 1819
rect 3108 1788 3249 1816
rect 3108 1776 3114 1788
rect 3237 1785 3249 1788
rect 3283 1785 3295 1819
rect 3344 1816 3372 1856
rect 4065 1853 4077 1856
rect 4111 1884 4123 1887
rect 5736 1884 5764 1924
rect 5994 1912 6000 1924
rect 6052 1952 6058 1964
rect 7650 1952 7656 1964
rect 6052 1924 7512 1952
rect 7611 1924 7656 1952
rect 6052 1912 6058 1924
rect 4111 1856 5764 1884
rect 5813 1887 5871 1893
rect 4111 1853 4123 1856
rect 4065 1847 4123 1853
rect 5813 1853 5825 1887
rect 5859 1884 5871 1887
rect 6362 1884 6368 1896
rect 5859 1856 6368 1884
rect 5859 1853 5871 1856
rect 5813 1847 5871 1853
rect 6362 1844 6368 1856
rect 6420 1844 6426 1896
rect 7484 1884 7512 1924
rect 7650 1912 7656 1924
rect 7708 1912 7714 1964
rect 7929 1955 7987 1961
rect 7929 1921 7941 1955
rect 7975 1952 7987 1955
rect 8110 1952 8116 1964
rect 7975 1924 8116 1952
rect 7975 1921 7987 1924
rect 7929 1915 7987 1921
rect 8110 1912 8116 1924
rect 8168 1912 8174 1964
rect 8220 1961 8248 1992
rect 8205 1955 8263 1961
rect 8205 1921 8217 1955
rect 8251 1921 8263 1955
rect 8205 1915 8263 1921
rect 8389 1955 8447 1961
rect 8389 1921 8401 1955
rect 8435 1921 8447 1955
rect 8496 1952 8524 1992
rect 8573 1989 8585 2023
rect 8619 2020 8631 2023
rect 8846 2020 8852 2032
rect 8619 1992 8852 2020
rect 8619 1989 8631 1992
rect 8573 1983 8631 1989
rect 8846 1980 8852 1992
rect 8904 1980 8910 2032
rect 10336 2020 10364 2048
rect 12253 2023 12311 2029
rect 12253 2020 12265 2023
rect 9876 1992 10364 2020
rect 10704 1992 12265 2020
rect 9876 1961 9904 1992
rect 8757 1955 8815 1961
rect 8757 1952 8769 1955
rect 8496 1924 8769 1952
rect 8389 1915 8447 1921
rect 8757 1921 8769 1924
rect 8803 1921 8815 1955
rect 8757 1915 8815 1921
rect 9861 1955 9919 1961
rect 9861 1921 9873 1955
rect 9907 1921 9919 1955
rect 9861 1915 9919 1921
rect 10321 1955 10379 1961
rect 10321 1921 10333 1955
rect 10367 1952 10379 1955
rect 10502 1952 10508 1964
rect 10367 1924 10508 1952
rect 10367 1921 10379 1924
rect 10321 1915 10379 1921
rect 8220 1884 8248 1915
rect 7484 1856 8248 1884
rect 3510 1816 3516 1828
rect 3344 1788 3516 1816
rect 3237 1779 3295 1785
rect 3510 1776 3516 1788
rect 3568 1776 3574 1828
rect 8404 1816 8432 1915
rect 10502 1912 10508 1924
rect 10560 1912 10566 1964
rect 10226 1884 10232 1896
rect 10187 1856 10232 1884
rect 10226 1844 10232 1856
rect 10284 1844 10290 1896
rect 10244 1816 10272 1844
rect 8404 1788 10272 1816
rect 3881 1751 3939 1757
rect 3881 1717 3893 1751
rect 3927 1748 3939 1751
rect 3970 1748 3976 1760
rect 3927 1720 3976 1748
rect 3927 1717 3939 1720
rect 3881 1711 3939 1717
rect 3970 1708 3976 1720
rect 4028 1708 4034 1760
rect 4341 1751 4399 1757
rect 4341 1717 4353 1751
rect 4387 1748 4399 1751
rect 4706 1748 4712 1760
rect 4387 1720 4712 1748
rect 4387 1717 4399 1720
rect 4341 1711 4399 1717
rect 4706 1708 4712 1720
rect 4764 1708 4770 1760
rect 5350 1748 5356 1760
rect 5311 1720 5356 1748
rect 5350 1708 5356 1720
rect 5408 1708 5414 1760
rect 7006 1708 7012 1760
rect 7064 1748 7070 1760
rect 8849 1751 8907 1757
rect 8849 1748 8861 1751
rect 7064 1720 8861 1748
rect 7064 1708 7070 1720
rect 8849 1717 8861 1720
rect 8895 1748 8907 1751
rect 9214 1748 9220 1760
rect 8895 1720 9220 1748
rect 8895 1717 8907 1720
rect 8849 1711 8907 1717
rect 9214 1708 9220 1720
rect 9272 1708 9278 1760
rect 9401 1751 9459 1757
rect 9401 1717 9413 1751
rect 9447 1748 9459 1751
rect 9490 1748 9496 1760
rect 9447 1720 9496 1748
rect 9447 1717 9459 1720
rect 9401 1711 9459 1717
rect 9490 1708 9496 1720
rect 9548 1708 9554 1760
rect 9582 1708 9588 1760
rect 9640 1748 9646 1760
rect 10704 1748 10732 1992
rect 12253 1989 12265 1992
rect 12299 1989 12311 2023
rect 12253 1983 12311 1989
rect 12360 1992 13860 2020
rect 10781 1955 10839 1961
rect 10781 1921 10793 1955
rect 10827 1952 10839 1955
rect 11054 1952 11060 1964
rect 10827 1924 11060 1952
rect 10827 1921 10839 1924
rect 10781 1915 10839 1921
rect 11054 1912 11060 1924
rect 11112 1912 11118 1964
rect 11238 1912 11244 1964
rect 11296 1952 11302 1964
rect 12360 1952 12388 1992
rect 11296 1924 12388 1952
rect 11296 1912 11302 1924
rect 12618 1912 12624 1964
rect 12676 1952 12682 1964
rect 12989 1955 13047 1961
rect 12989 1952 13001 1955
rect 12676 1924 13001 1952
rect 12676 1912 12682 1924
rect 12989 1921 13001 1924
rect 13035 1921 13047 1955
rect 12989 1915 13047 1921
rect 10962 1884 10968 1896
rect 10923 1856 10968 1884
rect 10962 1844 10968 1856
rect 11020 1844 11026 1896
rect 13004 1884 13032 1915
rect 13078 1912 13084 1964
rect 13136 1952 13142 1964
rect 13832 1961 13860 1992
rect 13209 1955 13267 1961
rect 13136 1924 13181 1952
rect 13136 1912 13142 1924
rect 13209 1921 13221 1955
rect 13255 1952 13267 1955
rect 13633 1955 13691 1961
rect 13633 1952 13645 1955
rect 13255 1924 13645 1952
rect 13255 1921 13267 1924
rect 13209 1915 13267 1921
rect 13633 1921 13645 1924
rect 13679 1952 13691 1955
rect 13817 1955 13875 1961
rect 13679 1924 13768 1952
rect 13679 1921 13691 1924
rect 13633 1915 13691 1921
rect 13740 1896 13768 1924
rect 13817 1921 13829 1955
rect 13863 1952 13875 1955
rect 14182 1952 14188 1964
rect 13863 1924 14188 1952
rect 13863 1921 13875 1924
rect 13817 1915 13875 1921
rect 14182 1912 14188 1924
rect 14240 1952 14246 1964
rect 14384 1961 14412 2060
rect 15562 2048 15568 2060
rect 15620 2048 15626 2100
rect 15657 2091 15715 2097
rect 15657 2057 15669 2091
rect 15703 2088 15715 2091
rect 17221 2091 17279 2097
rect 17221 2088 17233 2091
rect 15703 2060 17233 2088
rect 15703 2057 15715 2060
rect 15657 2051 15715 2057
rect 17221 2057 17233 2060
rect 17267 2057 17279 2091
rect 17681 2091 17739 2097
rect 17681 2088 17693 2091
rect 17221 2051 17279 2057
rect 17328 2060 17693 2088
rect 14553 2023 14611 2029
rect 14553 1989 14565 2023
rect 14599 2020 14611 2023
rect 14734 2020 14740 2032
rect 14599 1992 14740 2020
rect 14599 1989 14611 1992
rect 14553 1983 14611 1989
rect 14734 1980 14740 1992
rect 14792 1980 14798 2032
rect 15286 1980 15292 2032
rect 15344 2020 15350 2032
rect 15749 2023 15807 2029
rect 15749 2020 15761 2023
rect 15344 1992 15761 2020
rect 15344 1980 15350 1992
rect 15749 1989 15761 1992
rect 15795 2020 15807 2023
rect 17328 2020 17356 2060
rect 17681 2057 17693 2060
rect 17727 2057 17739 2091
rect 18138 2088 18144 2100
rect 18099 2060 18144 2088
rect 17681 2051 17739 2057
rect 18138 2048 18144 2060
rect 18196 2048 18202 2100
rect 15795 1992 17356 2020
rect 17589 2023 17647 2029
rect 15795 1989 15807 1992
rect 15749 1983 15807 1989
rect 17589 1989 17601 2023
rect 17635 2020 17647 2023
rect 18230 2020 18236 2032
rect 17635 1992 18236 2020
rect 17635 1989 17647 1992
rect 17589 1983 17647 1989
rect 18230 1980 18236 1992
rect 18288 1980 18294 2032
rect 14277 1955 14335 1961
rect 14277 1952 14289 1955
rect 14240 1924 14289 1952
rect 14240 1912 14246 1924
rect 14277 1921 14289 1924
rect 14323 1921 14335 1955
rect 14277 1915 14335 1921
rect 14369 1955 14427 1961
rect 14369 1921 14381 1955
rect 14415 1921 14427 1955
rect 14369 1915 14427 1921
rect 16485 1955 16543 1961
rect 16485 1921 16497 1955
rect 16531 1952 16543 1955
rect 17218 1952 17224 1964
rect 16531 1924 17224 1952
rect 16531 1921 16543 1924
rect 16485 1915 16543 1921
rect 17218 1912 17224 1924
rect 17276 1912 17282 1964
rect 18046 1952 18052 1964
rect 18007 1924 18052 1952
rect 18046 1912 18052 1924
rect 18104 1912 18110 1964
rect 18506 1952 18512 1964
rect 18467 1924 18512 1952
rect 18506 1912 18512 1924
rect 18564 1912 18570 1964
rect 13357 1887 13415 1893
rect 13357 1884 13369 1887
rect 13004 1856 13369 1884
rect 13357 1853 13369 1856
rect 13403 1853 13415 1887
rect 13357 1847 13415 1853
rect 13722 1844 13728 1896
rect 13780 1844 13786 1896
rect 15838 1884 15844 1896
rect 14384 1856 15844 1884
rect 9640 1720 10732 1748
rect 9640 1708 9646 1720
rect 11146 1708 11152 1760
rect 11204 1748 11210 1760
rect 11241 1751 11299 1757
rect 11241 1748 11253 1751
rect 11204 1720 11253 1748
rect 11204 1708 11210 1720
rect 11241 1717 11253 1720
rect 11287 1748 11299 1751
rect 11698 1748 11704 1760
rect 11287 1720 11704 1748
rect 11287 1717 11299 1720
rect 11241 1711 11299 1717
rect 11698 1708 11704 1720
rect 11756 1708 11762 1760
rect 12250 1748 12256 1760
rect 12163 1720 12256 1748
rect 12250 1708 12256 1720
rect 12308 1748 12314 1760
rect 14384 1748 14412 1856
rect 15838 1844 15844 1856
rect 15896 1884 15902 1896
rect 16574 1884 16580 1896
rect 15896 1856 16436 1884
rect 16535 1856 16580 1884
rect 15896 1844 15902 1856
rect 14918 1776 14924 1828
rect 14976 1816 14982 1828
rect 16117 1819 16175 1825
rect 16117 1816 16129 1819
rect 14976 1788 16129 1816
rect 14976 1776 14982 1788
rect 16117 1785 16129 1788
rect 16163 1785 16175 1819
rect 16408 1816 16436 1856
rect 16574 1844 16580 1856
rect 16632 1844 16638 1896
rect 16669 1887 16727 1893
rect 16669 1853 16681 1887
rect 16715 1853 16727 1887
rect 17862 1884 17868 1896
rect 17823 1856 17868 1884
rect 16669 1847 16727 1853
rect 16684 1816 16712 1847
rect 17862 1844 17868 1856
rect 17920 1844 17926 1896
rect 16408 1788 16712 1816
rect 16117 1779 16175 1785
rect 12308 1720 14412 1748
rect 14461 1751 14519 1757
rect 12308 1708 12314 1720
rect 14461 1717 14473 1751
rect 14507 1748 14519 1751
rect 14734 1748 14740 1760
rect 14507 1720 14740 1748
rect 14507 1717 14519 1720
rect 14461 1711 14519 1717
rect 14734 1708 14740 1720
rect 14792 1708 14798 1760
rect 15286 1748 15292 1760
rect 15247 1720 15292 1748
rect 15286 1708 15292 1720
rect 15344 1708 15350 1760
rect 18322 1748 18328 1760
rect 18283 1720 18328 1748
rect 18322 1708 18328 1720
rect 18380 1708 18386 1760
rect 368 1658 18860 1680
rect 368 1606 3478 1658
rect 3530 1606 3542 1658
rect 3594 1606 3606 1658
rect 3658 1606 3670 1658
rect 3722 1606 3734 1658
rect 3786 1606 6578 1658
rect 6630 1606 6642 1658
rect 6694 1606 6706 1658
rect 6758 1606 6770 1658
rect 6822 1606 6834 1658
rect 6886 1606 9678 1658
rect 9730 1606 9742 1658
rect 9794 1606 9806 1658
rect 9858 1606 9870 1658
rect 9922 1606 9934 1658
rect 9986 1606 12778 1658
rect 12830 1606 12842 1658
rect 12894 1606 12906 1658
rect 12958 1606 12970 1658
rect 13022 1606 13034 1658
rect 13086 1606 15878 1658
rect 15930 1606 15942 1658
rect 15994 1606 16006 1658
rect 16058 1606 16070 1658
rect 16122 1606 16134 1658
rect 16186 1606 18860 1658
rect 368 1584 18860 1606
rect 5353 1547 5411 1553
rect 5353 1513 5365 1547
rect 5399 1544 5411 1547
rect 5442 1544 5448 1556
rect 5399 1516 5448 1544
rect 5399 1513 5411 1516
rect 5353 1507 5411 1513
rect 5442 1504 5448 1516
rect 5500 1504 5506 1556
rect 7926 1504 7932 1556
rect 7984 1544 7990 1556
rect 7984 1516 8892 1544
rect 7984 1504 7990 1516
rect 4525 1479 4583 1485
rect 4525 1476 4537 1479
rect 3620 1448 4537 1476
rect 2130 1408 2136 1420
rect 2091 1380 2136 1408
rect 2130 1368 2136 1380
rect 2188 1368 2194 1420
rect 2409 1411 2467 1417
rect 2409 1377 2421 1411
rect 2455 1408 2467 1411
rect 3620 1408 3648 1448
rect 4525 1445 4537 1448
rect 4571 1445 4583 1479
rect 8294 1476 8300 1488
rect 4525 1439 4583 1445
rect 6012 1448 8300 1476
rect 2455 1380 3648 1408
rect 4433 1411 4491 1417
rect 2455 1377 2467 1380
rect 2409 1371 2467 1377
rect 4433 1377 4445 1411
rect 4479 1408 4491 1411
rect 5350 1408 5356 1420
rect 4479 1380 5356 1408
rect 4479 1377 4491 1380
rect 4433 1371 4491 1377
rect 5350 1368 5356 1380
rect 5408 1368 5414 1420
rect 5718 1368 5724 1420
rect 5776 1408 5782 1420
rect 6012 1417 6040 1448
rect 8294 1436 8300 1448
rect 8352 1476 8358 1488
rect 8864 1476 8892 1516
rect 9214 1504 9220 1556
rect 9272 1544 9278 1556
rect 12434 1544 12440 1556
rect 9272 1516 12440 1544
rect 9272 1504 9278 1516
rect 9306 1476 9312 1488
rect 8352 1448 8524 1476
rect 8864 1448 9312 1476
rect 8352 1436 8358 1448
rect 5813 1411 5871 1417
rect 5813 1408 5825 1411
rect 5776 1380 5825 1408
rect 5776 1368 5782 1380
rect 5813 1377 5825 1380
rect 5859 1377 5871 1411
rect 5813 1371 5871 1377
rect 5997 1411 6055 1417
rect 5997 1377 6009 1411
rect 6043 1377 6055 1411
rect 5997 1371 6055 1377
rect 7745 1411 7803 1417
rect 7745 1377 7757 1411
rect 7791 1408 7803 1411
rect 7926 1408 7932 1420
rect 7791 1380 7932 1408
rect 7791 1377 7803 1380
rect 7745 1371 7803 1377
rect 7926 1368 7932 1380
rect 7984 1368 7990 1420
rect 8496 1417 8524 1448
rect 9306 1436 9312 1448
rect 9364 1476 9370 1488
rect 9582 1476 9588 1488
rect 9364 1448 9588 1476
rect 9364 1436 9370 1448
rect 9582 1436 9588 1448
rect 9640 1436 9646 1488
rect 10318 1476 10324 1488
rect 9784 1448 10324 1476
rect 8481 1411 8539 1417
rect 8481 1377 8493 1411
rect 8527 1408 8539 1411
rect 8662 1408 8668 1420
rect 8527 1380 8668 1408
rect 8527 1377 8539 1380
rect 8481 1371 8539 1377
rect 8662 1368 8668 1380
rect 8720 1368 8726 1420
rect 9784 1417 9812 1448
rect 10318 1436 10324 1448
rect 10376 1436 10382 1488
rect 11241 1479 11299 1485
rect 11241 1476 11253 1479
rect 10980 1448 11253 1476
rect 9769 1411 9827 1417
rect 9769 1377 9781 1411
rect 9815 1377 9827 1411
rect 9769 1371 9827 1377
rect 9861 1411 9919 1417
rect 9861 1377 9873 1411
rect 9907 1377 9919 1411
rect 9861 1371 9919 1377
rect 3970 1340 3976 1352
rect 3542 1312 3976 1340
rect 3970 1300 3976 1312
rect 4028 1300 4034 1352
rect 4614 1340 4620 1352
rect 4575 1312 4620 1340
rect 4614 1300 4620 1312
rect 4672 1300 4678 1352
rect 4709 1343 4767 1349
rect 4709 1309 4721 1343
rect 4755 1309 4767 1343
rect 4709 1303 4767 1309
rect 4724 1272 4752 1303
rect 4798 1300 4804 1352
rect 4856 1340 4862 1352
rect 4985 1343 5043 1349
rect 4985 1340 4997 1343
rect 4856 1312 4997 1340
rect 4856 1300 4862 1312
rect 4985 1309 4997 1312
rect 5031 1309 5043 1343
rect 4985 1303 5043 1309
rect 6362 1300 6368 1352
rect 6420 1340 6426 1352
rect 6457 1343 6515 1349
rect 6457 1340 6469 1343
rect 6420 1312 6469 1340
rect 6420 1300 6426 1312
rect 6457 1309 6469 1312
rect 6503 1309 6515 1343
rect 6457 1303 6515 1309
rect 6641 1343 6699 1349
rect 6641 1309 6653 1343
rect 6687 1309 6699 1343
rect 6641 1303 6699 1309
rect 6917 1343 6975 1349
rect 6917 1309 6929 1343
rect 6963 1340 6975 1343
rect 7282 1340 7288 1352
rect 6963 1312 7288 1340
rect 6963 1309 6975 1312
rect 6917 1303 6975 1309
rect 4893 1275 4951 1281
rect 4893 1272 4905 1275
rect 3896 1244 4660 1272
rect 4724 1244 4905 1272
rect 3896 1213 3924 1244
rect 3881 1207 3939 1213
rect 3881 1173 3893 1207
rect 3927 1173 3939 1207
rect 3881 1167 3939 1173
rect 3970 1164 3976 1216
rect 4028 1204 4034 1216
rect 4157 1207 4215 1213
rect 4157 1204 4169 1207
rect 4028 1176 4169 1204
rect 4028 1164 4034 1176
rect 4157 1173 4169 1176
rect 4203 1173 4215 1207
rect 4632 1204 4660 1244
rect 4893 1241 4905 1244
rect 4939 1272 4951 1275
rect 5721 1275 5779 1281
rect 5721 1272 5733 1275
rect 4939 1244 5733 1272
rect 4939 1241 4951 1244
rect 4893 1235 4951 1241
rect 5721 1241 5733 1244
rect 5767 1241 5779 1275
rect 6656 1272 6684 1303
rect 7282 1300 7288 1312
rect 7340 1300 7346 1352
rect 8202 1340 8208 1352
rect 7392 1312 8208 1340
rect 6656 1244 7144 1272
rect 5721 1235 5779 1241
rect 4798 1204 4804 1216
rect 4632 1176 4804 1204
rect 4157 1167 4215 1173
rect 4798 1164 4804 1176
rect 4856 1164 4862 1216
rect 6086 1164 6092 1216
rect 6144 1204 6150 1216
rect 6457 1207 6515 1213
rect 6457 1204 6469 1207
rect 6144 1176 6469 1204
rect 6144 1164 6150 1176
rect 6457 1173 6469 1176
rect 6503 1173 6515 1207
rect 6457 1167 6515 1173
rect 6825 1207 6883 1213
rect 6825 1173 6837 1207
rect 6871 1204 6883 1207
rect 6914 1204 6920 1216
rect 6871 1176 6920 1204
rect 6871 1173 6883 1176
rect 6825 1167 6883 1173
rect 6914 1164 6920 1176
rect 6972 1164 6978 1216
rect 7116 1213 7144 1244
rect 7101 1207 7159 1213
rect 7101 1173 7113 1207
rect 7147 1173 7159 1207
rect 7101 1167 7159 1173
rect 7190 1164 7196 1216
rect 7248 1204 7254 1216
rect 7392 1204 7420 1312
rect 8202 1300 8208 1312
rect 8260 1340 8266 1352
rect 8389 1343 8447 1349
rect 8389 1340 8401 1343
rect 8260 1312 8401 1340
rect 8260 1300 8266 1312
rect 8389 1309 8401 1312
rect 8435 1309 8447 1343
rect 8680 1340 8708 1368
rect 9876 1340 9904 1371
rect 10594 1340 10600 1352
rect 8680 1312 9904 1340
rect 10555 1312 10600 1340
rect 8389 1303 8447 1309
rect 10594 1300 10600 1312
rect 10652 1300 10658 1352
rect 10689 1343 10747 1349
rect 10689 1309 10701 1343
rect 10735 1309 10747 1343
rect 10980 1340 11008 1448
rect 11241 1445 11253 1448
rect 11287 1445 11299 1479
rect 11241 1439 11299 1445
rect 11057 1343 11115 1349
rect 11057 1340 11069 1343
rect 10980 1312 11069 1340
rect 10689 1303 10747 1309
rect 11057 1309 11069 1312
rect 11103 1309 11115 1343
rect 11238 1340 11244 1352
rect 11199 1312 11244 1340
rect 11057 1303 11115 1309
rect 7469 1275 7527 1281
rect 7469 1241 7481 1275
rect 7515 1272 7527 1275
rect 8297 1275 8355 1281
rect 7515 1244 7972 1272
rect 7515 1241 7527 1244
rect 7469 1235 7527 1241
rect 7944 1213 7972 1244
rect 8297 1241 8309 1275
rect 8343 1272 8355 1275
rect 8478 1272 8484 1284
rect 8343 1244 8484 1272
rect 8343 1241 8355 1244
rect 8297 1235 8355 1241
rect 8478 1232 8484 1244
rect 8536 1232 8542 1284
rect 10704 1272 10732 1303
rect 11238 1300 11244 1312
rect 11296 1300 11302 1352
rect 11532 1349 11560 1516
rect 12434 1504 12440 1516
rect 12492 1504 12498 1556
rect 13722 1504 13728 1556
rect 13780 1544 13786 1556
rect 17862 1544 17868 1556
rect 13780 1516 17868 1544
rect 13780 1504 13786 1516
rect 17862 1504 17868 1516
rect 17920 1504 17926 1556
rect 17954 1504 17960 1556
rect 18012 1544 18018 1556
rect 18049 1547 18107 1553
rect 18049 1544 18061 1547
rect 18012 1516 18061 1544
rect 18012 1504 18018 1516
rect 18049 1513 18061 1516
rect 18095 1513 18107 1547
rect 18506 1544 18512 1556
rect 18467 1516 18512 1544
rect 18049 1507 18107 1513
rect 18506 1504 18512 1516
rect 18564 1504 18570 1556
rect 12250 1408 12256 1420
rect 12211 1380 12256 1408
rect 12250 1368 12256 1380
rect 12308 1368 12314 1420
rect 13078 1408 13084 1420
rect 13039 1380 13084 1408
rect 13078 1368 13084 1380
rect 13136 1368 13142 1420
rect 13265 1411 13323 1417
rect 13265 1377 13277 1411
rect 13311 1408 13323 1411
rect 13722 1408 13728 1420
rect 13311 1380 13728 1408
rect 13311 1377 13323 1380
rect 13265 1371 13323 1377
rect 13722 1368 13728 1380
rect 13780 1368 13786 1420
rect 13998 1408 14004 1420
rect 13959 1380 14004 1408
rect 13998 1368 14004 1380
rect 14056 1408 14062 1420
rect 15654 1408 15660 1420
rect 14056 1380 15660 1408
rect 14056 1368 14062 1380
rect 15654 1368 15660 1380
rect 15712 1368 15718 1420
rect 16577 1411 16635 1417
rect 16577 1377 16589 1411
rect 16623 1408 16635 1411
rect 18322 1408 18328 1420
rect 16623 1380 18328 1408
rect 16623 1377 16635 1380
rect 16577 1371 16635 1377
rect 18322 1368 18328 1380
rect 18380 1368 18386 1420
rect 11517 1343 11575 1349
rect 11517 1309 11529 1343
rect 11563 1309 11575 1343
rect 12066 1340 12072 1352
rect 12027 1312 12072 1340
rect 11517 1303 11575 1309
rect 12066 1300 12072 1312
rect 12124 1300 12130 1352
rect 12618 1300 12624 1352
rect 12676 1340 12682 1352
rect 13633 1343 13691 1349
rect 13633 1340 13645 1343
rect 12676 1312 13645 1340
rect 12676 1300 12682 1312
rect 13633 1309 13645 1312
rect 13679 1309 13691 1343
rect 13633 1303 13691 1309
rect 14090 1300 14096 1352
rect 14148 1340 14154 1352
rect 14369 1343 14427 1349
rect 14369 1340 14381 1343
rect 14148 1312 14381 1340
rect 14148 1300 14154 1312
rect 14369 1309 14381 1312
rect 14415 1309 14427 1343
rect 16298 1340 16304 1352
rect 16259 1312 16304 1340
rect 14369 1303 14427 1309
rect 16298 1300 16304 1312
rect 16356 1300 16362 1352
rect 11333 1275 11391 1281
rect 10704 1244 11284 1272
rect 7561 1207 7619 1213
rect 7561 1204 7573 1207
rect 7248 1176 7573 1204
rect 7248 1164 7254 1176
rect 7561 1173 7573 1176
rect 7607 1173 7619 1207
rect 7561 1167 7619 1173
rect 7929 1207 7987 1213
rect 7929 1173 7941 1207
rect 7975 1173 7987 1207
rect 7929 1167 7987 1173
rect 9309 1207 9367 1213
rect 9309 1173 9321 1207
rect 9355 1204 9367 1207
rect 9398 1204 9404 1216
rect 9355 1176 9404 1204
rect 9355 1173 9367 1176
rect 9309 1167 9367 1173
rect 9398 1164 9404 1176
rect 9456 1164 9462 1216
rect 9582 1164 9588 1216
rect 9640 1204 9646 1216
rect 9677 1207 9735 1213
rect 9677 1204 9689 1207
rect 9640 1176 9689 1204
rect 9640 1164 9646 1176
rect 9677 1173 9689 1176
rect 9723 1173 9735 1207
rect 9677 1167 9735 1173
rect 10413 1207 10471 1213
rect 10413 1173 10425 1207
rect 10459 1204 10471 1207
rect 10686 1204 10692 1216
rect 10459 1176 10692 1204
rect 10459 1173 10471 1176
rect 10413 1167 10471 1173
rect 10686 1164 10692 1176
rect 10744 1164 10750 1216
rect 11256 1204 11284 1244
rect 11333 1241 11345 1275
rect 11379 1272 11391 1275
rect 11422 1272 11428 1284
rect 11379 1244 11428 1272
rect 11379 1241 11391 1244
rect 11333 1235 11391 1241
rect 11422 1232 11428 1244
rect 11480 1232 11486 1284
rect 12989 1275 13047 1281
rect 12989 1241 13001 1275
rect 13035 1272 13047 1275
rect 13170 1272 13176 1284
rect 13035 1244 13176 1272
rect 13035 1241 13047 1244
rect 12989 1235 13047 1241
rect 13170 1232 13176 1244
rect 13228 1232 13234 1284
rect 13354 1232 13360 1284
rect 13412 1272 13418 1284
rect 13725 1275 13783 1281
rect 13725 1272 13737 1275
rect 13412 1244 13737 1272
rect 13412 1232 13418 1244
rect 13725 1241 13737 1244
rect 13771 1241 13783 1275
rect 13906 1272 13912 1284
rect 13867 1244 13912 1272
rect 13725 1235 13783 1241
rect 13906 1232 13912 1244
rect 13964 1232 13970 1284
rect 15102 1232 15108 1284
rect 15160 1232 15166 1284
rect 15562 1232 15568 1284
rect 15620 1272 15626 1284
rect 15795 1275 15853 1281
rect 15795 1272 15807 1275
rect 15620 1244 15807 1272
rect 15620 1232 15626 1244
rect 15795 1241 15807 1244
rect 15841 1272 15853 1275
rect 16206 1272 16212 1284
rect 15841 1244 16212 1272
rect 15841 1241 15853 1244
rect 15795 1235 15853 1241
rect 16206 1232 16212 1244
rect 16264 1232 16270 1284
rect 11609 1207 11667 1213
rect 11609 1204 11621 1207
rect 11256 1176 11621 1204
rect 11609 1173 11621 1176
rect 11655 1173 11667 1207
rect 11609 1167 11667 1173
rect 11977 1207 12035 1213
rect 11977 1173 11989 1207
rect 12023 1204 12035 1207
rect 12621 1207 12679 1213
rect 12621 1204 12633 1207
rect 12023 1176 12633 1204
rect 12023 1173 12035 1176
rect 11977 1167 12035 1173
rect 12621 1173 12633 1176
rect 12667 1173 12679 1207
rect 13630 1204 13636 1216
rect 13591 1176 13636 1204
rect 12621 1167 12679 1173
rect 13630 1164 13636 1176
rect 13688 1164 13694 1216
rect 15120 1204 15148 1232
rect 15930 1204 15936 1216
rect 15120 1176 15936 1204
rect 15930 1164 15936 1176
rect 15988 1204 15994 1216
rect 16117 1207 16175 1213
rect 16117 1204 16129 1207
rect 15988 1176 16129 1204
rect 15988 1164 15994 1176
rect 16117 1173 16129 1176
rect 16163 1204 16175 1207
rect 17052 1204 17080 1258
rect 16163 1176 17080 1204
rect 16163 1173 16175 1176
rect 16117 1167 16175 1173
rect 368 1114 18860 1136
rect 368 1062 5028 1114
rect 5080 1062 5092 1114
rect 5144 1062 5156 1114
rect 5208 1062 5220 1114
rect 5272 1062 5284 1114
rect 5336 1062 8128 1114
rect 8180 1062 8192 1114
rect 8244 1062 8256 1114
rect 8308 1062 8320 1114
rect 8372 1062 8384 1114
rect 8436 1062 11228 1114
rect 11280 1062 11292 1114
rect 11344 1062 11356 1114
rect 11408 1062 11420 1114
rect 11472 1062 11484 1114
rect 11536 1062 14328 1114
rect 14380 1062 14392 1114
rect 14444 1062 14456 1114
rect 14508 1062 14520 1114
rect 14572 1062 14584 1114
rect 14636 1062 17428 1114
rect 17480 1062 17492 1114
rect 17544 1062 17556 1114
rect 17608 1062 17620 1114
rect 17672 1062 17684 1114
rect 17736 1062 18860 1114
rect 368 1040 18860 1062
rect 2915 1003 2973 1009
rect 2915 969 2927 1003
rect 2961 1000 2973 1003
rect 7282 1000 7288 1012
rect 2961 972 7144 1000
rect 7243 972 7288 1000
rect 2961 969 2973 972
rect 2915 963 2973 969
rect 3970 892 3976 944
rect 4028 892 4034 944
rect 4706 864 4712 876
rect 4667 836 4712 864
rect 4706 824 4712 836
rect 4764 824 4770 876
rect 5276 873 5304 972
rect 5626 932 5632 944
rect 5552 904 5632 932
rect 5552 873 5580 904
rect 5626 892 5632 904
rect 5684 892 5690 944
rect 5902 892 5908 944
rect 5960 932 5966 944
rect 5960 904 6302 932
rect 5960 892 5966 904
rect 5077 867 5135 873
rect 5077 833 5089 867
rect 5123 833 5135 867
rect 5077 827 5135 833
rect 5261 867 5319 873
rect 5261 833 5273 867
rect 5307 833 5319 867
rect 5261 827 5319 833
rect 5537 867 5595 873
rect 5537 833 5549 867
rect 5583 833 5595 867
rect 7116 864 7144 972
rect 7282 960 7288 972
rect 7340 1000 7346 1012
rect 8018 1000 8024 1012
rect 7340 972 8024 1000
rect 7340 960 7346 972
rect 8018 960 8024 972
rect 8076 1000 8082 1012
rect 8662 1000 8668 1012
rect 8076 972 8156 1000
rect 8623 972 8668 1000
rect 8076 960 8082 972
rect 7837 867 7895 873
rect 7837 864 7849 867
rect 7116 836 7849 864
rect 5537 827 5595 833
rect 7837 833 7849 836
rect 7883 833 7895 867
rect 7837 827 7895 833
rect 2685 799 2743 805
rect 2685 765 2697 799
rect 2731 796 2743 799
rect 3970 796 3976 808
rect 2731 768 3976 796
rect 2731 765 2743 768
rect 2685 759 2743 765
rect 3970 756 3976 768
rect 4028 756 4034 808
rect 4341 799 4399 805
rect 4341 765 4353 799
rect 4387 796 4399 799
rect 4801 799 4859 805
rect 4387 768 4752 796
rect 4387 765 4399 768
rect 4341 759 4399 765
rect 4724 728 4752 768
rect 4801 765 4813 799
rect 4847 796 4859 799
rect 4982 796 4988 808
rect 4847 768 4988 796
rect 4847 765 4859 768
rect 4801 759 4859 765
rect 4982 756 4988 768
rect 5040 756 5046 808
rect 5092 796 5120 827
rect 5810 796 5816 808
rect 5092 768 5396 796
rect 5771 768 5816 796
rect 4893 731 4951 737
rect 4893 728 4905 731
rect 4724 700 4905 728
rect 4893 697 4905 700
rect 4939 697 4951 731
rect 4893 691 4951 697
rect 4985 663 5043 669
rect 4985 629 4997 663
rect 5031 660 5043 663
rect 5166 660 5172 672
rect 5031 632 5172 660
rect 5031 629 5043 632
rect 4985 623 5043 629
rect 5166 620 5172 632
rect 5224 620 5230 672
rect 5368 669 5396 768
rect 5810 756 5816 768
rect 5868 756 5874 808
rect 7852 796 7880 827
rect 7926 824 7932 876
rect 7984 864 7990 876
rect 8128 873 8156 972
rect 8662 960 8668 972
rect 8720 960 8726 1012
rect 9398 1000 9404 1012
rect 9359 972 9404 1000
rect 9398 960 9404 972
rect 9456 960 9462 1012
rect 9490 960 9496 1012
rect 9548 1000 9554 1012
rect 10321 1003 10379 1009
rect 9548 972 9593 1000
rect 9548 960 9554 972
rect 10321 969 10333 1003
rect 10367 1000 10379 1003
rect 10367 972 11192 1000
rect 10367 969 10379 972
rect 10321 963 10379 969
rect 11164 944 11192 972
rect 11606 960 11612 1012
rect 11664 1000 11670 1012
rect 12161 1003 12219 1009
rect 12161 1000 12173 1003
rect 11664 972 12173 1000
rect 11664 960 11670 972
rect 12161 969 12173 972
rect 12207 1000 12219 1003
rect 12618 1000 12624 1012
rect 12207 972 12434 1000
rect 12579 972 12624 1000
rect 12207 969 12219 972
rect 12161 963 12219 969
rect 10686 932 10692 944
rect 10647 904 10692 932
rect 10686 892 10692 904
rect 10744 892 10750 944
rect 11146 892 11152 944
rect 11204 892 11210 944
rect 8021 867 8079 873
rect 8021 864 8033 867
rect 7984 836 8033 864
rect 7984 824 7990 836
rect 8021 833 8033 836
rect 8067 833 8079 867
rect 8021 827 8079 833
rect 8113 867 8171 873
rect 8113 833 8125 867
rect 8159 833 8171 867
rect 8113 827 8171 833
rect 8389 867 8447 873
rect 8389 833 8401 867
rect 8435 833 8447 867
rect 8389 827 8447 833
rect 8941 867 8999 873
rect 8941 833 8953 867
rect 8987 833 8999 867
rect 12406 864 12434 972
rect 12618 960 12624 972
rect 12676 960 12682 1012
rect 13354 1000 13360 1012
rect 13315 972 13360 1000
rect 13354 960 13360 972
rect 13412 960 13418 1012
rect 13633 1003 13691 1009
rect 13633 969 13645 1003
rect 13679 1000 13691 1003
rect 13722 1000 13728 1012
rect 13679 972 13728 1000
rect 13679 969 13691 972
rect 13633 963 13691 969
rect 13722 960 13728 972
rect 13780 960 13786 1012
rect 14645 1003 14703 1009
rect 14645 969 14657 1003
rect 14691 1000 14703 1003
rect 14734 1000 14740 1012
rect 14691 972 14740 1000
rect 14691 969 14703 972
rect 14645 963 14703 969
rect 14734 960 14740 972
rect 14792 960 14798 1012
rect 15102 960 15108 1012
rect 15160 1000 15166 1012
rect 17218 1000 17224 1012
rect 15160 972 15205 1000
rect 17179 972 17224 1000
rect 15160 960 15166 972
rect 17218 960 17224 972
rect 17276 960 17282 1012
rect 18230 1000 18236 1012
rect 18191 972 18236 1000
rect 18230 960 18236 972
rect 18288 960 18294 1012
rect 13446 892 13452 944
rect 13504 932 13510 944
rect 13909 935 13967 941
rect 13909 932 13921 935
rect 13504 904 13921 932
rect 13504 892 13510 904
rect 13909 901 13921 904
rect 13955 901 13967 935
rect 13909 895 13967 901
rect 14826 892 14832 944
rect 14884 932 14890 944
rect 14884 904 14929 932
rect 14884 892 14890 904
rect 15010 892 15016 944
rect 15068 932 15074 944
rect 15068 904 15113 932
rect 15068 892 15074 904
rect 15930 892 15936 944
rect 15988 892 15994 944
rect 17862 892 17868 944
rect 17920 892 17926 944
rect 12526 864 12532 876
rect 12406 836 12532 864
rect 8941 827 8999 833
rect 8404 796 8432 827
rect 8846 796 8852 808
rect 7852 768 8852 796
rect 8846 756 8852 768
rect 8904 756 8910 808
rect 8956 740 8984 827
rect 12526 824 12532 836
rect 12584 824 12590 876
rect 13265 867 13323 873
rect 13265 833 13277 867
rect 13311 864 13323 867
rect 13538 864 13544 876
rect 13311 836 13544 864
rect 13311 833 13323 836
rect 13265 827 13323 833
rect 13538 824 13544 836
rect 13596 824 13602 876
rect 13630 824 13636 876
rect 13688 864 13694 876
rect 13725 867 13783 873
rect 13725 864 13737 867
rect 13688 836 13737 864
rect 13688 824 13694 836
rect 13725 833 13737 836
rect 13771 833 13783 867
rect 13725 827 13783 833
rect 13814 824 13820 876
rect 13872 864 13878 876
rect 13872 836 14228 864
rect 13872 824 13878 836
rect 14200 808 14228 836
rect 14366 824 14372 876
rect 14424 864 14430 876
rect 17586 864 17592 876
rect 14424 862 14872 864
rect 14424 854 14964 862
rect 15089 857 15147 863
rect 15089 854 15101 857
rect 14424 836 15101 854
rect 14424 824 14430 836
rect 14844 834 15101 836
rect 14936 826 15101 834
rect 15089 823 15101 826
rect 15135 823 15147 857
rect 17547 836 17592 864
rect 17586 824 17592 836
rect 17644 824 17650 876
rect 15089 817 15147 823
rect 9306 756 9312 808
rect 9364 796 9370 808
rect 9585 799 9643 805
rect 9585 796 9597 799
rect 9364 768 9597 796
rect 9364 756 9370 768
rect 9585 765 9597 768
rect 9631 765 9643 799
rect 9585 759 9643 765
rect 10413 799 10471 805
rect 10413 765 10425 799
rect 10459 796 10471 799
rect 10778 796 10784 808
rect 10459 768 10784 796
rect 10459 765 10471 768
rect 10413 759 10471 765
rect 10778 756 10784 768
rect 10836 756 10842 808
rect 14182 796 14188 808
rect 14143 768 14188 796
rect 14182 756 14188 768
rect 14240 756 14246 808
rect 14277 799 14335 805
rect 14277 765 14289 799
rect 14323 796 14335 799
rect 14734 796 14740 808
rect 14323 768 14740 796
rect 14323 765 14335 768
rect 14277 759 14335 765
rect 14734 756 14740 768
rect 14792 756 14798 808
rect 15197 799 15255 805
rect 15197 765 15209 799
rect 15243 765 15255 799
rect 15470 796 15476 808
rect 15431 768 15476 796
rect 15197 759 15255 765
rect 7926 688 7932 740
rect 7984 728 7990 740
rect 8938 728 8944 740
rect 7984 700 8944 728
rect 7984 688 7990 700
rect 8938 688 8944 700
rect 8996 688 9002 740
rect 5353 663 5411 669
rect 5353 629 5365 663
rect 5399 660 5411 663
rect 5442 660 5448 672
rect 5399 632 5448 660
rect 5399 629 5411 632
rect 5353 623 5411 629
rect 5442 620 5448 632
rect 5500 620 5506 672
rect 8021 663 8079 669
rect 8021 629 8033 663
rect 8067 660 8079 663
rect 8110 660 8116 672
rect 8067 632 8116 660
rect 8067 629 8079 632
rect 8021 623 8079 629
rect 8110 620 8116 632
rect 8168 620 8174 672
rect 9030 660 9036 672
rect 8991 632 9036 660
rect 9030 620 9036 632
rect 9088 620 9094 672
rect 14001 663 14059 669
rect 14001 629 14013 663
rect 14047 660 14059 663
rect 14090 660 14096 672
rect 14047 632 14096 660
rect 14047 629 14059 632
rect 14001 623 14059 629
rect 14090 620 14096 632
rect 14148 620 14154 672
rect 15212 660 15240 759
rect 15470 756 15476 768
rect 15528 756 15534 808
rect 16666 756 16672 808
rect 16724 796 16730 808
rect 17880 805 17908 892
rect 18049 867 18107 873
rect 18049 833 18061 867
rect 18095 833 18107 867
rect 18049 827 18107 833
rect 17681 799 17739 805
rect 17681 796 17693 799
rect 16724 768 17693 796
rect 16724 756 16730 768
rect 17681 765 17693 768
rect 17727 765 17739 799
rect 17681 759 17739 765
rect 17865 799 17923 805
rect 17865 765 17877 799
rect 17911 765 17923 799
rect 17865 759 17923 765
rect 16942 728 16948 740
rect 16903 700 16948 728
rect 16942 688 16948 700
rect 17000 728 17006 740
rect 18064 728 18092 827
rect 17000 700 18092 728
rect 17000 688 17006 700
rect 15654 660 15660 672
rect 15212 632 15660 660
rect 15654 620 15660 632
rect 15712 620 15718 672
rect 368 570 18860 592
rect 368 518 3478 570
rect 3530 518 3542 570
rect 3594 518 3606 570
rect 3658 518 3670 570
rect 3722 518 3734 570
rect 3786 518 6578 570
rect 6630 518 6642 570
rect 6694 518 6706 570
rect 6758 518 6770 570
rect 6822 518 6834 570
rect 6886 518 9678 570
rect 9730 518 9742 570
rect 9794 518 9806 570
rect 9858 518 9870 570
rect 9922 518 9934 570
rect 9986 518 12778 570
rect 12830 518 12842 570
rect 12894 518 12906 570
rect 12958 518 12970 570
rect 13022 518 13034 570
rect 13086 518 15878 570
rect 15930 518 15942 570
rect 15994 518 16006 570
rect 16058 518 16070 570
rect 16122 518 16134 570
rect 16186 518 18860 570
rect 368 496 18860 518
rect 4982 456 4988 468
rect 4943 428 4988 456
rect 4982 416 4988 428
rect 5040 416 5046 468
rect 5810 456 5816 468
rect 5771 428 5816 456
rect 5810 416 5816 428
rect 5868 416 5874 468
rect 5905 459 5963 465
rect 5905 425 5917 459
rect 5951 456 5963 459
rect 6362 456 6368 468
rect 5951 428 6368 456
rect 5951 425 5963 428
rect 5905 419 5963 425
rect 4614 348 4620 400
rect 4672 388 4678 400
rect 5166 388 5172 400
rect 4672 360 5172 388
rect 4672 348 4678 360
rect 4908 261 4936 360
rect 5166 348 5172 360
rect 5224 388 5230 400
rect 5920 388 5948 419
rect 6362 416 6368 428
rect 6420 416 6426 468
rect 6454 416 6460 468
rect 6512 456 6518 468
rect 6549 459 6607 465
rect 6549 456 6561 459
rect 6512 428 6561 456
rect 6512 416 6518 428
rect 6549 425 6561 428
rect 6595 425 6607 459
rect 6549 419 6607 425
rect 8389 459 8447 465
rect 8389 425 8401 459
rect 8435 456 8447 459
rect 8478 456 8484 468
rect 8435 428 8484 456
rect 8435 425 8447 428
rect 8389 419 8447 425
rect 8478 416 8484 428
rect 8536 416 8542 468
rect 12989 459 13047 465
rect 12989 425 13001 459
rect 13035 456 13047 459
rect 13170 456 13176 468
rect 13035 428 13176 456
rect 13035 425 13047 428
rect 12989 419 13047 425
rect 13170 416 13176 428
rect 13228 416 13234 468
rect 15013 459 15071 465
rect 15013 425 15025 459
rect 15059 456 15071 459
rect 15194 456 15200 468
rect 15059 428 15200 456
rect 15059 425 15071 428
rect 15013 419 15071 425
rect 15194 416 15200 428
rect 15252 416 15258 468
rect 15470 416 15476 468
rect 15528 456 15534 468
rect 15749 459 15807 465
rect 15749 456 15761 459
rect 15528 428 15761 456
rect 15528 416 15534 428
rect 15749 425 15761 428
rect 15795 425 15807 459
rect 15749 419 15807 425
rect 17586 416 17592 468
rect 17644 456 17650 468
rect 17681 459 17739 465
rect 17681 456 17693 459
rect 17644 428 17693 456
rect 17644 416 17650 428
rect 17681 425 17693 428
rect 17727 425 17739 459
rect 18046 456 18052 468
rect 18007 428 18052 456
rect 17681 419 17739 425
rect 18046 416 18052 428
rect 18104 416 18110 468
rect 18506 456 18512 468
rect 18467 428 18512 456
rect 18506 416 18512 428
rect 18564 416 18570 468
rect 5224 360 5948 388
rect 9401 391 9459 397
rect 5224 348 5230 360
rect 9401 357 9413 391
rect 9447 388 9459 391
rect 9582 388 9588 400
rect 9447 360 9588 388
rect 9447 357 9459 360
rect 9401 351 9459 357
rect 9582 348 9588 360
rect 9640 348 9646 400
rect 13906 348 13912 400
rect 13964 388 13970 400
rect 14918 388 14924 400
rect 13964 360 14924 388
rect 13964 348 13970 360
rect 14918 348 14924 360
rect 14976 388 14982 400
rect 16942 388 16948 400
rect 14976 360 16948 388
rect 14976 348 14982 360
rect 16942 348 16948 360
rect 17000 388 17006 400
rect 17000 360 17356 388
rect 17000 348 17006 360
rect 5721 323 5779 329
rect 5721 289 5733 323
rect 5767 320 5779 323
rect 6086 320 6092 332
rect 5767 292 6092 320
rect 5767 289 5779 292
rect 5721 283 5779 289
rect 6086 280 6092 292
rect 6144 280 6150 332
rect 6454 280 6460 332
rect 6512 320 6518 332
rect 7926 320 7932 332
rect 6512 292 7932 320
rect 6512 280 6518 292
rect 7926 280 7932 292
rect 7984 280 7990 332
rect 8110 320 8116 332
rect 8071 292 8116 320
rect 8110 280 8116 292
rect 8168 280 8174 332
rect 8938 320 8944 332
rect 8899 292 8944 320
rect 8938 280 8944 292
rect 8996 280 9002 332
rect 12713 323 12771 329
rect 12713 289 12725 323
rect 12759 320 12771 323
rect 13265 323 13323 329
rect 13265 320 13277 323
rect 12759 292 13277 320
rect 12759 289 12771 292
rect 12713 283 12771 289
rect 13265 289 13277 292
rect 13311 289 13323 323
rect 15102 320 15108 332
rect 15063 292 15108 320
rect 13265 283 13323 289
rect 15102 280 15108 292
rect 15160 280 15166 332
rect 15286 280 15292 332
rect 15344 320 15350 332
rect 17328 329 17356 360
rect 15473 323 15531 329
rect 15473 320 15485 323
rect 15344 292 15485 320
rect 15344 280 15350 292
rect 15473 289 15485 292
rect 15519 289 15531 323
rect 15473 283 15531 289
rect 17313 323 17371 329
rect 17313 289 17325 323
rect 17359 289 17371 323
rect 17313 283 17371 289
rect 4893 255 4951 261
rect 4893 221 4905 255
rect 4939 221 4951 255
rect 5074 252 5080 264
rect 5035 224 5080 252
rect 4893 215 4951 221
rect 5074 212 5080 224
rect 5132 212 5138 264
rect 5445 255 5503 261
rect 5445 221 5457 255
rect 5491 252 5503 255
rect 5902 252 5908 264
rect 5491 224 5908 252
rect 5491 221 5503 224
rect 5445 215 5503 221
rect 5902 212 5908 224
rect 5960 212 5966 264
rect 5997 255 6055 261
rect 5997 221 6009 255
rect 6043 252 6055 255
rect 6733 255 6791 261
rect 6733 252 6745 255
rect 6043 224 6745 252
rect 6043 221 6055 224
rect 5997 215 6055 221
rect 6733 221 6745 224
rect 6779 252 6791 255
rect 6822 252 6828 264
rect 6779 224 6828 252
rect 6779 221 6791 224
rect 6733 215 6791 221
rect 6822 212 6828 224
rect 6880 212 6886 264
rect 8018 252 8024 264
rect 7979 224 8024 252
rect 8018 212 8024 224
rect 8076 212 8082 264
rect 8846 212 8852 264
rect 8904 252 8910 264
rect 9033 255 9091 261
rect 9033 252 9045 255
rect 8904 224 9045 252
rect 8904 212 8910 224
rect 9033 221 9045 224
rect 9079 221 9091 255
rect 9033 215 9091 221
rect 12526 212 12532 264
rect 12584 252 12590 264
rect 12621 255 12679 261
rect 12621 252 12633 255
rect 12584 224 12633 252
rect 12584 212 12590 224
rect 12621 221 12633 224
rect 12667 221 12679 255
rect 12621 215 12679 221
rect 13173 255 13231 261
rect 13173 221 13185 255
rect 13219 221 13231 255
rect 13173 215 13231 221
rect 13357 255 13415 261
rect 13357 221 13369 255
rect 13403 252 13415 255
rect 13906 252 13912 264
rect 13403 224 13912 252
rect 13403 221 13415 224
rect 13357 215 13415 221
rect 4798 144 4804 196
rect 4856 184 4862 196
rect 6454 184 6460 196
rect 4856 156 6460 184
rect 4856 144 4862 156
rect 6454 144 6460 156
rect 6512 144 6518 196
rect 6641 187 6699 193
rect 6641 153 6653 187
rect 6687 153 6699 187
rect 13188 184 13216 215
rect 13906 212 13912 224
rect 13964 212 13970 264
rect 14182 212 14188 264
rect 14240 252 14246 264
rect 15565 255 15623 261
rect 15565 252 15577 255
rect 14240 224 15577 252
rect 14240 212 14246 224
rect 15565 221 15577 224
rect 15611 221 15623 255
rect 15565 215 15623 221
rect 16206 212 16212 264
rect 16264 252 16270 264
rect 17405 255 17463 261
rect 17405 252 17417 255
rect 16264 224 17417 252
rect 16264 212 16270 224
rect 17405 221 17417 224
rect 17451 221 17463 255
rect 17405 215 17463 221
rect 18233 255 18291 261
rect 18233 221 18245 255
rect 18279 252 18291 255
rect 18506 252 18512 264
rect 18279 224 18512 252
rect 18279 221 18291 224
rect 18233 215 18291 221
rect 18506 212 18512 224
rect 18564 212 18570 264
rect 13538 184 13544 196
rect 13188 156 13544 184
rect 6641 147 6699 153
rect 5442 76 5448 128
rect 5500 116 5506 128
rect 6656 116 6684 147
rect 13538 144 13544 156
rect 13596 144 13602 196
rect 5500 88 6684 116
rect 5500 76 5506 88
rect 368 26 18860 48
rect 368 -26 5028 26
rect 5080 -26 5092 26
rect 5144 -26 5156 26
rect 5208 -26 5220 26
rect 5272 -26 5284 26
rect 5336 -26 8128 26
rect 8180 -26 8192 26
rect 8244 -26 8256 26
rect 8308 -26 8320 26
rect 8372 -26 8384 26
rect 8436 -26 11228 26
rect 11280 -26 11292 26
rect 11344 -26 11356 26
rect 11408 -26 11420 26
rect 11472 -26 11484 26
rect 11536 -26 14328 26
rect 14380 -26 14392 26
rect 14444 -26 14456 26
rect 14508 -26 14520 26
rect 14572 -26 14584 26
rect 14636 -26 17428 26
rect 17480 -26 17492 26
rect 17544 -26 17556 26
rect 17608 -26 17620 26
rect 17672 -26 17684 26
rect 17736 -26 18860 26
rect 368 -48 18860 -26
<< via1 >>
rect 5028 10854 5080 10906
rect 5092 10854 5144 10906
rect 5156 10854 5208 10906
rect 5220 10854 5272 10906
rect 5284 10854 5336 10906
rect 8128 10854 8180 10906
rect 8192 10854 8244 10906
rect 8256 10854 8308 10906
rect 8320 10854 8372 10906
rect 8384 10854 8436 10906
rect 11228 10854 11280 10906
rect 11292 10854 11344 10906
rect 11356 10854 11408 10906
rect 11420 10854 11472 10906
rect 11484 10854 11536 10906
rect 14328 10854 14380 10906
rect 14392 10854 14444 10906
rect 14456 10854 14508 10906
rect 14520 10854 14572 10906
rect 14584 10854 14636 10906
rect 17428 10854 17480 10906
rect 17492 10854 17544 10906
rect 17556 10854 17608 10906
rect 17620 10854 17672 10906
rect 17684 10854 17736 10906
rect 6828 10795 6880 10804
rect 6828 10761 6837 10795
rect 6837 10761 6871 10795
rect 6871 10761 6880 10795
rect 6828 10752 6880 10761
rect 664 10616 716 10668
rect 2412 10616 2464 10668
rect 3056 10616 3108 10668
rect 5264 10659 5316 10668
rect 5264 10625 5273 10659
rect 5273 10625 5307 10659
rect 5307 10625 5316 10659
rect 5264 10616 5316 10625
rect 5448 10659 5500 10668
rect 5448 10625 5457 10659
rect 5457 10625 5491 10659
rect 5491 10625 5500 10659
rect 5448 10616 5500 10625
rect 9956 10752 10008 10804
rect 12900 10752 12952 10804
rect 3240 10548 3292 10600
rect 8760 10616 8812 10668
rect 2688 10480 2740 10532
rect 8576 10548 8628 10600
rect 8484 10480 8536 10532
rect 11152 10616 11204 10668
rect 12532 10684 12584 10736
rect 13176 10616 13228 10668
rect 18788 10752 18840 10804
rect 12440 10548 12492 10600
rect 13268 10548 13320 10600
rect 18052 10659 18104 10668
rect 18052 10625 18061 10659
rect 18061 10625 18095 10659
rect 18095 10625 18104 10659
rect 18052 10616 18104 10625
rect 2044 10412 2096 10464
rect 2596 10412 2648 10464
rect 2964 10455 3016 10464
rect 2964 10421 2973 10455
rect 2973 10421 3007 10455
rect 3007 10421 3016 10455
rect 2964 10412 3016 10421
rect 4436 10412 4488 10464
rect 7288 10412 7340 10464
rect 8576 10455 8628 10464
rect 8576 10421 8585 10455
rect 8585 10421 8619 10455
rect 8619 10421 8628 10455
rect 8576 10412 8628 10421
rect 9128 10412 9180 10464
rect 11980 10412 12032 10464
rect 13176 10455 13228 10464
rect 13176 10421 13185 10455
rect 13185 10421 13219 10455
rect 13219 10421 13228 10455
rect 13176 10412 13228 10421
rect 14004 10455 14056 10464
rect 14004 10421 14013 10455
rect 14013 10421 14047 10455
rect 14047 10421 14056 10455
rect 14004 10412 14056 10421
rect 15292 10412 15344 10464
rect 3478 10310 3530 10362
rect 3542 10310 3594 10362
rect 3606 10310 3658 10362
rect 3670 10310 3722 10362
rect 3734 10310 3786 10362
rect 6578 10310 6630 10362
rect 6642 10310 6694 10362
rect 6706 10310 6758 10362
rect 6770 10310 6822 10362
rect 6834 10310 6886 10362
rect 9678 10310 9730 10362
rect 9742 10310 9794 10362
rect 9806 10310 9858 10362
rect 9870 10310 9922 10362
rect 9934 10310 9986 10362
rect 12778 10310 12830 10362
rect 12842 10310 12894 10362
rect 12906 10310 12958 10362
rect 12970 10310 13022 10362
rect 13034 10310 13086 10362
rect 15878 10310 15930 10362
rect 15942 10310 15994 10362
rect 16006 10310 16058 10362
rect 16070 10310 16122 10362
rect 16134 10310 16186 10362
rect 2688 10208 2740 10260
rect 4252 10208 4304 10260
rect 5264 10140 5316 10192
rect 8484 10208 8536 10260
rect 8760 10208 8812 10260
rect 12624 10208 12676 10260
rect 18052 10208 18104 10260
rect 1676 10115 1728 10124
rect 1676 10081 1685 10115
rect 1685 10081 1719 10115
rect 1719 10081 1728 10115
rect 1676 10072 1728 10081
rect 2044 10115 2096 10124
rect 2044 10081 2053 10115
rect 2053 10081 2087 10115
rect 2087 10081 2096 10115
rect 2044 10072 2096 10081
rect 2964 10072 3016 10124
rect 3148 10072 3200 10124
rect 4436 10115 4488 10124
rect 4436 10081 4445 10115
rect 4445 10081 4479 10115
rect 4479 10081 4488 10115
rect 4436 10072 4488 10081
rect 5540 10072 5592 10124
rect 2504 10004 2556 10056
rect 2780 9936 2832 9988
rect 940 9868 992 9920
rect 2412 9868 2464 9920
rect 7196 10047 7248 10056
rect 3792 9868 3844 9920
rect 5448 9936 5500 9988
rect 7196 10013 7205 10047
rect 7205 10013 7239 10047
rect 7239 10013 7248 10047
rect 7196 10004 7248 10013
rect 7288 10004 7340 10056
rect 11980 10072 12032 10124
rect 11060 10004 11112 10056
rect 13176 10072 13228 10124
rect 11612 9936 11664 9988
rect 11980 9936 12032 9988
rect 5356 9911 5408 9920
rect 5356 9877 5365 9911
rect 5365 9877 5399 9911
rect 5399 9877 5408 9911
rect 5356 9868 5408 9877
rect 6276 9911 6328 9920
rect 6276 9877 6285 9911
rect 6285 9877 6319 9911
rect 6319 9877 6328 9911
rect 6276 9868 6328 9877
rect 12440 9868 12492 9920
rect 12808 9868 12860 9920
rect 14096 10004 14148 10056
rect 15292 9868 15344 9920
rect 5028 9766 5080 9818
rect 5092 9766 5144 9818
rect 5156 9766 5208 9818
rect 5220 9766 5272 9818
rect 5284 9766 5336 9818
rect 8128 9766 8180 9818
rect 8192 9766 8244 9818
rect 8256 9766 8308 9818
rect 8320 9766 8372 9818
rect 8384 9766 8436 9818
rect 11228 9766 11280 9818
rect 11292 9766 11344 9818
rect 11356 9766 11408 9818
rect 11420 9766 11472 9818
rect 11484 9766 11536 9818
rect 14328 9766 14380 9818
rect 14392 9766 14444 9818
rect 14456 9766 14508 9818
rect 14520 9766 14572 9818
rect 14584 9766 14636 9818
rect 17428 9766 17480 9818
rect 17492 9766 17544 9818
rect 17556 9766 17608 9818
rect 17620 9766 17672 9818
rect 17684 9766 17736 9818
rect 1676 9664 1728 9716
rect 3240 9707 3292 9716
rect 940 9639 992 9648
rect 940 9605 949 9639
rect 949 9605 983 9639
rect 983 9605 992 9639
rect 940 9596 992 9605
rect 2596 9596 2648 9648
rect 2964 9639 3016 9648
rect 664 9571 716 9580
rect 664 9537 673 9571
rect 673 9537 707 9571
rect 707 9537 716 9571
rect 664 9528 716 9537
rect 2504 9571 2556 9580
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 2504 9528 2556 9537
rect 2964 9605 2973 9639
rect 2973 9605 3007 9639
rect 3007 9605 3016 9639
rect 2964 9596 3016 9605
rect 3240 9673 3249 9707
rect 3249 9673 3283 9707
rect 3283 9673 3292 9707
rect 3240 9664 3292 9673
rect 6276 9664 6328 9716
rect 11152 9664 11204 9716
rect 14096 9664 14148 9716
rect 5264 9596 5316 9648
rect 5540 9596 5592 9648
rect 12624 9639 12676 9648
rect 12624 9605 12633 9639
rect 12633 9605 12667 9639
rect 12667 9605 12676 9639
rect 12624 9596 12676 9605
rect 14188 9596 14240 9648
rect 15568 9596 15620 9648
rect 3148 9571 3200 9580
rect 2412 9503 2464 9512
rect 2412 9469 2421 9503
rect 2421 9469 2455 9503
rect 2455 9469 2464 9503
rect 2412 9460 2464 9469
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 3240 9571 3292 9580
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 3792 9571 3844 9580
rect 3792 9537 3801 9571
rect 3801 9537 3835 9571
rect 3835 9537 3844 9571
rect 3792 9528 3844 9537
rect 2504 9392 2556 9444
rect 2688 9392 2740 9444
rect 3240 9392 3292 9444
rect 4620 9460 4672 9512
rect 6000 9528 6052 9580
rect 6368 9528 6420 9580
rect 8760 9571 8812 9580
rect 8760 9537 8794 9571
rect 8794 9537 8812 9571
rect 8760 9528 8812 9537
rect 2872 9324 2924 9376
rect 3056 9324 3108 9376
rect 4068 9367 4120 9376
rect 4068 9333 4077 9367
rect 4077 9333 4111 9367
rect 4111 9333 4120 9367
rect 4068 9324 4120 9333
rect 5448 9392 5500 9444
rect 10324 9460 10376 9512
rect 11612 9528 11664 9580
rect 10784 9503 10836 9512
rect 10784 9469 10793 9503
rect 10793 9469 10827 9503
rect 10827 9469 10836 9503
rect 10784 9460 10836 9469
rect 12532 9528 12584 9580
rect 13084 9528 13136 9580
rect 18696 9528 18748 9580
rect 6276 9324 6328 9376
rect 6460 9324 6512 9376
rect 7104 9367 7156 9376
rect 7104 9333 7113 9367
rect 7113 9333 7147 9367
rect 7147 9333 7156 9367
rect 7104 9324 7156 9333
rect 10508 9324 10560 9376
rect 14004 9460 14056 9512
rect 14832 9503 14884 9512
rect 14832 9469 14841 9503
rect 14841 9469 14875 9503
rect 14875 9469 14884 9503
rect 14832 9460 14884 9469
rect 16580 9503 16632 9512
rect 16580 9469 16589 9503
rect 16589 9469 16623 9503
rect 16623 9469 16632 9503
rect 16580 9460 16632 9469
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 12808 9392 12860 9444
rect 14096 9324 14148 9376
rect 14372 9324 14424 9376
rect 3478 9222 3530 9274
rect 3542 9222 3594 9274
rect 3606 9222 3658 9274
rect 3670 9222 3722 9274
rect 3734 9222 3786 9274
rect 6578 9222 6630 9274
rect 6642 9222 6694 9274
rect 6706 9222 6758 9274
rect 6770 9222 6822 9274
rect 6834 9222 6886 9274
rect 9678 9222 9730 9274
rect 9742 9222 9794 9274
rect 9806 9222 9858 9274
rect 9870 9222 9922 9274
rect 9934 9222 9986 9274
rect 12778 9222 12830 9274
rect 12842 9222 12894 9274
rect 12906 9222 12958 9274
rect 12970 9222 13022 9274
rect 13034 9222 13086 9274
rect 15878 9222 15930 9274
rect 15942 9222 15994 9274
rect 16006 9222 16058 9274
rect 16070 9222 16122 9274
rect 16134 9222 16186 9274
rect 1400 9120 1452 9172
rect 4620 9120 4672 9172
rect 9588 9120 9640 9172
rect 1308 8984 1360 9036
rect 1492 9052 1544 9104
rect 2504 9052 2556 9104
rect 10784 9120 10836 9172
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 2780 8984 2832 9036
rect 3148 8984 3200 9036
rect 6276 8984 6328 9036
rect 10140 8984 10192 9036
rect 11060 8984 11112 9036
rect 14832 9120 14884 9172
rect 16580 9120 16632 9172
rect 14096 9027 14148 9036
rect 14096 8993 14105 9027
rect 14105 8993 14139 9027
rect 14139 8993 14148 9027
rect 14096 8984 14148 8993
rect 16856 8984 16908 9036
rect 1216 8823 1268 8832
rect 1216 8789 1225 8823
rect 1225 8789 1259 8823
rect 1259 8789 1268 8823
rect 1216 8780 1268 8789
rect 4160 8916 4212 8968
rect 4896 8916 4948 8968
rect 6460 8916 6512 8968
rect 11152 8916 11204 8968
rect 16396 8959 16448 8968
rect 16396 8925 16405 8959
rect 16405 8925 16439 8959
rect 16439 8925 16448 8959
rect 16396 8916 16448 8925
rect 2872 8891 2924 8900
rect 2872 8857 2881 8891
rect 2881 8857 2915 8891
rect 2915 8857 2924 8891
rect 2872 8848 2924 8857
rect 3976 8848 4028 8900
rect 7104 8848 7156 8900
rect 9128 8891 9180 8900
rect 3240 8823 3292 8832
rect 3240 8789 3249 8823
rect 3249 8789 3283 8823
rect 3283 8789 3292 8823
rect 3240 8780 3292 8789
rect 3332 8780 3384 8832
rect 6368 8780 6420 8832
rect 8852 8780 8904 8832
rect 9128 8857 9137 8891
rect 9137 8857 9171 8891
rect 9171 8857 9180 8891
rect 9128 8848 9180 8857
rect 9220 8780 9272 8832
rect 9312 8780 9364 8832
rect 11612 8848 11664 8900
rect 12072 8848 12124 8900
rect 14372 8891 14424 8900
rect 12164 8780 12216 8832
rect 14372 8857 14381 8891
rect 14381 8857 14415 8891
rect 14415 8857 14424 8891
rect 14372 8848 14424 8857
rect 14188 8780 14240 8832
rect 17132 8848 17184 8900
rect 18144 8823 18196 8832
rect 18144 8789 18153 8823
rect 18153 8789 18187 8823
rect 18187 8789 18196 8823
rect 18144 8780 18196 8789
rect 5028 8678 5080 8730
rect 5092 8678 5144 8730
rect 5156 8678 5208 8730
rect 5220 8678 5272 8730
rect 5284 8678 5336 8730
rect 8128 8678 8180 8730
rect 8192 8678 8244 8730
rect 8256 8678 8308 8730
rect 8320 8678 8372 8730
rect 8384 8678 8436 8730
rect 11228 8678 11280 8730
rect 11292 8678 11344 8730
rect 11356 8678 11408 8730
rect 11420 8678 11472 8730
rect 11484 8678 11536 8730
rect 14328 8678 14380 8730
rect 14392 8678 14444 8730
rect 14456 8678 14508 8730
rect 14520 8678 14572 8730
rect 14584 8678 14636 8730
rect 17428 8678 17480 8730
rect 17492 8678 17544 8730
rect 17556 8678 17608 8730
rect 17620 8678 17672 8730
rect 17684 8678 17736 8730
rect 1308 8576 1360 8628
rect 3240 8576 3292 8628
rect 1216 8508 1268 8560
rect 2504 8508 2556 8560
rect 664 8483 716 8492
rect 664 8449 673 8483
rect 673 8449 707 8483
rect 707 8449 716 8483
rect 664 8440 716 8449
rect 3056 8483 3108 8492
rect 2780 8372 2832 8424
rect 3056 8449 3065 8483
rect 3065 8449 3099 8483
rect 3099 8449 3108 8483
rect 3056 8440 3108 8449
rect 3332 8440 3384 8492
rect 5448 8576 5500 8628
rect 4896 8508 4948 8560
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 4344 8415 4396 8424
rect 4344 8381 4353 8415
rect 4353 8381 4387 8415
rect 4387 8381 4396 8415
rect 6184 8505 6236 8526
rect 6184 8474 6191 8505
rect 6191 8474 6225 8505
rect 6225 8474 6236 8505
rect 8392 8508 8444 8560
rect 8576 8508 8628 8560
rect 9312 8576 9364 8628
rect 4344 8372 4396 8381
rect 2872 8304 2924 8356
rect 4804 8279 4856 8288
rect 4804 8245 4813 8279
rect 4813 8245 4847 8279
rect 4847 8245 4856 8279
rect 4804 8236 4856 8245
rect 7564 8440 7616 8492
rect 8484 8440 8536 8492
rect 8852 8483 8904 8492
rect 8852 8449 8861 8483
rect 8861 8449 8895 8483
rect 8895 8449 8904 8483
rect 8852 8440 8904 8449
rect 9220 8440 9272 8492
rect 7104 8304 7156 8356
rect 9772 8440 9824 8492
rect 10048 8372 10100 8424
rect 11612 8576 11664 8628
rect 14096 8508 14148 8560
rect 10416 8483 10468 8492
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 10784 8440 10836 8492
rect 11244 8440 11296 8492
rect 13820 8483 13872 8492
rect 15568 8508 15620 8560
rect 16396 8576 16448 8628
rect 18144 8508 18196 8560
rect 13820 8449 13838 8483
rect 13838 8449 13872 8483
rect 13820 8440 13872 8449
rect 11612 8372 11664 8424
rect 11888 8372 11940 8424
rect 6920 8236 6972 8288
rect 8208 8236 8260 8288
rect 10508 8279 10560 8288
rect 10508 8245 10517 8279
rect 10517 8245 10551 8279
rect 10551 8245 10560 8279
rect 10508 8236 10560 8245
rect 10784 8236 10836 8288
rect 10968 8236 11020 8288
rect 11336 8236 11388 8288
rect 11796 8236 11848 8288
rect 12072 8236 12124 8288
rect 13452 8236 13504 8288
rect 17132 8304 17184 8356
rect 18604 8304 18656 8356
rect 14188 8236 14240 8288
rect 15384 8236 15436 8288
rect 16856 8236 16908 8288
rect 3478 8134 3530 8186
rect 3542 8134 3594 8186
rect 3606 8134 3658 8186
rect 3670 8134 3722 8186
rect 3734 8134 3786 8186
rect 6578 8134 6630 8186
rect 6642 8134 6694 8186
rect 6706 8134 6758 8186
rect 6770 8134 6822 8186
rect 6834 8134 6886 8186
rect 9678 8134 9730 8186
rect 9742 8134 9794 8186
rect 9806 8134 9858 8186
rect 9870 8134 9922 8186
rect 9934 8134 9986 8186
rect 12778 8134 12830 8186
rect 12842 8134 12894 8186
rect 12906 8134 12958 8186
rect 12970 8134 13022 8186
rect 13034 8134 13086 8186
rect 15878 8134 15930 8186
rect 15942 8134 15994 8186
rect 16006 8134 16058 8186
rect 16070 8134 16122 8186
rect 16134 8134 16186 8186
rect 3056 8032 3108 8084
rect 4896 8075 4948 8084
rect 4896 8041 4905 8075
rect 4905 8041 4939 8075
rect 4939 8041 4948 8075
rect 4896 8032 4948 8041
rect 6000 8032 6052 8084
rect 6368 8032 6420 8084
rect 4160 7896 4212 7948
rect 4712 7939 4764 7948
rect 1492 7828 1544 7880
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 2596 7871 2648 7880
rect 2596 7837 2605 7871
rect 2605 7837 2639 7871
rect 2639 7837 2648 7871
rect 2596 7828 2648 7837
rect 3148 7828 3200 7880
rect 3332 7828 3384 7880
rect 4712 7905 4721 7939
rect 4721 7905 4755 7939
rect 4755 7905 4764 7939
rect 4712 7896 4764 7905
rect 6828 7964 6880 8016
rect 9496 8032 9548 8084
rect 10968 8032 11020 8084
rect 9772 7964 9824 8016
rect 10416 7964 10468 8016
rect 4804 7828 4856 7880
rect 2688 7760 2740 7812
rect 4344 7760 4396 7812
rect 6368 7828 6420 7880
rect 6828 7871 6880 7880
rect 6828 7837 6837 7871
rect 6837 7837 6871 7871
rect 6871 7837 6880 7871
rect 6828 7828 6880 7837
rect 7104 7896 7156 7948
rect 9588 7896 9640 7948
rect 18512 8032 18564 8084
rect 14096 7964 14148 8016
rect 11152 7896 11204 7948
rect 13452 7896 13504 7948
rect 14740 7939 14792 7948
rect 14740 7905 14749 7939
rect 14749 7905 14783 7939
rect 14783 7905 14792 7939
rect 14740 7896 14792 7905
rect 14924 7896 14976 7948
rect 17040 7896 17092 7948
rect 11060 7871 11112 7880
rect 11060 7837 11069 7871
rect 11069 7837 11103 7871
rect 11103 7837 11112 7871
rect 11060 7828 11112 7837
rect 11612 7871 11664 7880
rect 11612 7837 11621 7871
rect 11621 7837 11655 7871
rect 11655 7837 11664 7871
rect 11612 7828 11664 7837
rect 12808 7828 12860 7880
rect 14004 7871 14056 7880
rect 14004 7837 14013 7871
rect 14013 7837 14047 7871
rect 14047 7837 14056 7871
rect 14004 7828 14056 7837
rect 14188 7871 14240 7880
rect 14188 7837 14197 7871
rect 14197 7837 14231 7871
rect 14231 7837 14240 7871
rect 14188 7828 14240 7837
rect 5908 7803 5960 7812
rect 5908 7769 5917 7803
rect 5917 7769 5951 7803
rect 5951 7769 5960 7803
rect 5908 7760 5960 7769
rect 6460 7803 6512 7812
rect 6460 7769 6469 7803
rect 6469 7769 6503 7803
rect 6503 7769 6512 7803
rect 6460 7760 6512 7769
rect 2412 7692 2464 7744
rect 5540 7692 5592 7744
rect 8208 7760 8260 7812
rect 8484 7692 8536 7744
rect 9128 7692 9180 7744
rect 12348 7760 12400 7812
rect 13452 7803 13504 7812
rect 13452 7769 13461 7803
rect 13461 7769 13495 7803
rect 13495 7769 13504 7803
rect 13452 7760 13504 7769
rect 15384 7828 15436 7880
rect 13728 7735 13780 7744
rect 13728 7701 13737 7735
rect 13737 7701 13771 7735
rect 13771 7701 13780 7735
rect 13728 7692 13780 7701
rect 16396 7760 16448 7812
rect 15200 7692 15252 7744
rect 16120 7692 16172 7744
rect 17132 7760 17184 7812
rect 17868 7760 17920 7812
rect 5028 7590 5080 7642
rect 5092 7590 5144 7642
rect 5156 7590 5208 7642
rect 5220 7590 5272 7642
rect 5284 7590 5336 7642
rect 8128 7590 8180 7642
rect 8192 7590 8244 7642
rect 8256 7590 8308 7642
rect 8320 7590 8372 7642
rect 8384 7590 8436 7642
rect 11228 7590 11280 7642
rect 11292 7590 11344 7642
rect 11356 7590 11408 7642
rect 11420 7590 11472 7642
rect 11484 7590 11536 7642
rect 14328 7590 14380 7642
rect 14392 7590 14444 7642
rect 14456 7590 14508 7642
rect 14520 7590 14572 7642
rect 14584 7590 14636 7642
rect 17428 7590 17480 7642
rect 17492 7590 17544 7642
rect 17556 7590 17608 7642
rect 17620 7590 17672 7642
rect 17684 7590 17736 7642
rect 2228 7488 2280 7540
rect 2688 7488 2740 7540
rect 4160 7488 4212 7540
rect 2412 7420 2464 7472
rect 6184 7488 6236 7540
rect 6828 7488 6880 7540
rect 8760 7488 8812 7540
rect 9496 7488 9548 7540
rect 10048 7488 10100 7540
rect 664 7395 716 7404
rect 664 7361 673 7395
rect 673 7361 707 7395
rect 707 7361 716 7395
rect 664 7352 716 7361
rect 2044 7352 2096 7404
rect 1308 7284 1360 7336
rect 1952 7148 2004 7200
rect 2596 7352 2648 7404
rect 3148 7352 3200 7404
rect 4068 7352 4120 7404
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 5908 7352 5960 7404
rect 8760 7395 8812 7404
rect 3976 7284 4028 7336
rect 4712 7284 4764 7336
rect 5724 7327 5776 7336
rect 5724 7293 5733 7327
rect 5733 7293 5767 7327
rect 5767 7293 5776 7327
rect 5724 7284 5776 7293
rect 2964 7216 3016 7268
rect 3884 7216 3936 7268
rect 6460 7284 6512 7336
rect 8760 7361 8769 7395
rect 8769 7361 8803 7395
rect 8803 7361 8812 7395
rect 8760 7352 8812 7361
rect 7932 7284 7984 7336
rect 9312 7352 9364 7404
rect 9588 7352 9640 7404
rect 10048 7352 10100 7404
rect 10416 7420 10468 7472
rect 11612 7488 11664 7540
rect 11704 7488 11756 7540
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 14188 7488 14240 7540
rect 10600 7395 10652 7404
rect 9220 7284 9272 7336
rect 9772 7284 9824 7336
rect 7564 7216 7616 7268
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 10876 7352 10928 7404
rect 11336 7395 11388 7404
rect 11336 7361 11345 7395
rect 11345 7361 11379 7395
rect 11379 7361 11388 7395
rect 11336 7352 11388 7361
rect 12072 7420 12124 7472
rect 14740 7488 14792 7540
rect 14924 7531 14976 7540
rect 14924 7497 14933 7531
rect 14933 7497 14967 7531
rect 14967 7497 14976 7531
rect 14924 7488 14976 7497
rect 16120 7488 16172 7540
rect 11796 7395 11848 7404
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 12808 7395 12860 7404
rect 11796 7352 11848 7361
rect 12808 7361 12817 7395
rect 12817 7361 12851 7395
rect 12851 7361 12860 7395
rect 12808 7352 12860 7361
rect 12716 7327 12768 7336
rect 12716 7293 12725 7327
rect 12725 7293 12759 7327
rect 12759 7293 12768 7327
rect 12716 7284 12768 7293
rect 14280 7352 14332 7404
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 15108 7420 15160 7472
rect 15384 7420 15436 7472
rect 14464 7352 14516 7361
rect 14924 7352 14976 7404
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 17316 7352 17368 7404
rect 16672 7284 16724 7336
rect 18328 7284 18380 7336
rect 3240 7148 3292 7200
rect 5264 7191 5316 7200
rect 5264 7157 5273 7191
rect 5273 7157 5307 7191
rect 5307 7157 5316 7191
rect 5264 7148 5316 7157
rect 5632 7148 5684 7200
rect 8024 7148 8076 7200
rect 8392 7191 8444 7200
rect 8392 7157 8401 7191
rect 8401 7157 8435 7191
rect 8435 7157 8444 7191
rect 8392 7148 8444 7157
rect 13728 7216 13780 7268
rect 14832 7216 14884 7268
rect 11336 7148 11388 7200
rect 12256 7148 12308 7200
rect 14096 7191 14148 7200
rect 14096 7157 14105 7191
rect 14105 7157 14139 7191
rect 14139 7157 14148 7191
rect 14096 7148 14148 7157
rect 14372 7148 14424 7200
rect 15384 7148 15436 7200
rect 17224 7191 17276 7200
rect 17224 7157 17233 7191
rect 17233 7157 17267 7191
rect 17267 7157 17276 7191
rect 17224 7148 17276 7157
rect 3478 7046 3530 7098
rect 3542 7046 3594 7098
rect 3606 7046 3658 7098
rect 3670 7046 3722 7098
rect 3734 7046 3786 7098
rect 6578 7046 6630 7098
rect 6642 7046 6694 7098
rect 6706 7046 6758 7098
rect 6770 7046 6822 7098
rect 6834 7046 6886 7098
rect 9678 7046 9730 7098
rect 9742 7046 9794 7098
rect 9806 7046 9858 7098
rect 9870 7046 9922 7098
rect 9934 7046 9986 7098
rect 12778 7046 12830 7098
rect 12842 7046 12894 7098
rect 12906 7046 12958 7098
rect 12970 7046 13022 7098
rect 13034 7046 13086 7098
rect 15878 7046 15930 7098
rect 15942 7046 15994 7098
rect 16006 7046 16058 7098
rect 16070 7046 16122 7098
rect 16134 7046 16186 7098
rect 2412 6987 2464 6996
rect 2412 6953 2421 6987
rect 2421 6953 2455 6987
rect 2455 6953 2464 6987
rect 2412 6944 2464 6953
rect 5724 6944 5776 6996
rect 6276 6944 6328 6996
rect 8760 6944 8812 6996
rect 9128 6944 9180 6996
rect 3056 6919 3108 6928
rect 3056 6885 3065 6919
rect 3065 6885 3099 6919
rect 3099 6885 3108 6919
rect 3056 6876 3108 6885
rect 940 6783 992 6792
rect 940 6749 949 6783
rect 949 6749 983 6783
rect 983 6749 992 6783
rect 940 6740 992 6749
rect 1492 6783 1544 6792
rect 1492 6749 1501 6783
rect 1501 6749 1535 6783
rect 1535 6749 1544 6783
rect 1492 6740 1544 6749
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 3240 6808 3292 6860
rect 2504 6783 2556 6792
rect 1308 6672 1360 6724
rect 1032 6604 1084 6656
rect 2504 6749 2513 6783
rect 2513 6749 2547 6783
rect 2547 6749 2556 6783
rect 2504 6740 2556 6749
rect 2964 6783 3016 6792
rect 2964 6749 2973 6783
rect 2973 6749 3007 6783
rect 3007 6749 3016 6783
rect 2964 6740 3016 6749
rect 3424 6740 3476 6792
rect 3608 6783 3660 6792
rect 3608 6749 3617 6783
rect 3617 6749 3651 6783
rect 3651 6749 3660 6783
rect 3608 6740 3660 6749
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 3976 6740 4028 6792
rect 4160 6740 4212 6792
rect 5632 6808 5684 6860
rect 5816 6808 5868 6860
rect 3884 6672 3936 6724
rect 5264 6740 5316 6792
rect 5908 6740 5960 6792
rect 7012 6851 7064 6860
rect 7012 6817 7021 6851
rect 7021 6817 7055 6851
rect 7055 6817 7064 6851
rect 7012 6808 7064 6817
rect 10416 6876 10468 6928
rect 7840 6808 7892 6860
rect 8392 6808 8444 6860
rect 8484 6808 8536 6860
rect 10692 6876 10744 6928
rect 11060 6944 11112 6996
rect 13452 6944 13504 6996
rect 12992 6876 13044 6928
rect 16396 6944 16448 6996
rect 15200 6876 15252 6928
rect 13912 6808 13964 6860
rect 14464 6808 14516 6860
rect 15016 6808 15068 6860
rect 3516 6604 3568 6656
rect 5540 6672 5592 6724
rect 7380 6715 7432 6724
rect 7380 6681 7389 6715
rect 7389 6681 7423 6715
rect 7423 6681 7432 6715
rect 7380 6672 7432 6681
rect 7564 6715 7616 6724
rect 7564 6681 7573 6715
rect 7573 6681 7607 6715
rect 7607 6681 7616 6715
rect 7564 6672 7616 6681
rect 8024 6740 8076 6792
rect 10232 6740 10284 6792
rect 10876 6740 10928 6792
rect 11060 6740 11112 6792
rect 12624 6740 12676 6792
rect 14004 6783 14056 6792
rect 14004 6749 14013 6783
rect 14013 6749 14047 6783
rect 14047 6749 14056 6783
rect 14004 6740 14056 6749
rect 16304 6808 16356 6860
rect 17224 6808 17276 6860
rect 17776 6808 17828 6860
rect 8944 6672 8996 6724
rect 10416 6715 10468 6724
rect 10416 6681 10425 6715
rect 10425 6681 10459 6715
rect 10459 6681 10468 6715
rect 10416 6672 10468 6681
rect 11336 6672 11388 6724
rect 14372 6672 14424 6724
rect 4804 6604 4856 6656
rect 5724 6604 5776 6656
rect 7472 6604 7524 6656
rect 8576 6604 8628 6656
rect 9404 6647 9456 6656
rect 9404 6613 9413 6647
rect 9413 6613 9447 6647
rect 9447 6613 9456 6647
rect 9404 6604 9456 6613
rect 9496 6647 9548 6656
rect 9496 6613 9505 6647
rect 9505 6613 9539 6647
rect 9539 6613 9548 6647
rect 9496 6604 9548 6613
rect 10784 6604 10836 6656
rect 12808 6604 12860 6656
rect 13360 6647 13412 6656
rect 13360 6613 13369 6647
rect 13369 6613 13403 6647
rect 13403 6613 13412 6647
rect 15752 6647 15804 6656
rect 13360 6604 13412 6613
rect 15752 6613 15761 6647
rect 15761 6613 15795 6647
rect 15795 6613 15804 6647
rect 15752 6604 15804 6613
rect 16212 6647 16264 6656
rect 16212 6613 16221 6647
rect 16221 6613 16255 6647
rect 16255 6613 16264 6647
rect 16212 6604 16264 6613
rect 16396 6783 16448 6792
rect 16396 6749 16405 6783
rect 16405 6749 16439 6783
rect 16439 6749 16448 6783
rect 16396 6740 16448 6749
rect 17132 6672 17184 6724
rect 16672 6604 16724 6656
rect 5028 6502 5080 6554
rect 5092 6502 5144 6554
rect 5156 6502 5208 6554
rect 5220 6502 5272 6554
rect 5284 6502 5336 6554
rect 8128 6502 8180 6554
rect 8192 6502 8244 6554
rect 8256 6502 8308 6554
rect 8320 6502 8372 6554
rect 8384 6502 8436 6554
rect 11228 6502 11280 6554
rect 11292 6502 11344 6554
rect 11356 6502 11408 6554
rect 11420 6502 11472 6554
rect 11484 6502 11536 6554
rect 14328 6502 14380 6554
rect 14392 6502 14444 6554
rect 14456 6502 14508 6554
rect 14520 6502 14572 6554
rect 14584 6502 14636 6554
rect 17428 6502 17480 6554
rect 17492 6502 17544 6554
rect 17556 6502 17608 6554
rect 17620 6502 17672 6554
rect 17684 6502 17736 6554
rect 2504 6400 2556 6452
rect 3516 6443 3568 6452
rect 3516 6409 3525 6443
rect 3525 6409 3559 6443
rect 3559 6409 3568 6443
rect 3516 6400 3568 6409
rect 5724 6443 5776 6452
rect 5724 6409 5733 6443
rect 5733 6409 5767 6443
rect 5767 6409 5776 6443
rect 5724 6400 5776 6409
rect 5908 6443 5960 6452
rect 5908 6409 5917 6443
rect 5917 6409 5951 6443
rect 5951 6409 5960 6443
rect 5908 6400 5960 6409
rect 7012 6400 7064 6452
rect 2044 6332 2096 6384
rect 1032 6307 1084 6316
rect 1032 6273 1041 6307
rect 1041 6273 1075 6307
rect 1075 6273 1084 6307
rect 1032 6264 1084 6273
rect 3056 6332 3108 6384
rect 7564 6400 7616 6452
rect 10048 6400 10100 6452
rect 10784 6400 10836 6452
rect 12808 6443 12860 6452
rect 12808 6409 12817 6443
rect 12817 6409 12851 6443
rect 12851 6409 12860 6443
rect 12808 6400 12860 6409
rect 5540 6307 5592 6316
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 5816 6307 5868 6316
rect 5816 6273 5825 6307
rect 5825 6273 5859 6307
rect 5859 6273 5868 6307
rect 5816 6264 5868 6273
rect 6000 6264 6052 6316
rect 2780 6196 2832 6248
rect 3056 6239 3108 6248
rect 3056 6205 3065 6239
rect 3065 6205 3099 6239
rect 3099 6205 3108 6239
rect 3056 6196 3108 6205
rect 6276 6196 6328 6248
rect 8484 6332 8536 6384
rect 9588 6332 9640 6384
rect 7472 6264 7524 6316
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 11152 6307 11204 6316
rect 3148 6128 3200 6180
rect 3608 6128 3660 6180
rect 2872 6103 2924 6112
rect 2872 6069 2881 6103
rect 2881 6069 2915 6103
rect 2915 6069 2924 6103
rect 2872 6060 2924 6069
rect 4068 6060 4120 6112
rect 7380 6196 7432 6248
rect 8484 6196 8536 6248
rect 7932 6128 7984 6180
rect 8024 6128 8076 6180
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 11060 6239 11112 6248
rect 11060 6205 11069 6239
rect 11069 6205 11103 6239
rect 11103 6205 11112 6239
rect 11060 6196 11112 6205
rect 9220 6128 9272 6180
rect 12164 6196 12216 6248
rect 11520 6128 11572 6180
rect 12992 6239 13044 6248
rect 12992 6205 13001 6239
rect 13001 6205 13035 6239
rect 13035 6205 13044 6239
rect 12992 6196 13044 6205
rect 13820 6400 13872 6452
rect 14004 6443 14056 6452
rect 14004 6409 14013 6443
rect 14013 6409 14047 6443
rect 14047 6409 14056 6443
rect 14004 6400 14056 6409
rect 14832 6400 14884 6452
rect 14188 6332 14240 6384
rect 14096 6307 14148 6316
rect 14096 6273 14105 6307
rect 14105 6273 14139 6307
rect 14139 6273 14148 6307
rect 14096 6264 14148 6273
rect 16212 6400 16264 6452
rect 16856 6400 16908 6452
rect 17776 6400 17828 6452
rect 18328 6443 18380 6452
rect 18328 6409 18337 6443
rect 18337 6409 18371 6443
rect 18371 6409 18380 6443
rect 18328 6400 18380 6409
rect 16304 6332 16356 6384
rect 14740 6264 14792 6316
rect 15200 6264 15252 6316
rect 14924 6196 14976 6248
rect 18512 6307 18564 6316
rect 18512 6273 18521 6307
rect 18521 6273 18555 6307
rect 18555 6273 18564 6307
rect 18512 6264 18564 6273
rect 15476 6196 15528 6248
rect 15752 6239 15804 6248
rect 15752 6205 15761 6239
rect 15761 6205 15795 6239
rect 15795 6205 15804 6239
rect 15752 6196 15804 6205
rect 17868 6239 17920 6248
rect 17868 6205 17877 6239
rect 17877 6205 17911 6239
rect 17911 6205 17920 6239
rect 17868 6196 17920 6205
rect 14464 6128 14516 6180
rect 17316 6128 17368 6180
rect 11060 6060 11112 6112
rect 15752 6060 15804 6112
rect 3478 5958 3530 6010
rect 3542 5958 3594 6010
rect 3606 5958 3658 6010
rect 3670 5958 3722 6010
rect 3734 5958 3786 6010
rect 6578 5958 6630 6010
rect 6642 5958 6694 6010
rect 6706 5958 6758 6010
rect 6770 5958 6822 6010
rect 6834 5958 6886 6010
rect 9678 5958 9730 6010
rect 9742 5958 9794 6010
rect 9806 5958 9858 6010
rect 9870 5958 9922 6010
rect 9934 5958 9986 6010
rect 12778 5958 12830 6010
rect 12842 5958 12894 6010
rect 12906 5958 12958 6010
rect 12970 5958 13022 6010
rect 13034 5958 13086 6010
rect 15878 5958 15930 6010
rect 15942 5958 15994 6010
rect 16006 5958 16058 6010
rect 16070 5958 16122 6010
rect 16134 5958 16186 6010
rect 2872 5856 2924 5908
rect 3056 5856 3108 5908
rect 3884 5856 3936 5908
rect 5632 5856 5684 5908
rect 7196 5856 7248 5908
rect 7748 5856 7800 5908
rect 5816 5788 5868 5840
rect 7380 5788 7432 5840
rect 940 5720 992 5772
rect 6460 5720 6512 5772
rect 2780 5584 2832 5636
rect 4804 5584 4856 5636
rect 9680 5720 9732 5772
rect 8576 5652 8628 5704
rect 15660 5856 15712 5908
rect 12624 5788 12676 5840
rect 15476 5831 15528 5840
rect 15476 5797 15485 5831
rect 15485 5797 15519 5831
rect 15519 5797 15528 5831
rect 15476 5788 15528 5797
rect 17868 5856 17920 5908
rect 16396 5788 16448 5840
rect 13452 5720 13504 5772
rect 14832 5720 14884 5772
rect 14464 5695 14516 5704
rect 4068 5516 4120 5568
rect 5540 5516 5592 5568
rect 7012 5516 7064 5568
rect 7932 5584 7984 5636
rect 11520 5627 11572 5636
rect 11520 5593 11529 5627
rect 11529 5593 11563 5627
rect 11563 5593 11572 5627
rect 11520 5584 11572 5593
rect 12256 5584 12308 5636
rect 10416 5516 10468 5568
rect 13176 5516 13228 5568
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 14740 5584 14792 5636
rect 16212 5584 16264 5636
rect 16764 5627 16816 5636
rect 16764 5593 16773 5627
rect 16773 5593 16807 5627
rect 16807 5593 16816 5627
rect 16764 5584 16816 5593
rect 16856 5584 16908 5636
rect 17224 5584 17276 5636
rect 14832 5516 14884 5568
rect 15752 5559 15804 5568
rect 15752 5525 15761 5559
rect 15761 5525 15795 5559
rect 15795 5525 15804 5559
rect 15752 5516 15804 5525
rect 15844 5516 15896 5568
rect 16580 5516 16632 5568
rect 16672 5516 16724 5568
rect 5028 5414 5080 5466
rect 5092 5414 5144 5466
rect 5156 5414 5208 5466
rect 5220 5414 5272 5466
rect 5284 5414 5336 5466
rect 8128 5414 8180 5466
rect 8192 5414 8244 5466
rect 8256 5414 8308 5466
rect 8320 5414 8372 5466
rect 8384 5414 8436 5466
rect 11228 5414 11280 5466
rect 11292 5414 11344 5466
rect 11356 5414 11408 5466
rect 11420 5414 11472 5466
rect 11484 5414 11536 5466
rect 14328 5414 14380 5466
rect 14392 5414 14444 5466
rect 14456 5414 14508 5466
rect 14520 5414 14572 5466
rect 14584 5414 14636 5466
rect 17428 5414 17480 5466
rect 17492 5414 17544 5466
rect 17556 5414 17608 5466
rect 17620 5414 17672 5466
rect 17684 5414 17736 5466
rect 4068 5355 4120 5364
rect 4068 5321 4077 5355
rect 4077 5321 4111 5355
rect 4111 5321 4120 5355
rect 4068 5312 4120 5321
rect 5540 5355 5592 5364
rect 5540 5321 5549 5355
rect 5549 5321 5583 5355
rect 5583 5321 5592 5355
rect 5540 5312 5592 5321
rect 7840 5312 7892 5364
rect 9404 5355 9456 5364
rect 9404 5321 9413 5355
rect 9413 5321 9447 5355
rect 9447 5321 9456 5355
rect 9404 5312 9456 5321
rect 10692 5312 10744 5364
rect 7012 5244 7064 5296
rect 7196 5244 7248 5296
rect 7932 5244 7984 5296
rect 9680 5287 9732 5296
rect 5632 5219 5684 5228
rect 5632 5185 5641 5219
rect 5641 5185 5675 5219
rect 5675 5185 5684 5219
rect 5632 5176 5684 5185
rect 8484 5176 8536 5228
rect 9680 5253 9689 5287
rect 9689 5253 9723 5287
rect 9723 5253 9732 5287
rect 9680 5244 9732 5253
rect 10140 5244 10192 5296
rect 5908 5108 5960 5160
rect 10416 5176 10468 5228
rect 12256 5244 12308 5296
rect 13360 5312 13412 5364
rect 12624 5176 12676 5228
rect 13452 5244 13504 5296
rect 14740 5312 14792 5364
rect 16304 5355 16356 5364
rect 16304 5321 16313 5355
rect 16313 5321 16347 5355
rect 16347 5321 16356 5355
rect 16304 5312 16356 5321
rect 16580 5312 16632 5364
rect 16212 5219 16264 5228
rect 16212 5185 16221 5219
rect 16221 5185 16255 5219
rect 16255 5185 16264 5219
rect 16212 5176 16264 5185
rect 16672 5219 16724 5228
rect 16672 5185 16681 5219
rect 16681 5185 16715 5219
rect 16715 5185 16724 5219
rect 16672 5176 16724 5185
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 8944 5151 8996 5160
rect 8944 5117 8953 5151
rect 8953 5117 8987 5151
rect 8987 5117 8996 5151
rect 8944 5108 8996 5117
rect 10324 5108 10376 5160
rect 13176 5151 13228 5160
rect 6920 4972 6972 5024
rect 13176 5117 13185 5151
rect 13185 5117 13219 5151
rect 13219 5117 13228 5151
rect 13176 5108 13228 5117
rect 15844 5151 15896 5160
rect 15844 5117 15853 5151
rect 15853 5117 15887 5151
rect 15887 5117 15896 5151
rect 15844 5108 15896 5117
rect 16764 5108 16816 5160
rect 18144 4972 18196 5024
rect 18328 5015 18380 5024
rect 18328 4981 18337 5015
rect 18337 4981 18371 5015
rect 18371 4981 18380 5015
rect 18328 4972 18380 4981
rect 3478 4870 3530 4922
rect 3542 4870 3594 4922
rect 3606 4870 3658 4922
rect 3670 4870 3722 4922
rect 3734 4870 3786 4922
rect 6578 4870 6630 4922
rect 6642 4870 6694 4922
rect 6706 4870 6758 4922
rect 6770 4870 6822 4922
rect 6834 4870 6886 4922
rect 9678 4870 9730 4922
rect 9742 4870 9794 4922
rect 9806 4870 9858 4922
rect 9870 4870 9922 4922
rect 9934 4870 9986 4922
rect 12778 4870 12830 4922
rect 12842 4870 12894 4922
rect 12906 4870 12958 4922
rect 12970 4870 13022 4922
rect 13034 4870 13086 4922
rect 15878 4870 15930 4922
rect 15942 4870 15994 4922
rect 16006 4870 16058 4922
rect 16070 4870 16122 4922
rect 16134 4870 16186 4922
rect 940 4675 992 4684
rect 940 4641 949 4675
rect 949 4641 983 4675
rect 983 4641 992 4675
rect 940 4632 992 4641
rect 5908 4811 5960 4820
rect 5908 4777 5917 4811
rect 5917 4777 5951 4811
rect 5951 4777 5960 4811
rect 5908 4768 5960 4777
rect 7932 4811 7984 4820
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 9404 4768 9456 4820
rect 4068 4700 4120 4752
rect 2136 4675 2188 4684
rect 2136 4641 2145 4675
rect 2145 4641 2179 4675
rect 2179 4641 2188 4675
rect 5632 4700 5684 4752
rect 2136 4632 2188 4641
rect 1308 4607 1360 4616
rect 1308 4573 1317 4607
rect 1317 4573 1351 4607
rect 1351 4573 1360 4607
rect 1308 4564 1360 4573
rect 4068 4564 4120 4616
rect 3884 4496 3936 4548
rect 2780 4428 2832 4480
rect 3976 4428 4028 4480
rect 4436 4471 4488 4480
rect 4436 4437 4445 4471
rect 4445 4437 4479 4471
rect 4479 4437 4488 4471
rect 4436 4428 4488 4437
rect 4804 4428 4856 4480
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 6920 4675 6972 4684
rect 6920 4641 6929 4675
rect 6929 4641 6963 4675
rect 6963 4641 6972 4675
rect 6920 4632 6972 4641
rect 7932 4632 7984 4684
rect 18328 4768 18380 4820
rect 10416 4632 10468 4684
rect 12256 4632 12308 4684
rect 12624 4632 12676 4684
rect 14096 4675 14148 4684
rect 14096 4641 14105 4675
rect 14105 4641 14139 4675
rect 14139 4641 14148 4675
rect 14096 4632 14148 4641
rect 13268 4564 13320 4616
rect 13360 4564 13412 4616
rect 17960 4564 18012 4616
rect 18236 4607 18288 4616
rect 18236 4573 18245 4607
rect 18245 4573 18279 4607
rect 18279 4573 18288 4607
rect 18236 4564 18288 4573
rect 7104 4496 7156 4548
rect 12256 4496 12308 4548
rect 13452 4496 13504 4548
rect 14188 4496 14240 4548
rect 15752 4496 15804 4548
rect 16856 4496 16908 4548
rect 6920 4428 6972 4480
rect 12716 4428 12768 4480
rect 15476 4471 15528 4480
rect 15476 4437 15485 4471
rect 15485 4437 15519 4471
rect 15519 4437 15528 4471
rect 15476 4428 15528 4437
rect 16212 4471 16264 4480
rect 16212 4437 16221 4471
rect 16221 4437 16255 4471
rect 16255 4437 16264 4471
rect 16212 4428 16264 4437
rect 17868 4428 17920 4480
rect 5028 4326 5080 4378
rect 5092 4326 5144 4378
rect 5156 4326 5208 4378
rect 5220 4326 5272 4378
rect 5284 4326 5336 4378
rect 8128 4326 8180 4378
rect 8192 4326 8244 4378
rect 8256 4326 8308 4378
rect 8320 4326 8372 4378
rect 8384 4326 8436 4378
rect 11228 4326 11280 4378
rect 11292 4326 11344 4378
rect 11356 4326 11408 4378
rect 11420 4326 11472 4378
rect 11484 4326 11536 4378
rect 14328 4326 14380 4378
rect 14392 4326 14444 4378
rect 14456 4326 14508 4378
rect 14520 4326 14572 4378
rect 14584 4326 14636 4378
rect 17428 4326 17480 4378
rect 17492 4326 17544 4378
rect 17556 4326 17608 4378
rect 17620 4326 17672 4378
rect 17684 4326 17736 4378
rect 2780 4224 2832 4276
rect 4436 4224 4488 4276
rect 7104 4267 7156 4276
rect 7104 4233 7113 4267
rect 7113 4233 7147 4267
rect 7147 4233 7156 4267
rect 7104 4224 7156 4233
rect 10692 4267 10744 4276
rect 940 4199 992 4208
rect 940 4165 949 4199
rect 949 4165 983 4199
rect 983 4165 992 4199
rect 940 4156 992 4165
rect 2780 4088 2832 4140
rect 3976 4156 4028 4208
rect 9404 4156 9456 4208
rect 10692 4233 10701 4267
rect 10701 4233 10735 4267
rect 10735 4233 10744 4267
rect 10692 4224 10744 4233
rect 14188 4224 14240 4276
rect 17960 4224 18012 4276
rect 4068 4131 4120 4140
rect 1308 4020 1360 4072
rect 4068 4097 4077 4131
rect 4077 4097 4111 4131
rect 4111 4097 4120 4131
rect 4068 4088 4120 4097
rect 4896 4088 4948 4140
rect 6092 4088 6144 4140
rect 6920 4088 6972 4140
rect 7748 4131 7800 4140
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 4804 4063 4856 4072
rect 4804 4029 4813 4063
rect 4813 4029 4847 4063
rect 4847 4029 4856 4063
rect 4804 4020 4856 4029
rect 6460 4063 6512 4072
rect 6460 4029 6469 4063
rect 6469 4029 6503 4063
rect 6503 4029 6512 4063
rect 6460 4020 6512 4029
rect 8208 4020 8260 4072
rect 10048 4088 10100 4140
rect 12256 4156 12308 4208
rect 11244 4131 11296 4140
rect 11244 4097 11253 4131
rect 11253 4097 11287 4131
rect 11287 4097 11296 4131
rect 11244 4088 11296 4097
rect 15476 4131 15528 4140
rect 10692 4020 10744 4072
rect 12716 4063 12768 4072
rect 12716 4029 12725 4063
rect 12725 4029 12759 4063
rect 12759 4029 12768 4063
rect 12716 4020 12768 4029
rect 13360 4020 13412 4072
rect 2780 3884 2832 3936
rect 6368 3884 6420 3936
rect 8024 3884 8076 3936
rect 10048 3884 10100 3936
rect 10232 3927 10284 3936
rect 10232 3893 10241 3927
rect 10241 3893 10275 3927
rect 10275 3893 10284 3927
rect 10232 3884 10284 3893
rect 12256 3927 12308 3936
rect 12256 3893 12265 3927
rect 12265 3893 12299 3927
rect 12299 3893 12308 3927
rect 12256 3884 12308 3893
rect 12440 3884 12492 3936
rect 13268 3884 13320 3936
rect 15476 4097 15485 4131
rect 15485 4097 15519 4131
rect 15519 4097 15528 4131
rect 15476 4088 15528 4097
rect 16396 4088 16448 4140
rect 18512 4131 18564 4140
rect 18512 4097 18521 4131
rect 18521 4097 18555 4131
rect 18555 4097 18564 4131
rect 18512 4088 18564 4097
rect 15384 3952 15436 4004
rect 15200 3927 15252 3936
rect 15200 3893 15209 3927
rect 15209 3893 15243 3927
rect 15243 3893 15252 3927
rect 15200 3884 15252 3893
rect 15476 3884 15528 3936
rect 3478 3782 3530 3834
rect 3542 3782 3594 3834
rect 3606 3782 3658 3834
rect 3670 3782 3722 3834
rect 3734 3782 3786 3834
rect 6578 3782 6630 3834
rect 6642 3782 6694 3834
rect 6706 3782 6758 3834
rect 6770 3782 6822 3834
rect 6834 3782 6886 3834
rect 9678 3782 9730 3834
rect 9742 3782 9794 3834
rect 9806 3782 9858 3834
rect 9870 3782 9922 3834
rect 9934 3782 9986 3834
rect 12778 3782 12830 3834
rect 12842 3782 12894 3834
rect 12906 3782 12958 3834
rect 12970 3782 13022 3834
rect 13034 3782 13086 3834
rect 15878 3782 15930 3834
rect 15942 3782 15994 3834
rect 16006 3782 16058 3834
rect 16070 3782 16122 3834
rect 16134 3782 16186 3834
rect 3884 3680 3936 3732
rect 6460 3680 6512 3732
rect 7564 3680 7616 3732
rect 7932 3680 7984 3732
rect 8208 3723 8260 3732
rect 8208 3689 8217 3723
rect 8217 3689 8251 3723
rect 8251 3689 8260 3723
rect 8208 3680 8260 3689
rect 13268 3680 13320 3732
rect 16304 3680 16356 3732
rect 10232 3655 10284 3664
rect 2136 3587 2188 3596
rect 2136 3553 2145 3587
rect 2145 3553 2179 3587
rect 2179 3553 2188 3587
rect 2136 3544 2188 3553
rect 4436 3544 4488 3596
rect 4068 3519 4120 3528
rect 4068 3485 4077 3519
rect 4077 3485 4111 3519
rect 4111 3485 4120 3519
rect 4068 3476 4120 3485
rect 2412 3451 2464 3460
rect 2412 3417 2421 3451
rect 2421 3417 2455 3451
rect 2455 3417 2464 3451
rect 2412 3408 2464 3417
rect 2780 3340 2832 3392
rect 3884 3408 3936 3460
rect 4712 3408 4764 3460
rect 6368 3476 6420 3528
rect 6920 3476 6972 3528
rect 7555 3519 7607 3528
rect 7555 3485 7571 3519
rect 7571 3485 7607 3519
rect 7555 3476 7607 3485
rect 10232 3621 10241 3655
rect 10241 3621 10275 3655
rect 10275 3621 10284 3655
rect 10232 3612 10284 3621
rect 10048 3544 10100 3596
rect 10692 3544 10744 3596
rect 8852 3519 8904 3528
rect 8852 3485 8861 3519
rect 8861 3485 8895 3519
rect 8895 3485 8904 3519
rect 8852 3476 8904 3485
rect 7932 3408 7984 3460
rect 10508 3476 10560 3528
rect 11244 3476 11296 3528
rect 12072 3476 12124 3528
rect 4344 3340 4396 3392
rect 5816 3340 5868 3392
rect 10600 3408 10652 3460
rect 13452 3519 13504 3528
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 14096 3544 14148 3596
rect 16304 3544 16356 3596
rect 18236 3587 18288 3596
rect 18236 3553 18245 3587
rect 18245 3553 18279 3587
rect 18279 3553 18288 3587
rect 18236 3544 18288 3553
rect 13728 3476 13780 3528
rect 15200 3476 15252 3528
rect 16488 3476 16540 3528
rect 17868 3519 17920 3528
rect 17868 3485 17877 3519
rect 17877 3485 17911 3519
rect 17911 3485 17920 3519
rect 17868 3476 17920 3485
rect 15292 3408 15344 3460
rect 16212 3408 16264 3460
rect 10416 3383 10468 3392
rect 10416 3349 10425 3383
rect 10425 3349 10459 3383
rect 10459 3349 10468 3383
rect 10416 3340 10468 3349
rect 15200 3340 15252 3392
rect 15660 3340 15712 3392
rect 15752 3383 15804 3392
rect 15752 3349 15761 3383
rect 15761 3349 15795 3383
rect 15795 3349 15804 3383
rect 16120 3383 16172 3392
rect 15752 3340 15804 3349
rect 16120 3349 16129 3383
rect 16129 3349 16163 3383
rect 16163 3349 16172 3383
rect 16120 3340 16172 3349
rect 16396 3340 16448 3392
rect 5028 3238 5080 3290
rect 5092 3238 5144 3290
rect 5156 3238 5208 3290
rect 5220 3238 5272 3290
rect 5284 3238 5336 3290
rect 8128 3238 8180 3290
rect 8192 3238 8244 3290
rect 8256 3238 8308 3290
rect 8320 3238 8372 3290
rect 8384 3238 8436 3290
rect 11228 3238 11280 3290
rect 11292 3238 11344 3290
rect 11356 3238 11408 3290
rect 11420 3238 11472 3290
rect 11484 3238 11536 3290
rect 14328 3238 14380 3290
rect 14392 3238 14444 3290
rect 14456 3238 14508 3290
rect 14520 3238 14572 3290
rect 14584 3238 14636 3290
rect 17428 3238 17480 3290
rect 17492 3238 17544 3290
rect 17556 3238 17608 3290
rect 17620 3238 17672 3290
rect 17684 3238 17736 3290
rect 2412 3136 2464 3188
rect 7196 3136 7248 3188
rect 2780 3068 2832 3120
rect 3056 3000 3108 3052
rect 3332 3000 3384 3052
rect 4068 3068 4120 3120
rect 4344 3111 4396 3120
rect 4344 3077 4353 3111
rect 4353 3077 4387 3111
rect 4387 3077 4396 3111
rect 4344 3068 4396 3077
rect 5724 3068 5776 3120
rect 3976 3043 4028 3052
rect 3976 3009 3985 3043
rect 3985 3009 4019 3043
rect 4019 3009 4028 3043
rect 3976 3000 4028 3009
rect 4436 3043 4488 3052
rect 4436 3009 4445 3043
rect 4445 3009 4479 3043
rect 4479 3009 4488 3043
rect 4436 3000 4488 3009
rect 4712 3043 4764 3052
rect 4712 3009 4721 3043
rect 4721 3009 4755 3043
rect 4755 3009 4764 3043
rect 4712 3000 4764 3009
rect 5816 3043 5868 3052
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 5816 3000 5868 3009
rect 7380 3068 7432 3120
rect 6092 3000 6144 3052
rect 7196 3000 7248 3052
rect 10232 3136 10284 3188
rect 10508 3136 10560 3188
rect 9220 3068 9272 3120
rect 13176 3136 13228 3188
rect 13728 3136 13780 3188
rect 15292 3136 15344 3188
rect 16488 3179 16540 3188
rect 16488 3145 16497 3179
rect 16497 3145 16531 3179
rect 16531 3145 16540 3179
rect 16488 3136 16540 3145
rect 7932 3000 7984 3052
rect 10048 3000 10100 3052
rect 10232 3000 10284 3052
rect 10416 3043 10468 3052
rect 10416 3009 10425 3043
rect 10425 3009 10459 3043
rect 10459 3009 10468 3043
rect 10416 3000 10468 3009
rect 10784 3043 10836 3052
rect 10784 3009 10793 3043
rect 10793 3009 10827 3043
rect 10827 3009 10836 3043
rect 10784 3000 10836 3009
rect 11152 3043 11204 3052
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 11796 3000 11848 3052
rect 13452 3000 13504 3052
rect 14004 3000 14056 3052
rect 15200 3043 15252 3052
rect 15200 3009 15209 3043
rect 15209 3009 15243 3043
rect 15243 3009 15252 3043
rect 15200 3000 15252 3009
rect 15476 3111 15528 3120
rect 15476 3077 15485 3111
rect 15485 3077 15519 3111
rect 15519 3077 15528 3111
rect 15660 3111 15712 3120
rect 15476 3068 15528 3077
rect 15660 3077 15669 3111
rect 15669 3077 15703 3111
rect 15703 3077 15712 3111
rect 15660 3068 15712 3077
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 7472 2975 7524 2984
rect 3516 2864 3568 2916
rect 3700 2864 3752 2916
rect 7472 2941 7481 2975
rect 7481 2941 7515 2975
rect 7515 2941 7524 2975
rect 7472 2932 7524 2941
rect 2504 2796 2556 2848
rect 2780 2796 2832 2848
rect 5816 2839 5868 2848
rect 5816 2805 5825 2839
rect 5825 2805 5859 2839
rect 5859 2805 5868 2839
rect 5816 2796 5868 2805
rect 7104 2864 7156 2916
rect 7288 2864 7340 2916
rect 8576 2932 8628 2984
rect 12440 2932 12492 2984
rect 11060 2864 11112 2916
rect 7656 2796 7708 2848
rect 12624 2796 12676 2848
rect 16120 2932 16172 2984
rect 14188 2796 14240 2848
rect 3478 2694 3530 2746
rect 3542 2694 3594 2746
rect 3606 2694 3658 2746
rect 3670 2694 3722 2746
rect 3734 2694 3786 2746
rect 6578 2694 6630 2746
rect 6642 2694 6694 2746
rect 6706 2694 6758 2746
rect 6770 2694 6822 2746
rect 6834 2694 6886 2746
rect 9678 2694 9730 2746
rect 9742 2694 9794 2746
rect 9806 2694 9858 2746
rect 9870 2694 9922 2746
rect 9934 2694 9986 2746
rect 12778 2694 12830 2746
rect 12842 2694 12894 2746
rect 12906 2694 12958 2746
rect 12970 2694 13022 2746
rect 13034 2694 13086 2746
rect 15878 2694 15930 2746
rect 15942 2694 15994 2746
rect 16006 2694 16058 2746
rect 16070 2694 16122 2746
rect 16134 2694 16186 2746
rect 3976 2592 4028 2644
rect 3148 2524 3200 2576
rect 664 2456 716 2508
rect 2688 2456 2740 2508
rect 3332 2499 3384 2508
rect 3332 2465 3341 2499
rect 3341 2465 3375 2499
rect 3375 2465 3384 2499
rect 3332 2456 3384 2465
rect 2964 2388 3016 2440
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 3884 2431 3936 2440
rect 3884 2397 3893 2431
rect 3893 2397 3927 2431
rect 3927 2397 3936 2431
rect 5908 2524 5960 2576
rect 6920 2567 6972 2576
rect 6920 2533 6929 2567
rect 6929 2533 6963 2567
rect 6963 2533 6972 2567
rect 6920 2524 6972 2533
rect 7288 2567 7340 2576
rect 7288 2533 7297 2567
rect 7297 2533 7331 2567
rect 7331 2533 7340 2567
rect 7288 2524 7340 2533
rect 3884 2388 3936 2397
rect 3056 2320 3108 2372
rect 3608 2320 3660 2372
rect 5448 2388 5500 2440
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 6000 2431 6052 2440
rect 6000 2397 6009 2431
rect 6009 2397 6043 2431
rect 6043 2397 6052 2431
rect 6000 2388 6052 2397
rect 6460 2431 6512 2440
rect 6460 2397 6469 2431
rect 6469 2397 6503 2431
rect 6503 2397 6512 2431
rect 6460 2388 6512 2397
rect 7012 2431 7064 2440
rect 1676 2295 1728 2304
rect 1676 2261 1685 2295
rect 1685 2261 1719 2295
rect 1719 2261 1728 2295
rect 1676 2252 1728 2261
rect 2044 2252 2096 2304
rect 2780 2252 2832 2304
rect 3976 2252 4028 2304
rect 4896 2252 4948 2304
rect 5724 2320 5776 2372
rect 7012 2397 7021 2431
rect 7021 2397 7055 2431
rect 7055 2397 7064 2431
rect 7012 2388 7064 2397
rect 8852 2456 8904 2508
rect 7288 2431 7340 2440
rect 7288 2397 7297 2431
rect 7297 2397 7331 2431
rect 7331 2397 7340 2431
rect 7288 2388 7340 2397
rect 7472 2388 7524 2440
rect 5540 2252 5592 2304
rect 5908 2252 5960 2304
rect 7932 2388 7984 2440
rect 11796 2592 11848 2644
rect 10784 2524 10836 2576
rect 11704 2524 11756 2576
rect 12256 2592 12308 2644
rect 13452 2592 13504 2644
rect 14556 2592 14608 2644
rect 15108 2592 15160 2644
rect 15752 2592 15804 2644
rect 13084 2524 13136 2576
rect 10048 2456 10100 2508
rect 11060 2499 11112 2508
rect 11060 2465 11069 2499
rect 11069 2465 11103 2499
rect 11103 2465 11112 2499
rect 11060 2456 11112 2465
rect 7104 2252 7156 2304
rect 12992 2388 13044 2440
rect 13360 2388 13412 2440
rect 14188 2456 14240 2508
rect 15292 2456 15344 2508
rect 18236 2499 18288 2508
rect 18236 2465 18245 2499
rect 18245 2465 18279 2499
rect 18279 2465 18288 2499
rect 18236 2456 18288 2465
rect 10232 2320 10284 2372
rect 11704 2320 11756 2372
rect 10324 2252 10376 2304
rect 12440 2252 12492 2304
rect 13544 2320 13596 2372
rect 14096 2320 14148 2372
rect 14556 2320 14608 2372
rect 15844 2363 15896 2372
rect 15844 2329 15853 2363
rect 15853 2329 15887 2363
rect 15887 2329 15896 2363
rect 15844 2320 15896 2329
rect 17960 2363 18012 2372
rect 17960 2329 17969 2363
rect 17969 2329 18003 2363
rect 18003 2329 18012 2363
rect 17960 2320 18012 2329
rect 14740 2252 14792 2304
rect 5028 2150 5080 2202
rect 5092 2150 5144 2202
rect 5156 2150 5208 2202
rect 5220 2150 5272 2202
rect 5284 2150 5336 2202
rect 8128 2150 8180 2202
rect 8192 2150 8244 2202
rect 8256 2150 8308 2202
rect 8320 2150 8372 2202
rect 8384 2150 8436 2202
rect 11228 2150 11280 2202
rect 11292 2150 11344 2202
rect 11356 2150 11408 2202
rect 11420 2150 11472 2202
rect 11484 2150 11536 2202
rect 14328 2150 14380 2202
rect 14392 2150 14444 2202
rect 14456 2150 14508 2202
rect 14520 2150 14572 2202
rect 14584 2150 14636 2202
rect 17428 2150 17480 2202
rect 17492 2150 17544 2202
rect 17556 2150 17608 2202
rect 17620 2150 17672 2202
rect 17684 2150 17736 2202
rect 664 2091 716 2100
rect 664 2057 673 2091
rect 673 2057 707 2091
rect 707 2057 716 2091
rect 664 2048 716 2057
rect 2964 2091 3016 2100
rect 2044 1980 2096 2032
rect 2136 1980 2188 2032
rect 2964 2057 2973 2091
rect 2973 2057 3007 2091
rect 3007 2057 3016 2091
rect 2964 2048 3016 2057
rect 3240 1980 3292 2032
rect 2504 1955 2556 1964
rect 2504 1921 2513 1955
rect 2513 1921 2547 1955
rect 2547 1921 2556 1955
rect 2504 1912 2556 1921
rect 2688 1955 2740 1964
rect 2688 1921 2697 1955
rect 2697 1921 2731 1955
rect 2731 1921 2740 1955
rect 2688 1912 2740 1921
rect 3148 1912 3200 1964
rect 3608 2048 3660 2100
rect 7288 2048 7340 2100
rect 1676 1844 1728 1896
rect 3608 1955 3660 1964
rect 3608 1921 3617 1955
rect 3617 1921 3651 1955
rect 3651 1921 3660 1955
rect 3608 1912 3660 1921
rect 3884 1912 3936 1964
rect 5632 1980 5684 2032
rect 6920 1980 6972 2032
rect 8484 2048 8536 2100
rect 10324 2048 10376 2100
rect 13360 2048 13412 2100
rect 13544 2091 13596 2100
rect 13544 2057 13553 2091
rect 13553 2057 13587 2091
rect 13587 2057 13596 2091
rect 13544 2048 13596 2057
rect 13636 2048 13688 2100
rect 4896 1912 4948 1964
rect 5540 1955 5592 1964
rect 5540 1921 5549 1955
rect 5549 1921 5583 1955
rect 5583 1921 5592 1955
rect 5540 1912 5592 1921
rect 3056 1776 3108 1828
rect 6000 1912 6052 1964
rect 7656 1955 7708 1964
rect 6368 1844 6420 1896
rect 7656 1921 7665 1955
rect 7665 1921 7699 1955
rect 7699 1921 7708 1955
rect 7656 1912 7708 1921
rect 8116 1912 8168 1964
rect 8852 1980 8904 2032
rect 3516 1776 3568 1828
rect 10508 1912 10560 1964
rect 10232 1887 10284 1896
rect 10232 1853 10241 1887
rect 10241 1853 10275 1887
rect 10275 1853 10284 1887
rect 10232 1844 10284 1853
rect 3976 1708 4028 1760
rect 4712 1708 4764 1760
rect 5356 1751 5408 1760
rect 5356 1717 5365 1751
rect 5365 1717 5399 1751
rect 5399 1717 5408 1751
rect 5356 1708 5408 1717
rect 7012 1708 7064 1760
rect 9220 1708 9272 1760
rect 9496 1708 9548 1760
rect 9588 1708 9640 1760
rect 11060 1912 11112 1964
rect 11244 1912 11296 1964
rect 12624 1912 12676 1964
rect 10968 1887 11020 1896
rect 10968 1853 10977 1887
rect 10977 1853 11011 1887
rect 11011 1853 11020 1887
rect 10968 1844 11020 1853
rect 13084 1955 13136 1964
rect 13084 1921 13093 1955
rect 13093 1921 13127 1955
rect 13127 1921 13136 1955
rect 13084 1912 13136 1921
rect 14188 1912 14240 1964
rect 15568 2048 15620 2100
rect 14740 1980 14792 2032
rect 15292 1980 15344 2032
rect 18144 2091 18196 2100
rect 18144 2057 18153 2091
rect 18153 2057 18187 2091
rect 18187 2057 18196 2091
rect 18144 2048 18196 2057
rect 18236 1980 18288 2032
rect 17224 1912 17276 1964
rect 18052 1955 18104 1964
rect 18052 1921 18061 1955
rect 18061 1921 18095 1955
rect 18095 1921 18104 1955
rect 18052 1912 18104 1921
rect 18512 1955 18564 1964
rect 18512 1921 18521 1955
rect 18521 1921 18555 1955
rect 18555 1921 18564 1955
rect 18512 1912 18564 1921
rect 13728 1844 13780 1896
rect 15844 1887 15896 1896
rect 11152 1708 11204 1760
rect 11704 1708 11756 1760
rect 12256 1751 12308 1760
rect 12256 1717 12265 1751
rect 12265 1717 12299 1751
rect 12299 1717 12308 1751
rect 15844 1853 15853 1887
rect 15853 1853 15887 1887
rect 15887 1853 15896 1887
rect 16580 1887 16632 1896
rect 15844 1844 15896 1853
rect 14924 1776 14976 1828
rect 16580 1853 16589 1887
rect 16589 1853 16623 1887
rect 16623 1853 16632 1887
rect 16580 1844 16632 1853
rect 17868 1887 17920 1896
rect 17868 1853 17877 1887
rect 17877 1853 17911 1887
rect 17911 1853 17920 1887
rect 17868 1844 17920 1853
rect 12256 1708 12308 1717
rect 14740 1708 14792 1760
rect 15292 1751 15344 1760
rect 15292 1717 15301 1751
rect 15301 1717 15335 1751
rect 15335 1717 15344 1751
rect 15292 1708 15344 1717
rect 18328 1751 18380 1760
rect 18328 1717 18337 1751
rect 18337 1717 18371 1751
rect 18371 1717 18380 1751
rect 18328 1708 18380 1717
rect 3478 1606 3530 1658
rect 3542 1606 3594 1658
rect 3606 1606 3658 1658
rect 3670 1606 3722 1658
rect 3734 1606 3786 1658
rect 6578 1606 6630 1658
rect 6642 1606 6694 1658
rect 6706 1606 6758 1658
rect 6770 1606 6822 1658
rect 6834 1606 6886 1658
rect 9678 1606 9730 1658
rect 9742 1606 9794 1658
rect 9806 1606 9858 1658
rect 9870 1606 9922 1658
rect 9934 1606 9986 1658
rect 12778 1606 12830 1658
rect 12842 1606 12894 1658
rect 12906 1606 12958 1658
rect 12970 1606 13022 1658
rect 13034 1606 13086 1658
rect 15878 1606 15930 1658
rect 15942 1606 15994 1658
rect 16006 1606 16058 1658
rect 16070 1606 16122 1658
rect 16134 1606 16186 1658
rect 5448 1504 5500 1556
rect 7932 1504 7984 1556
rect 2136 1411 2188 1420
rect 2136 1377 2145 1411
rect 2145 1377 2179 1411
rect 2179 1377 2188 1411
rect 2136 1368 2188 1377
rect 5356 1368 5408 1420
rect 5724 1368 5776 1420
rect 8300 1436 8352 1488
rect 9220 1504 9272 1556
rect 7932 1368 7984 1420
rect 9312 1436 9364 1488
rect 9588 1436 9640 1488
rect 8668 1368 8720 1420
rect 10324 1436 10376 1488
rect 3976 1300 4028 1352
rect 4620 1343 4672 1352
rect 4620 1309 4629 1343
rect 4629 1309 4663 1343
rect 4663 1309 4672 1343
rect 4620 1300 4672 1309
rect 4804 1300 4856 1352
rect 6368 1300 6420 1352
rect 3976 1164 4028 1216
rect 7288 1300 7340 1352
rect 4804 1164 4856 1216
rect 6092 1164 6144 1216
rect 6920 1164 6972 1216
rect 7196 1164 7248 1216
rect 8208 1300 8260 1352
rect 10600 1343 10652 1352
rect 10600 1309 10609 1343
rect 10609 1309 10643 1343
rect 10643 1309 10652 1343
rect 10600 1300 10652 1309
rect 11244 1343 11296 1352
rect 8484 1232 8536 1284
rect 11244 1309 11253 1343
rect 11253 1309 11287 1343
rect 11287 1309 11296 1343
rect 11244 1300 11296 1309
rect 12440 1504 12492 1556
rect 13728 1504 13780 1556
rect 17868 1504 17920 1556
rect 17960 1504 18012 1556
rect 18512 1547 18564 1556
rect 18512 1513 18521 1547
rect 18521 1513 18555 1547
rect 18555 1513 18564 1547
rect 18512 1504 18564 1513
rect 12256 1411 12308 1420
rect 12256 1377 12265 1411
rect 12265 1377 12299 1411
rect 12299 1377 12308 1411
rect 12256 1368 12308 1377
rect 13084 1411 13136 1420
rect 13084 1377 13093 1411
rect 13093 1377 13127 1411
rect 13127 1377 13136 1411
rect 13084 1368 13136 1377
rect 13728 1368 13780 1420
rect 14004 1411 14056 1420
rect 14004 1377 14013 1411
rect 14013 1377 14047 1411
rect 14047 1377 14056 1411
rect 14004 1368 14056 1377
rect 15660 1368 15712 1420
rect 18328 1368 18380 1420
rect 12072 1343 12124 1352
rect 12072 1309 12081 1343
rect 12081 1309 12115 1343
rect 12115 1309 12124 1343
rect 12072 1300 12124 1309
rect 12624 1300 12676 1352
rect 14096 1300 14148 1352
rect 16304 1343 16356 1352
rect 16304 1309 16313 1343
rect 16313 1309 16347 1343
rect 16347 1309 16356 1343
rect 16304 1300 16356 1309
rect 9404 1164 9456 1216
rect 9588 1164 9640 1216
rect 10692 1164 10744 1216
rect 11428 1232 11480 1284
rect 13176 1232 13228 1284
rect 13360 1232 13412 1284
rect 13912 1275 13964 1284
rect 13912 1241 13921 1275
rect 13921 1241 13955 1275
rect 13955 1241 13964 1275
rect 13912 1232 13964 1241
rect 15108 1232 15160 1284
rect 15568 1232 15620 1284
rect 16212 1232 16264 1284
rect 13636 1207 13688 1216
rect 13636 1173 13645 1207
rect 13645 1173 13679 1207
rect 13679 1173 13688 1207
rect 13636 1164 13688 1173
rect 15936 1164 15988 1216
rect 5028 1062 5080 1114
rect 5092 1062 5144 1114
rect 5156 1062 5208 1114
rect 5220 1062 5272 1114
rect 5284 1062 5336 1114
rect 8128 1062 8180 1114
rect 8192 1062 8244 1114
rect 8256 1062 8308 1114
rect 8320 1062 8372 1114
rect 8384 1062 8436 1114
rect 11228 1062 11280 1114
rect 11292 1062 11344 1114
rect 11356 1062 11408 1114
rect 11420 1062 11472 1114
rect 11484 1062 11536 1114
rect 14328 1062 14380 1114
rect 14392 1062 14444 1114
rect 14456 1062 14508 1114
rect 14520 1062 14572 1114
rect 14584 1062 14636 1114
rect 17428 1062 17480 1114
rect 17492 1062 17544 1114
rect 17556 1062 17608 1114
rect 17620 1062 17672 1114
rect 17684 1062 17736 1114
rect 7288 1003 7340 1012
rect 3976 892 4028 944
rect 4712 867 4764 876
rect 4712 833 4721 867
rect 4721 833 4755 867
rect 4755 833 4764 867
rect 4712 824 4764 833
rect 5632 892 5684 944
rect 5908 892 5960 944
rect 7288 969 7297 1003
rect 7297 969 7331 1003
rect 7331 969 7340 1003
rect 7288 960 7340 969
rect 8024 960 8076 1012
rect 8668 1003 8720 1012
rect 3976 756 4028 808
rect 4988 756 5040 808
rect 5816 799 5868 808
rect 5172 620 5224 672
rect 5816 765 5825 799
rect 5825 765 5859 799
rect 5859 765 5868 799
rect 5816 756 5868 765
rect 7932 824 7984 876
rect 8668 969 8677 1003
rect 8677 969 8711 1003
rect 8711 969 8720 1003
rect 8668 960 8720 969
rect 9404 1003 9456 1012
rect 9404 969 9413 1003
rect 9413 969 9447 1003
rect 9447 969 9456 1003
rect 9404 960 9456 969
rect 9496 1003 9548 1012
rect 9496 969 9505 1003
rect 9505 969 9539 1003
rect 9539 969 9548 1003
rect 9496 960 9548 969
rect 11612 960 11664 1012
rect 12624 1003 12676 1012
rect 10692 935 10744 944
rect 10692 901 10701 935
rect 10701 901 10735 935
rect 10735 901 10744 935
rect 10692 892 10744 901
rect 11152 892 11204 944
rect 12624 969 12633 1003
rect 12633 969 12667 1003
rect 12667 969 12676 1003
rect 12624 960 12676 969
rect 13360 1003 13412 1012
rect 13360 969 13369 1003
rect 13369 969 13403 1003
rect 13403 969 13412 1003
rect 13360 960 13412 969
rect 13728 960 13780 1012
rect 14740 960 14792 1012
rect 15108 1003 15160 1012
rect 15108 969 15117 1003
rect 15117 969 15151 1003
rect 15151 969 15160 1003
rect 17224 1003 17276 1012
rect 15108 960 15160 969
rect 17224 969 17233 1003
rect 17233 969 17267 1003
rect 17267 969 17276 1003
rect 17224 960 17276 969
rect 18236 1003 18288 1012
rect 18236 969 18245 1003
rect 18245 969 18279 1003
rect 18279 969 18288 1003
rect 18236 960 18288 969
rect 13452 892 13504 944
rect 14832 935 14884 944
rect 14832 901 14841 935
rect 14841 901 14875 935
rect 14875 901 14884 935
rect 14832 892 14884 901
rect 15016 935 15068 944
rect 15016 901 15025 935
rect 15025 901 15059 935
rect 15059 901 15068 935
rect 15016 892 15068 901
rect 15936 892 15988 944
rect 17868 892 17920 944
rect 12532 867 12584 876
rect 8852 756 8904 808
rect 12532 833 12541 867
rect 12541 833 12575 867
rect 12575 833 12584 867
rect 12532 824 12584 833
rect 13544 824 13596 876
rect 13636 824 13688 876
rect 13820 824 13872 876
rect 14372 824 14424 876
rect 17592 867 17644 876
rect 17592 833 17601 867
rect 17601 833 17635 867
rect 17635 833 17644 867
rect 17592 824 17644 833
rect 9312 756 9364 808
rect 10784 756 10836 808
rect 14188 799 14240 808
rect 14188 765 14197 799
rect 14197 765 14231 799
rect 14231 765 14240 799
rect 14188 756 14240 765
rect 14740 756 14792 808
rect 15476 799 15528 808
rect 7932 688 7984 740
rect 8944 688 8996 740
rect 5448 620 5500 672
rect 8116 620 8168 672
rect 9036 663 9088 672
rect 9036 629 9045 663
rect 9045 629 9079 663
rect 9079 629 9088 663
rect 9036 620 9088 629
rect 14096 620 14148 672
rect 15476 765 15485 799
rect 15485 765 15519 799
rect 15519 765 15528 799
rect 15476 756 15528 765
rect 16672 756 16724 808
rect 16948 731 17000 740
rect 16948 697 16957 731
rect 16957 697 16991 731
rect 16991 697 17000 731
rect 16948 688 17000 697
rect 15660 620 15712 672
rect 3478 518 3530 570
rect 3542 518 3594 570
rect 3606 518 3658 570
rect 3670 518 3722 570
rect 3734 518 3786 570
rect 6578 518 6630 570
rect 6642 518 6694 570
rect 6706 518 6758 570
rect 6770 518 6822 570
rect 6834 518 6886 570
rect 9678 518 9730 570
rect 9742 518 9794 570
rect 9806 518 9858 570
rect 9870 518 9922 570
rect 9934 518 9986 570
rect 12778 518 12830 570
rect 12842 518 12894 570
rect 12906 518 12958 570
rect 12970 518 13022 570
rect 13034 518 13086 570
rect 15878 518 15930 570
rect 15942 518 15994 570
rect 16006 518 16058 570
rect 16070 518 16122 570
rect 16134 518 16186 570
rect 4988 459 5040 468
rect 4988 425 4997 459
rect 4997 425 5031 459
rect 5031 425 5040 459
rect 4988 416 5040 425
rect 5816 459 5868 468
rect 5816 425 5825 459
rect 5825 425 5859 459
rect 5859 425 5868 459
rect 5816 416 5868 425
rect 4620 348 4672 400
rect 5172 348 5224 400
rect 6368 416 6420 468
rect 6460 416 6512 468
rect 8484 416 8536 468
rect 13176 416 13228 468
rect 15200 416 15252 468
rect 15476 416 15528 468
rect 17592 416 17644 468
rect 18052 459 18104 468
rect 18052 425 18061 459
rect 18061 425 18095 459
rect 18095 425 18104 459
rect 18052 416 18104 425
rect 18512 459 18564 468
rect 18512 425 18521 459
rect 18521 425 18555 459
rect 18555 425 18564 459
rect 18512 416 18564 425
rect 9588 348 9640 400
rect 13912 348 13964 400
rect 14924 348 14976 400
rect 16948 348 17000 400
rect 6092 280 6144 332
rect 6460 280 6512 332
rect 7932 280 7984 332
rect 8116 323 8168 332
rect 8116 289 8125 323
rect 8125 289 8159 323
rect 8159 289 8168 323
rect 8116 280 8168 289
rect 8944 323 8996 332
rect 8944 289 8953 323
rect 8953 289 8987 323
rect 8987 289 8996 323
rect 8944 280 8996 289
rect 15108 323 15160 332
rect 15108 289 15117 323
rect 15117 289 15151 323
rect 15151 289 15160 323
rect 15108 280 15160 289
rect 15292 280 15344 332
rect 5080 255 5132 264
rect 5080 221 5089 255
rect 5089 221 5123 255
rect 5123 221 5132 255
rect 5080 212 5132 221
rect 5908 212 5960 264
rect 6828 212 6880 264
rect 8024 255 8076 264
rect 8024 221 8033 255
rect 8033 221 8067 255
rect 8067 221 8076 255
rect 8024 212 8076 221
rect 8852 212 8904 264
rect 12532 212 12584 264
rect 4804 144 4856 196
rect 6460 187 6512 196
rect 6460 153 6469 187
rect 6469 153 6503 187
rect 6503 153 6512 187
rect 6460 144 6512 153
rect 13912 212 13964 264
rect 14188 212 14240 264
rect 16212 212 16264 264
rect 18512 212 18564 264
rect 5448 76 5500 128
rect 13544 144 13596 196
rect 5028 -26 5080 26
rect 5092 -26 5144 26
rect 5156 -26 5208 26
rect 5220 -26 5272 26
rect 5284 -26 5336 26
rect 8128 -26 8180 26
rect 8192 -26 8244 26
rect 8256 -26 8308 26
rect 8320 -26 8372 26
rect 8384 -26 8436 26
rect 11228 -26 11280 26
rect 11292 -26 11344 26
rect 11356 -26 11408 26
rect 11420 -26 11472 26
rect 11484 -26 11536 26
rect 14328 -26 14380 26
rect 14392 -26 14444 26
rect 14456 -26 14508 26
rect 14520 -26 14572 26
rect 14584 -26 14636 26
rect 17428 -26 17480 26
rect 17492 -26 17544 26
rect 17556 -26 17608 26
rect 17620 -26 17672 26
rect 17684 -26 17736 26
<< metal2 >>
rect 1398 11200 1454 12000
rect 4250 11200 4306 12000
rect 6840 11206 7052 11234
rect 664 10668 716 10674
rect 664 10610 716 10616
rect 676 9586 704 10610
rect 940 9920 992 9926
rect 940 9862 992 9868
rect 952 9654 980 9862
rect 940 9648 992 9654
rect 940 9590 992 9596
rect 664 9580 716 9586
rect 664 9522 716 9528
rect 676 8498 704 9522
rect 1412 9178 1440 11200
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 2056 10130 2084 10406
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 1688 9722 1716 10066
rect 2424 9926 2452 10610
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2504 10056 2556 10062
rect 2608 10044 2636 10406
rect 2700 10266 2728 10474
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2556 10016 2636 10044
rect 2504 9998 2556 10004
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 2424 9518 2452 9862
rect 2608 9654 2636 10016
rect 2596 9648 2648 9654
rect 2596 9590 2648 9596
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2516 9450 2544 9522
rect 2700 9450 2728 10202
rect 2976 10130 3004 10406
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 2688 9444 2740 9450
rect 2688 9386 2740 9392
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 2516 9110 2544 9386
rect 2792 9330 2820 9930
rect 2964 9648 3016 9654
rect 3068 9636 3096 10610
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3016 9608 3096 9636
rect 2964 9590 3016 9596
rect 3068 9382 3096 9608
rect 3160 9586 3188 10066
rect 3252 9722 3280 10542
rect 3478 10364 3786 10384
rect 3478 10362 3484 10364
rect 3540 10362 3564 10364
rect 3620 10362 3644 10364
rect 3700 10362 3724 10364
rect 3780 10362 3786 10364
rect 3540 10310 3542 10362
rect 3722 10310 3724 10362
rect 3478 10308 3484 10310
rect 3540 10308 3564 10310
rect 3620 10308 3644 10310
rect 3700 10308 3724 10310
rect 3780 10308 3786 10310
rect 3478 10288 3786 10308
rect 4264 10266 4292 11200
rect 5028 10908 5336 10928
rect 5028 10906 5034 10908
rect 5090 10906 5114 10908
rect 5170 10906 5194 10908
rect 5250 10906 5274 10908
rect 5330 10906 5336 10908
rect 5090 10854 5092 10906
rect 5272 10854 5274 10906
rect 5028 10852 5034 10854
rect 5090 10852 5114 10854
rect 5170 10852 5194 10854
rect 5250 10852 5274 10854
rect 5330 10852 5336 10854
rect 5028 10832 5336 10852
rect 6840 10810 6868 11206
rect 7024 11098 7052 11206
rect 7102 11200 7158 12000
rect 9954 11200 10010 12000
rect 12806 11200 12862 12000
rect 15658 11200 15714 12000
rect 18510 11200 18566 12000
rect 18786 11248 18842 11257
rect 7116 11098 7144 11200
rect 7024 11070 7144 11098
rect 8128 10908 8436 10928
rect 8128 10906 8134 10908
rect 8190 10906 8214 10908
rect 8270 10906 8294 10908
rect 8350 10906 8374 10908
rect 8430 10906 8436 10908
rect 8190 10854 8192 10906
rect 8372 10854 8374 10906
rect 8128 10852 8134 10854
rect 8190 10852 8214 10854
rect 8270 10852 8294 10854
rect 8350 10852 8374 10854
rect 8430 10852 8436 10854
rect 8128 10832 8436 10852
rect 9968 10810 9996 11200
rect 11228 10908 11536 10928
rect 11228 10906 11234 10908
rect 11290 10906 11314 10908
rect 11370 10906 11394 10908
rect 11450 10906 11474 10908
rect 11530 10906 11536 10908
rect 11290 10854 11292 10906
rect 11472 10854 11474 10906
rect 11228 10852 11234 10854
rect 11290 10852 11314 10854
rect 11370 10852 11394 10854
rect 11450 10852 11474 10854
rect 11530 10852 11536 10854
rect 11228 10832 11536 10852
rect 12820 10826 12848 11200
rect 14328 10908 14636 10928
rect 14328 10906 14334 10908
rect 14390 10906 14414 10908
rect 14470 10906 14494 10908
rect 14550 10906 14574 10908
rect 14630 10906 14636 10908
rect 14390 10854 14392 10906
rect 14572 10854 14574 10906
rect 14328 10852 14334 10854
rect 14390 10852 14414 10854
rect 14470 10852 14494 10854
rect 14550 10852 14574 10854
rect 14630 10852 14636 10854
rect 14328 10832 14636 10852
rect 12820 10810 12940 10826
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 9956 10804 10008 10810
rect 12820 10804 12952 10810
rect 12820 10798 12900 10804
rect 9956 10746 10008 10752
rect 12900 10746 12952 10752
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4448 10130 4476 10406
rect 5276 10198 5304 10610
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 5460 9994 5488 10610
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8484 10532 8536 10538
rect 8484 10474 8536 10480
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 6578 10364 6886 10384
rect 6578 10362 6584 10364
rect 6640 10362 6664 10364
rect 6720 10362 6744 10364
rect 6800 10362 6824 10364
rect 6880 10362 6886 10364
rect 6640 10310 6642 10362
rect 6822 10310 6824 10362
rect 6578 10308 6584 10310
rect 6640 10308 6664 10310
rect 6720 10308 6744 10310
rect 6800 10308 6824 10310
rect 6880 10308 6886 10310
rect 6578 10288 6886 10308
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3804 9586 3832 9862
rect 5028 9820 5336 9840
rect 5028 9818 5034 9820
rect 5090 9818 5114 9820
rect 5170 9818 5194 9820
rect 5250 9818 5274 9820
rect 5330 9818 5336 9820
rect 5090 9766 5092 9818
rect 5272 9766 5274 9818
rect 5028 9764 5034 9766
rect 5090 9764 5114 9766
rect 5170 9764 5194 9766
rect 5250 9764 5274 9766
rect 5330 9764 5336 9766
rect 5028 9744 5336 9764
rect 5264 9648 5316 9654
rect 5264 9590 5316 9596
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 2872 9376 2924 9382
rect 2792 9324 2872 9330
rect 2792 9318 2924 9324
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2792 9302 2912 9318
rect 1492 9104 1544 9110
rect 1412 9052 1492 9058
rect 1412 9046 1544 9052
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 1308 9036 1360 9042
rect 1308 8978 1360 8984
rect 1412 9030 1532 9046
rect 1216 8832 1268 8838
rect 1216 8774 1268 8780
rect 1228 8566 1256 8774
rect 1320 8634 1348 8978
rect 1412 8974 1440 9030
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1308 8628 1360 8634
rect 1308 8570 1360 8576
rect 2516 8566 2544 9046
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 1216 8560 1268 8566
rect 1216 8502 1268 8508
rect 2504 8560 2556 8566
rect 2504 8502 2556 8508
rect 664 8492 716 8498
rect 664 8434 716 8440
rect 676 7410 704 8434
rect 2792 8430 2820 8978
rect 2884 8906 2912 9302
rect 3160 9042 3188 9522
rect 3252 9450 3280 9522
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3478 9276 3786 9296
rect 3478 9274 3484 9276
rect 3540 9274 3564 9276
rect 3620 9274 3644 9276
rect 3700 9274 3724 9276
rect 3780 9274 3786 9276
rect 3540 9222 3542 9274
rect 3722 9222 3724 9274
rect 3478 9220 3484 9222
rect 3540 9220 3564 9222
rect 3620 9220 3644 9222
rect 3700 9220 3724 9222
rect 3780 9220 3786 9222
rect 3478 9200 3786 9220
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 4080 8922 4108 9318
rect 4632 9178 4660 9454
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 3988 8906 4108 8922
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 5276 8922 5304 9590
rect 5368 9432 5396 9862
rect 5552 9654 5580 10066
rect 7300 10062 7328 10406
rect 8496 10266 8524 10474
rect 8588 10470 8616 10542
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6288 9722 6316 9862
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 5448 9444 5500 9450
rect 5368 9404 5448 9432
rect 5448 9386 5500 9392
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 3976 8900 4108 8906
rect 4028 8894 4108 8900
rect 3976 8842 4028 8848
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2884 8362 2912 8842
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3252 8634 3280 8774
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3344 8498 3372 8774
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 3068 8090 3096 8434
rect 3478 8188 3786 8208
rect 3478 8186 3484 8188
rect 3540 8186 3564 8188
rect 3620 8186 3644 8188
rect 3700 8186 3724 8188
rect 3780 8186 3786 8188
rect 3540 8134 3542 8186
rect 3722 8134 3724 8186
rect 3478 8132 3484 8134
rect 3540 8132 3564 8134
rect 3620 8132 3644 8134
rect 3700 8132 3724 8134
rect 3780 8132 3786 8134
rect 3478 8112 3786 8132
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 664 7404 716 7410
rect 664 7346 716 7352
rect 676 6914 704 7346
rect 1308 7336 1360 7342
rect 1308 7278 1360 7284
rect 676 6886 980 6914
rect 952 6798 980 6886
rect 940 6792 992 6798
rect 940 6734 992 6740
rect 952 5778 980 6734
rect 1320 6730 1348 7278
rect 1504 6798 1532 7822
rect 2240 7546 2268 7822
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2424 7478 2452 7686
rect 2412 7472 2464 7478
rect 2412 7414 2464 7420
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1964 6798 1992 7142
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1308 6724 1360 6730
rect 1308 6666 1360 6672
rect 1032 6656 1084 6662
rect 1032 6598 1084 6604
rect 1044 6322 1072 6598
rect 2056 6390 2084 7346
rect 2424 7002 2452 7414
rect 2608 7410 2636 7822
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2700 7546 2728 7754
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 3160 7410 3188 7822
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2976 6798 3004 7210
rect 3056 6928 3108 6934
rect 3056 6870 3108 6876
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2516 6458 2544 6734
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 3068 6390 3096 6870
rect 2044 6384 2096 6390
rect 2044 6326 2096 6332
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 1032 6316 1084 6322
rect 1032 6258 1084 6264
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 940 5772 992 5778
rect 940 5714 992 5720
rect 2792 5642 2820 6190
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2884 5914 2912 6054
rect 3068 5914 3096 6190
rect 3160 6186 3188 7346
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3252 6866 3280 7142
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3344 6780 3372 7822
rect 4080 7410 4108 8894
rect 4172 7954 4200 8910
rect 4908 8566 4936 8910
rect 5276 8894 5396 8922
rect 5028 8732 5336 8752
rect 5028 8730 5034 8732
rect 5090 8730 5114 8732
rect 5170 8730 5194 8732
rect 5250 8730 5274 8732
rect 5330 8730 5336 8732
rect 5090 8678 5092 8730
rect 5272 8678 5274 8730
rect 5028 8676 5034 8678
rect 5090 8676 5114 8678
rect 5170 8676 5194 8678
rect 5250 8676 5274 8678
rect 5330 8676 5336 8678
rect 5028 8656 5336 8676
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4172 7546 4200 7890
rect 4356 7818 4384 8366
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 3478 7100 3786 7120
rect 3478 7098 3484 7100
rect 3540 7098 3564 7100
rect 3620 7098 3644 7100
rect 3700 7098 3724 7100
rect 3780 7098 3786 7100
rect 3540 7046 3542 7098
rect 3722 7046 3724 7098
rect 3478 7044 3484 7046
rect 3540 7044 3564 7046
rect 3620 7044 3644 7046
rect 3700 7044 3724 7046
rect 3780 7044 3786 7046
rect 3478 7024 3786 7044
rect 3424 6792 3476 6798
rect 3344 6752 3424 6780
rect 3424 6734 3476 6740
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3528 6458 3556 6598
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3620 6186 3648 6734
rect 3804 6474 3832 6734
rect 3896 6730 3924 7210
rect 3988 6798 4016 7278
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3884 6724 3936 6730
rect 3884 6666 3936 6672
rect 3804 6446 3924 6474
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 3478 6012 3786 6032
rect 3478 6010 3484 6012
rect 3540 6010 3564 6012
rect 3620 6010 3644 6012
rect 3700 6010 3724 6012
rect 3780 6010 3786 6012
rect 3540 5958 3542 6010
rect 3722 5958 3724 6010
rect 3478 5956 3484 5958
rect 3540 5956 3564 5958
rect 3620 5956 3644 5958
rect 3700 5956 3724 5958
rect 3780 5956 3786 5958
rect 3478 5936 3786 5956
rect 3896 5914 3924 6446
rect 4080 6118 4108 7346
rect 4172 6798 4200 7482
rect 4724 7342 4752 7890
rect 4816 7886 4844 8230
rect 4908 8090 4936 8502
rect 5368 8498 5396 8894
rect 5460 8634 5488 9386
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 6012 8090 6040 9522
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6288 9042 6316 9318
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6184 8526 6236 8532
rect 6184 8468 6236 8474
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5028 7644 5336 7664
rect 5028 7642 5034 7644
rect 5090 7642 5114 7644
rect 5170 7642 5194 7644
rect 5250 7642 5274 7644
rect 5330 7642 5336 7644
rect 5090 7590 5092 7642
rect 5272 7590 5274 7642
rect 5028 7588 5034 7590
rect 5090 7588 5114 7590
rect 5170 7588 5194 7590
rect 5250 7588 5274 7590
rect 5330 7588 5336 7590
rect 5028 7568 5336 7588
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5276 6798 5304 7142
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5552 6730 5580 7686
rect 5920 7410 5948 7754
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5644 7206 5672 7346
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5644 6866 5672 7142
rect 5736 7002 5764 7278
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 2780 5636 2832 5642
rect 2780 5578 2832 5584
rect 4080 5574 4108 6054
rect 4816 5642 4844 6598
rect 5028 6556 5336 6576
rect 5028 6554 5034 6556
rect 5090 6554 5114 6556
rect 5170 6554 5194 6556
rect 5250 6554 5274 6556
rect 5330 6554 5336 6556
rect 5090 6502 5092 6554
rect 5272 6502 5274 6554
rect 5028 6500 5034 6502
rect 5090 6500 5114 6502
rect 5170 6500 5194 6502
rect 5250 6500 5274 6502
rect 5330 6500 5336 6502
rect 5028 6480 5336 6500
rect 5552 6322 5580 6666
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5736 6458 5764 6598
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5828 6322 5856 6802
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5920 6458 5948 6734
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 6012 6322 6040 8026
rect 6196 7546 6224 8468
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6288 7002 6316 8978
rect 6380 8838 6408 9522
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 6472 8974 6500 9318
rect 6578 9276 6886 9296
rect 6578 9274 6584 9276
rect 6640 9274 6664 9276
rect 6720 9274 6744 9276
rect 6800 9274 6824 9276
rect 6880 9274 6886 9276
rect 6640 9222 6642 9274
rect 6822 9222 6824 9274
rect 6578 9220 6584 9222
rect 6640 9220 6664 9222
rect 6720 9220 6744 9222
rect 6800 9220 6824 9222
rect 6880 9220 6886 9222
rect 6578 9200 6886 9220
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6380 8090 6408 8774
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6380 7886 6408 8026
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6472 7818 6500 8910
rect 7116 8906 7144 9318
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6578 8188 6886 8208
rect 6578 8186 6584 8188
rect 6640 8186 6664 8188
rect 6720 8186 6744 8188
rect 6800 8186 6824 8188
rect 6880 8186 6886 8188
rect 6640 8134 6642 8186
rect 6822 8134 6824 8186
rect 6578 8132 6584 8134
rect 6640 8132 6664 8134
rect 6720 8132 6744 8134
rect 6800 8132 6824 8134
rect 6880 8132 6886 8134
rect 6578 8112 6886 8132
rect 6828 8016 6880 8022
rect 6932 7970 6960 8230
rect 6880 7964 6960 7970
rect 6828 7958 6960 7964
rect 6840 7942 6960 7958
rect 7116 7954 7144 8298
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6460 7812 6512 7818
rect 6460 7754 6512 7760
rect 6472 7342 6500 7754
rect 6840 7546 6868 7822
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 4080 5370 4108 5510
rect 5028 5468 5336 5488
rect 5028 5466 5034 5468
rect 5090 5466 5114 5468
rect 5170 5466 5194 5468
rect 5250 5466 5274 5468
rect 5330 5466 5336 5468
rect 5090 5414 5092 5466
rect 5272 5414 5274 5466
rect 5028 5412 5034 5414
rect 5090 5412 5114 5414
rect 5170 5412 5194 5414
rect 5250 5412 5274 5414
rect 5330 5412 5336 5414
rect 5028 5392 5336 5412
rect 5552 5370 5580 5510
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 3478 4924 3786 4944
rect 3478 4922 3484 4924
rect 3540 4922 3564 4924
rect 3620 4922 3644 4924
rect 3700 4922 3724 4924
rect 3780 4922 3786 4924
rect 3540 4870 3542 4922
rect 3722 4870 3724 4922
rect 3478 4868 3484 4870
rect 3540 4868 3564 4870
rect 3620 4868 3644 4870
rect 3700 4868 3724 4870
rect 3780 4868 3786 4870
rect 3478 4848 3786 4868
rect 4080 4842 4108 5306
rect 5644 5234 5672 5850
rect 5828 5846 5856 6258
rect 6288 6254 6316 6938
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 5816 5840 5868 5846
rect 5816 5782 5868 5788
rect 6472 5778 6500 7278
rect 6578 7100 6886 7120
rect 6578 7098 6584 7100
rect 6640 7098 6664 7100
rect 6720 7098 6744 7100
rect 6800 7098 6824 7100
rect 6880 7098 6886 7100
rect 6640 7046 6642 7098
rect 6822 7046 6824 7098
rect 6578 7044 6584 7046
rect 6640 7044 6664 7046
rect 6720 7044 6744 7046
rect 6800 7044 6824 7046
rect 6880 7044 6886 7046
rect 6578 7024 6886 7044
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 7024 6458 7052 6802
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6578 6012 6886 6032
rect 6578 6010 6584 6012
rect 6640 6010 6664 6012
rect 6720 6010 6744 6012
rect 6800 6010 6824 6012
rect 6880 6010 6886 6012
rect 6640 5958 6642 6010
rect 6822 5958 6824 6010
rect 6578 5956 6584 5958
rect 6640 5956 6664 5958
rect 6720 5956 6744 5958
rect 6800 5956 6824 5958
rect 6880 5956 6886 5958
rect 6578 5936 6886 5956
rect 7208 5914 7236 9998
rect 8128 9820 8436 9840
rect 8128 9818 8134 9820
rect 8190 9818 8214 9820
rect 8270 9818 8294 9820
rect 8350 9818 8374 9820
rect 8430 9818 8436 9820
rect 8190 9766 8192 9818
rect 8372 9766 8374 9818
rect 8128 9764 8134 9766
rect 8190 9764 8214 9766
rect 8270 9764 8294 9766
rect 8350 9764 8374 9766
rect 8430 9764 8436 9766
rect 8128 9744 8436 9764
rect 8128 8732 8436 8752
rect 8128 8730 8134 8732
rect 8190 8730 8214 8732
rect 8270 8730 8294 8732
rect 8350 8730 8374 8732
rect 8430 8730 8436 8732
rect 8190 8678 8192 8730
rect 8372 8678 8374 8730
rect 8128 8676 8134 8678
rect 8190 8676 8214 8678
rect 8270 8676 8294 8678
rect 8350 8676 8374 8678
rect 8430 8676 8436 8678
rect 8128 8656 8436 8676
rect 8588 8566 8616 10406
rect 8772 10266 8800 10610
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8392 8560 8444 8566
rect 8312 8520 8392 8548
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7576 7274 7604 8434
rect 8312 8378 8340 8520
rect 8392 8502 8444 8508
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8220 8350 8340 8378
rect 8220 8294 8248 8350
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8220 7818 8248 8230
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 8496 7750 8524 8434
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8128 7644 8436 7664
rect 8128 7642 8134 7644
rect 8190 7642 8214 7644
rect 8270 7642 8294 7644
rect 8350 7642 8374 7644
rect 8430 7642 8436 7644
rect 8190 7590 8192 7642
rect 8372 7590 8374 7642
rect 8128 7588 8134 7590
rect 8190 7588 8214 7590
rect 8270 7588 8294 7590
rect 8350 7588 8374 7590
rect 8430 7588 8436 7590
rect 8128 7568 8436 7588
rect 8772 7546 8800 9522
rect 9140 8906 9168 10406
rect 9678 10364 9986 10384
rect 9678 10362 9684 10364
rect 9740 10362 9764 10364
rect 9820 10362 9844 10364
rect 9900 10362 9924 10364
rect 9980 10362 9986 10364
rect 9740 10310 9742 10362
rect 9922 10310 9924 10362
rect 9678 10308 9684 10310
rect 9740 10308 9764 10310
rect 9820 10308 9844 10310
rect 9900 10308 9924 10310
rect 9980 10308 9986 10310
rect 9678 10288 9986 10308
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 9678 9276 9986 9296
rect 9678 9274 9684 9276
rect 9740 9274 9764 9276
rect 9820 9274 9844 9276
rect 9900 9274 9924 9276
rect 9980 9274 9986 9276
rect 9740 9222 9742 9274
rect 9922 9222 9924 9274
rect 9678 9220 9684 9222
rect 9740 9220 9764 9222
rect 9820 9220 9844 9222
rect 9900 9220 9924 9222
rect 9980 9220 9986 9222
rect 9678 9200 9986 9220
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 8864 8498 8892 8774
rect 9232 8514 9260 8774
rect 9324 8634 9352 8774
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9600 8514 9628 9114
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 9232 8498 9812 8514
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 9220 8492 9824 8498
rect 9272 8486 9772 8492
rect 9220 8434 9272 8440
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7576 6730 7604 7210
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7392 6254 7420 6666
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7484 6322 7512 6598
rect 7576 6458 7604 6666
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7392 5846 7420 6190
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7024 5302 7052 5510
rect 7012 5296 7064 5302
rect 7012 5238 7064 5244
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 3896 4814 4108 4842
rect 940 4684 992 4690
rect 940 4626 992 4632
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 952 4214 980 4626
rect 1308 4616 1360 4622
rect 1308 4558 1360 4564
rect 940 4208 992 4214
rect 940 4150 992 4156
rect 1320 4078 1348 4558
rect 1308 4072 1360 4078
rect 1308 4014 1360 4020
rect 2148 3602 2176 4626
rect 3896 4554 3924 4814
rect 5644 4758 5672 5170
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5920 4826 5948 5102
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6578 4924 6886 4944
rect 6578 4922 6584 4924
rect 6640 4922 6664 4924
rect 6720 4922 6744 4924
rect 6800 4922 6824 4924
rect 6880 4922 6886 4924
rect 6640 4870 6642 4922
rect 6822 4870 6824 4922
rect 6578 4868 6584 4870
rect 6640 4868 6664 4870
rect 6720 4868 6744 4870
rect 6800 4868 6824 4870
rect 6880 4868 6886 4870
rect 6578 4848 6886 4868
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 4080 4622 4108 4694
rect 4068 4616 4120 4622
rect 4988 4616 5040 4622
rect 4068 4558 4120 4564
rect 4908 4576 4988 4604
rect 3884 4548 3936 4554
rect 3884 4490 3936 4496
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2792 4282 2820 4422
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2792 3942 2820 4082
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2136 3596 2188 3602
rect 2136 3538 2188 3544
rect 664 2508 716 2514
rect 664 2450 716 2456
rect 676 2106 704 2450
rect 1676 2304 1728 2310
rect 1676 2246 1728 2252
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 664 2100 716 2106
rect 664 2042 716 2048
rect 1688 1902 1716 2246
rect 2056 2038 2084 2246
rect 2148 2038 2176 3538
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 2424 3194 2452 3402
rect 2792 3398 2820 3878
rect 3478 3836 3786 3856
rect 3478 3834 3484 3836
rect 3540 3834 3564 3836
rect 3620 3834 3644 3836
rect 3700 3834 3724 3836
rect 3780 3834 3786 3836
rect 3540 3782 3542 3834
rect 3722 3782 3724 3834
rect 3478 3780 3484 3782
rect 3540 3780 3564 3782
rect 3620 3780 3644 3782
rect 3700 3780 3724 3782
rect 3780 3780 3786 3782
rect 3478 3760 3786 3780
rect 3896 3738 3924 4490
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3988 4214 4016 4422
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 4080 4146 4108 4558
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4448 4282 4476 4422
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4816 4078 4844 4422
rect 4908 4146 4936 4576
rect 4988 4558 5040 4564
rect 5028 4380 5336 4400
rect 5028 4378 5034 4380
rect 5090 4378 5114 4380
rect 5170 4378 5194 4380
rect 5250 4378 5274 4380
rect 5330 4378 5336 4380
rect 5090 4326 5092 4378
rect 5272 4326 5274 4378
rect 5028 4324 5034 4326
rect 5090 4324 5114 4326
rect 5170 4324 5194 4326
rect 5250 4324 5274 4326
rect 5330 4324 5336 4326
rect 5028 4304 5336 4324
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3896 3466 3924 3674
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 3884 3460 3936 3466
rect 3884 3402 3936 3408
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2792 3126 2820 3334
rect 4080 3126 4108 3470
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4356 3126 4384 3334
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 2792 2854 2820 3062
rect 4448 3058 4476 3538
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4724 3058 4752 3402
rect 5028 3292 5336 3312
rect 5028 3290 5034 3292
rect 5090 3290 5114 3292
rect 5170 3290 5194 3292
rect 5250 3290 5274 3292
rect 5330 3290 5336 3292
rect 5090 3238 5092 3290
rect 5272 3238 5274 3290
rect 5028 3236 5034 3238
rect 5090 3236 5114 3238
rect 5170 3236 5194 3238
rect 5250 3236 5274 3238
rect 5330 3236 5336 3238
rect 5028 3216 5336 3236
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2044 2032 2096 2038
rect 2044 1974 2096 1980
rect 2136 2032 2188 2038
rect 2516 2009 2544 2790
rect 2688 2508 2740 2514
rect 2688 2450 2740 2456
rect 2136 1974 2188 1980
rect 2502 2000 2558 2009
rect 1676 1896 1728 1902
rect 1676 1838 1728 1844
rect 2148 1426 2176 1974
rect 2700 1970 2728 2450
rect 2792 2310 2820 2790
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 2976 2106 3004 2382
rect 3068 2378 3096 2994
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 3056 2372 3108 2378
rect 3056 2314 3108 2320
rect 2964 2100 3016 2106
rect 2964 2042 3016 2048
rect 2502 1935 2504 1944
rect 2556 1935 2558 1944
rect 2688 1964 2740 1970
rect 2504 1906 2556 1912
rect 2688 1906 2740 1912
rect 3068 1834 3096 2314
rect 3160 1970 3188 2518
rect 3344 2514 3372 2994
rect 3516 2916 3568 2922
rect 3700 2916 3752 2922
rect 3568 2876 3700 2904
rect 3516 2858 3568 2864
rect 3700 2858 3752 2864
rect 3478 2748 3786 2768
rect 3478 2746 3484 2748
rect 3540 2746 3564 2748
rect 3620 2746 3644 2748
rect 3700 2746 3724 2748
rect 3780 2746 3786 2748
rect 3540 2694 3542 2746
rect 3722 2694 3724 2746
rect 3478 2692 3484 2694
rect 3540 2692 3564 2694
rect 3620 2692 3644 2694
rect 3700 2692 3724 2694
rect 3780 2692 3786 2694
rect 3478 2672 3786 2692
rect 3988 2650 4016 2994
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 3252 2038 3280 2382
rect 3608 2372 3660 2378
rect 3608 2314 3660 2320
rect 3620 2106 3648 2314
rect 3608 2100 3660 2106
rect 3608 2042 3660 2048
rect 3240 2032 3292 2038
rect 3240 1974 3292 1980
rect 3896 1970 3924 2382
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3148 1964 3200 1970
rect 3148 1906 3200 1912
rect 3608 1964 3660 1970
rect 3608 1906 3660 1912
rect 3884 1964 3936 1970
rect 3884 1906 3936 1912
rect 3056 1828 3108 1834
rect 3056 1770 3108 1776
rect 3516 1828 3568 1834
rect 3620 1816 3648 1906
rect 3568 1788 3648 1816
rect 3516 1770 3568 1776
rect 3988 1766 4016 2246
rect 4724 2009 4752 2994
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 4710 2000 4766 2009
rect 4908 1970 4936 2246
rect 5028 2204 5336 2224
rect 5028 2202 5034 2204
rect 5090 2202 5114 2204
rect 5170 2202 5194 2204
rect 5250 2202 5274 2204
rect 5330 2202 5336 2204
rect 5090 2150 5092 2202
rect 5272 2150 5274 2202
rect 5028 2148 5034 2150
rect 5090 2148 5114 2150
rect 5170 2148 5194 2150
rect 5250 2148 5274 2150
rect 5330 2148 5336 2150
rect 5028 2128 5336 2148
rect 4710 1935 4766 1944
rect 4896 1964 4948 1970
rect 4896 1906 4948 1912
rect 3976 1760 4028 1766
rect 3976 1702 4028 1708
rect 4712 1760 4764 1766
rect 4712 1702 4764 1708
rect 5356 1760 5408 1766
rect 5356 1702 5408 1708
rect 3478 1660 3786 1680
rect 3478 1658 3484 1660
rect 3540 1658 3564 1660
rect 3620 1658 3644 1660
rect 3700 1658 3724 1660
rect 3780 1658 3786 1660
rect 3540 1606 3542 1658
rect 3722 1606 3724 1658
rect 3478 1604 3484 1606
rect 3540 1604 3564 1606
rect 3620 1604 3644 1606
rect 3700 1604 3724 1606
rect 3780 1604 3786 1606
rect 3478 1584 3786 1604
rect 2136 1420 2188 1426
rect 2136 1362 2188 1368
rect 3988 1358 4016 1702
rect 3976 1352 4028 1358
rect 3976 1294 4028 1300
rect 4620 1352 4672 1358
rect 4620 1294 4672 1300
rect 3988 1222 4016 1294
rect 3976 1216 4028 1222
rect 3976 1158 4028 1164
rect 3988 950 4016 1158
rect 3976 944 4028 950
rect 3974 912 3976 921
rect 4028 912 4030 921
rect 3974 847 4030 856
rect 3988 814 4016 847
rect 3976 808 4028 814
rect 3976 750 4028 756
rect 3478 572 3786 592
rect 3478 570 3484 572
rect 3540 570 3564 572
rect 3620 570 3644 572
rect 3700 570 3724 572
rect 3780 570 3786 572
rect 3540 518 3542 570
rect 3722 518 3724 570
rect 3478 516 3484 518
rect 3540 516 3564 518
rect 3620 516 3644 518
rect 3700 516 3724 518
rect 3780 516 3786 518
rect 3478 496 3786 516
rect 4632 406 4660 1294
rect 4724 882 4752 1702
rect 5368 1426 5396 1702
rect 5460 1562 5488 2382
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5552 1970 5580 2246
rect 5644 2038 5672 4694
rect 6932 4690 6960 4966
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6932 4486 6960 4626
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6932 4146 6960 4422
rect 7116 4282 7144 4490
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5724 3120 5776 3126
rect 5724 3062 5776 3068
rect 5736 2378 5764 3062
rect 5828 3058 5856 3334
rect 6104 3058 6132 4082
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6380 3534 6408 3878
rect 6472 3738 6500 4014
rect 6578 3836 6886 3856
rect 6578 3834 6584 3836
rect 6640 3834 6664 3836
rect 6720 3834 6744 3836
rect 6800 3834 6824 3836
rect 6880 3834 6886 3836
rect 6640 3782 6642 3834
rect 6822 3782 6824 3834
rect 6578 3780 6584 3782
rect 6640 3780 6664 3782
rect 6720 3780 6744 3782
rect 6800 3780 6824 3782
rect 6880 3780 6886 3782
rect 6578 3760 6886 3780
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6932 3534 6960 4082
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 7208 3194 7236 5238
rect 7760 4146 7788 5850
rect 7852 5370 7880 6802
rect 7944 6186 7972 7278
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 8036 6798 8064 7142
rect 8404 6866 8432 7142
rect 8772 7002 8800 7346
rect 9140 7002 9168 7686
rect 9324 7410 9352 8486
rect 9772 8434 9824 8440
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 9678 8188 9986 8208
rect 9678 8186 9684 8188
rect 9740 8186 9764 8188
rect 9820 8186 9844 8188
rect 9900 8186 9924 8188
rect 9980 8186 9986 8188
rect 9740 8134 9742 8186
rect 9922 8134 9924 8186
rect 9678 8132 9684 8134
rect 9740 8132 9764 8134
rect 9820 8132 9844 8134
rect 9900 8132 9924 8134
rect 9980 8132 9986 8134
rect 9678 8112 9986 8132
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9508 7546 9536 8026
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8036 6186 8064 6734
rect 8128 6556 8436 6576
rect 8128 6554 8134 6556
rect 8190 6554 8214 6556
rect 8270 6554 8294 6556
rect 8350 6554 8374 6556
rect 8430 6554 8436 6556
rect 8190 6502 8192 6554
rect 8372 6502 8374 6554
rect 8128 6500 8134 6502
rect 8190 6500 8214 6502
rect 8270 6500 8294 6502
rect 8350 6500 8374 6502
rect 8430 6500 8436 6502
rect 8128 6480 8436 6500
rect 8496 6390 8524 6802
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 7932 5636 7984 5642
rect 7932 5578 7984 5584
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7944 5302 7972 5578
rect 8128 5468 8436 5488
rect 8128 5466 8134 5468
rect 8190 5466 8214 5468
rect 8270 5466 8294 5468
rect 8350 5466 8374 5468
rect 8430 5466 8436 5468
rect 8190 5414 8192 5466
rect 8372 5414 8374 5466
rect 8128 5412 8134 5414
rect 8190 5412 8214 5414
rect 8270 5412 8294 5414
rect 8350 5412 8374 5414
rect 8430 5412 8436 5414
rect 8128 5392 8436 5412
rect 7932 5296 7984 5302
rect 7932 5238 7984 5244
rect 7944 4826 7972 5238
rect 8496 5234 8524 6190
rect 8588 5710 8616 6598
rect 8956 6322 8984 6666
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8956 5166 8984 6258
rect 9232 6186 9260 7278
rect 9508 6662 9536 7482
rect 9600 7410 9628 7890
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9220 6180 9272 6186
rect 9220 6122 9272 6128
rect 9416 5370 9444 6598
rect 9600 6390 9628 7346
rect 9784 7342 9812 7958
rect 10060 7546 10088 8366
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10046 7440 10102 7449
rect 10046 7375 10048 7384
rect 10100 7375 10102 7384
rect 10048 7346 10100 7352
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9678 7100 9986 7120
rect 9678 7098 9684 7100
rect 9740 7098 9764 7100
rect 9820 7098 9844 7100
rect 9900 7098 9924 7100
rect 9980 7098 9986 7100
rect 9740 7046 9742 7098
rect 9922 7046 9924 7098
rect 9678 7044 9684 7046
rect 9740 7044 9764 7046
rect 9820 7044 9844 7046
rect 9900 7044 9924 7046
rect 9980 7044 9986 7046
rect 9678 7024 9986 7044
rect 10060 6458 10088 7346
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 9678 6012 9986 6032
rect 9678 6010 9684 6012
rect 9740 6010 9764 6012
rect 9820 6010 9844 6012
rect 9900 6010 9924 6012
rect 9980 6010 9986 6012
rect 9740 5958 9742 6010
rect 9922 5958 9924 6010
rect 9678 5956 9684 5958
rect 9740 5956 9764 5958
rect 9820 5956 9844 5958
rect 9900 5956 9924 5958
rect 9980 5956 9986 5958
rect 9678 5936 9986 5956
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9692 5302 9720 5714
rect 10152 5302 10180 8978
rect 10230 6896 10286 6905
rect 10230 6831 10286 6840
rect 10244 6798 10272 6831
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 10336 5166 10364 9454
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10428 8022 10456 8434
rect 10520 8294 10548 9318
rect 10796 9178 10824 9454
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 11072 9042 11100 9998
rect 11164 9722 11192 10610
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11992 10130 12020 10406
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11992 9994 12020 10066
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 11228 9820 11536 9840
rect 11228 9818 11234 9820
rect 11290 9818 11314 9820
rect 11370 9818 11394 9820
rect 11450 9818 11474 9820
rect 11530 9818 11536 9820
rect 11290 9766 11292 9818
rect 11472 9766 11474 9818
rect 11228 9764 11234 9766
rect 11290 9764 11314 9766
rect 11370 9764 11394 9766
rect 11450 9764 11474 9766
rect 11530 9764 11536 9766
rect 11228 9744 11536 9764
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11624 9586 11652 9930
rect 12452 9926 12480 10542
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12544 9586 12572 10678
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13188 10470 13216 10610
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 12778 10364 13086 10384
rect 12778 10362 12784 10364
rect 12840 10362 12864 10364
rect 12920 10362 12944 10364
rect 13000 10362 13024 10364
rect 13080 10362 13086 10364
rect 12840 10310 12842 10362
rect 13022 10310 13024 10362
rect 12778 10308 12784 10310
rect 12840 10308 12864 10310
rect 12920 10308 12944 10310
rect 13000 10308 13024 10310
rect 13080 10308 13086 10310
rect 12778 10288 13086 10308
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12636 9654 12664 10202
rect 13188 10130 13216 10406
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12820 9450 12848 9862
rect 13188 9602 13216 10066
rect 13096 9586 13216 9602
rect 13084 9580 13216 9586
rect 13136 9574 13216 9580
rect 13084 9522 13136 9528
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12778 9276 13086 9296
rect 12778 9274 12784 9276
rect 12840 9274 12864 9276
rect 12920 9274 12944 9276
rect 13000 9274 13024 9276
rect 13080 9274 13086 9276
rect 12840 9222 12842 9274
rect 13022 9222 13024 9274
rect 12778 9220 12784 9222
rect 12840 9220 12864 9222
rect 12920 9220 12944 9222
rect 13000 9220 13024 9222
rect 13080 9220 13086 9222
rect 12778 9200 13086 9220
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10796 8294 10824 8434
rect 10508 8288 10560 8294
rect 10508 8230 10560 8236
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10980 8090 11008 8230
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 11164 7954 11192 8910
rect 12084 8906 12296 8922
rect 11612 8900 11664 8906
rect 11612 8842 11664 8848
rect 12072 8900 12296 8906
rect 12124 8894 12296 8900
rect 12072 8842 12124 8848
rect 11228 8732 11536 8752
rect 11228 8730 11234 8732
rect 11290 8730 11314 8732
rect 11370 8730 11394 8732
rect 11450 8730 11474 8732
rect 11530 8730 11536 8732
rect 11290 8678 11292 8730
rect 11472 8678 11474 8730
rect 11228 8676 11234 8678
rect 11290 8676 11314 8678
rect 11370 8676 11394 8678
rect 11450 8676 11474 8678
rect 11530 8676 11536 8678
rect 11228 8656 11536 8676
rect 11624 8634 11652 8842
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10416 7472 10468 7478
rect 10414 7440 10416 7449
rect 10468 7440 10470 7449
rect 10414 7375 10470 7384
rect 10598 7440 10654 7449
rect 10876 7404 10928 7410
rect 10654 7384 10732 7392
rect 10598 7375 10600 7384
rect 10652 7364 10732 7384
rect 10600 7346 10652 7352
rect 10414 7304 10470 7313
rect 10414 7239 10470 7248
rect 10428 6934 10456 7239
rect 10704 6934 10732 7364
rect 10876 7346 10928 7352
rect 10416 6928 10468 6934
rect 10692 6928 10744 6934
rect 10416 6870 10468 6876
rect 10690 6896 10692 6905
rect 10744 6896 10746 6905
rect 10690 6831 10746 6840
rect 10888 6798 10916 7346
rect 11072 7002 11100 7822
rect 11256 7732 11284 8434
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11348 7993 11376 8230
rect 11334 7984 11390 7993
rect 11624 7970 11652 8366
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11624 7942 11744 7970
rect 11334 7919 11390 7928
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11164 7704 11284 7732
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 10876 6792 10928 6798
rect 10414 6760 10470 6769
rect 11060 6792 11112 6798
rect 10876 6734 10928 6740
rect 11058 6760 11060 6769
rect 11112 6760 11114 6769
rect 10414 6695 10416 6704
rect 10468 6695 10470 6704
rect 11058 6695 11114 6704
rect 10416 6666 10468 6672
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10796 6458 10824 6598
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 11164 6322 11192 7704
rect 11228 7644 11536 7664
rect 11228 7642 11234 7644
rect 11290 7642 11314 7644
rect 11370 7642 11394 7644
rect 11450 7642 11474 7644
rect 11530 7642 11536 7644
rect 11290 7590 11292 7642
rect 11472 7590 11474 7642
rect 11228 7588 11234 7590
rect 11290 7588 11314 7590
rect 11370 7588 11394 7590
rect 11450 7588 11474 7590
rect 11530 7588 11536 7590
rect 11228 7568 11536 7588
rect 11624 7546 11652 7822
rect 11716 7546 11744 7942
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11808 7410 11836 8230
rect 11900 7546 11928 8366
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 12084 7478 12112 8230
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11348 7206 11376 7346
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11348 6730 11376 7142
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 11228 6556 11536 6576
rect 11228 6554 11234 6556
rect 11290 6554 11314 6556
rect 11370 6554 11394 6556
rect 11450 6554 11474 6556
rect 11530 6554 11536 6556
rect 11290 6502 11292 6554
rect 11472 6502 11474 6554
rect 11228 6500 11234 6502
rect 11290 6500 11314 6502
rect 11370 6500 11394 6502
rect 11450 6500 11474 6502
rect 11530 6500 11536 6502
rect 11228 6480 11536 6500
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 12176 6254 12204 8774
rect 12268 7800 12296 8894
rect 12778 8188 13086 8208
rect 12778 8186 12784 8188
rect 12840 8186 12864 8188
rect 12920 8186 12944 8188
rect 13000 8186 13024 8188
rect 13080 8186 13086 8188
rect 12840 8134 12842 8186
rect 13022 8134 13024 8186
rect 12778 8132 12784 8134
rect 12840 8132 12864 8134
rect 12920 8132 12944 8134
rect 13000 8132 13024 8134
rect 13080 8132 13086 8134
rect 12778 8112 13086 8132
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12348 7812 12400 7818
rect 12268 7772 12348 7800
rect 12348 7754 12400 7760
rect 12256 7200 12308 7206
rect 12360 7188 12388 7754
rect 12820 7410 12848 7822
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12716 7336 12768 7342
rect 12714 7304 12716 7313
rect 12768 7304 12770 7313
rect 12714 7239 12770 7248
rect 12308 7160 12388 7188
rect 12256 7142 12308 7148
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 11072 6118 11100 6190
rect 11520 6180 11572 6186
rect 11520 6122 11572 6128
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11532 5642 11560 6122
rect 12268 5642 12296 7142
rect 12778 7100 13086 7120
rect 12778 7098 12784 7100
rect 12840 7098 12864 7100
rect 12920 7098 12944 7100
rect 13000 7098 13024 7100
rect 13080 7098 13086 7100
rect 12840 7046 12842 7098
rect 13022 7046 13024 7098
rect 12778 7044 12784 7046
rect 12840 7044 12864 7046
rect 12920 7044 12944 7046
rect 13000 7044 13024 7046
rect 13080 7044 13086 7046
rect 12778 7024 13086 7044
rect 12992 6928 13044 6934
rect 12992 6870 13044 6876
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12636 5846 12664 6734
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12820 6458 12848 6598
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 13004 6254 13032 6870
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 12778 6012 13086 6032
rect 12778 6010 12784 6012
rect 12840 6010 12864 6012
rect 12920 6010 12944 6012
rect 13000 6010 13024 6012
rect 13080 6010 13086 6012
rect 12840 5958 12842 6010
rect 13022 5958 13024 6010
rect 12778 5956 12784 5958
rect 12840 5956 12864 5958
rect 12920 5956 12944 5958
rect 13000 5956 13024 5958
rect 13080 5956 13086 5958
rect 12778 5936 13086 5956
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 11520 5636 11572 5642
rect 11520 5578 11572 5584
rect 12256 5636 12308 5642
rect 12256 5578 12308 5584
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10428 5234 10456 5510
rect 11228 5468 11536 5488
rect 11228 5466 11234 5468
rect 11290 5466 11314 5468
rect 11370 5466 11394 5468
rect 11450 5466 11474 5468
rect 11530 5466 11536 5468
rect 11290 5414 11292 5466
rect 11472 5414 11474 5466
rect 11228 5412 11234 5414
rect 11290 5412 11314 5414
rect 11370 5412 11394 5414
rect 11450 5412 11474 5414
rect 11530 5412 11536 5414
rect 11228 5392 11536 5412
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 9678 4924 9986 4944
rect 9678 4922 9684 4924
rect 9740 4922 9764 4924
rect 9820 4922 9844 4924
rect 9900 4922 9924 4924
rect 9980 4922 9986 4924
rect 9740 4870 9742 4922
rect 9922 4870 9924 4922
rect 9678 4868 9684 4870
rect 9740 4868 9764 4870
rect 9820 4868 9844 4870
rect 9900 4868 9924 4870
rect 9980 4868 9986 4870
rect 9678 4848 9986 4868
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7944 3738 7972 4626
rect 8128 4380 8436 4400
rect 8128 4378 8134 4380
rect 8190 4378 8214 4380
rect 8270 4378 8294 4380
rect 8350 4378 8374 4380
rect 8430 4378 8436 4380
rect 8190 4326 8192 4378
rect 8372 4326 8374 4378
rect 8128 4324 8134 4326
rect 8190 4324 8214 4326
rect 8270 4324 8294 4326
rect 8350 4324 8374 4326
rect 8430 4324 8436 4326
rect 8128 4304 8436 4324
rect 9416 4214 9444 4762
rect 10428 4690 10456 5170
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10704 4282 10732 5306
rect 12268 5302 12296 5578
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 12268 4690 12296 5238
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12636 4690 12664 5170
rect 13188 5166 13216 5510
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 12778 4924 13086 4944
rect 12778 4922 12784 4924
rect 12840 4922 12864 4924
rect 12920 4922 12944 4924
rect 13000 4922 13024 4924
rect 13080 4922 13086 4924
rect 12840 4870 12842 4922
rect 13022 4870 13024 4922
rect 12778 4868 12784 4870
rect 12840 4868 12864 4870
rect 12920 4868 12944 4870
rect 13000 4868 13024 4870
rect 13080 4868 13086 4870
rect 12778 4848 13086 4868
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 12268 4554 12296 4626
rect 13280 4622 13308 10542
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 14016 9518 14044 10406
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 14108 9722 14136 9998
rect 15304 9926 15332 10406
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 14328 9820 14636 9840
rect 14328 9818 14334 9820
rect 14390 9818 14414 9820
rect 14470 9818 14494 9820
rect 14550 9818 14574 9820
rect 14630 9818 14636 9820
rect 14390 9766 14392 9818
rect 14572 9766 14574 9818
rect 14328 9764 14334 9766
rect 14390 9764 14414 9766
rect 14470 9764 14494 9766
rect 14550 9764 14574 9766
rect 14630 9764 14636 9766
rect 14328 9744 14636 9764
rect 14096 9716 14148 9722
rect 14096 9658 14148 9664
rect 15304 9674 15332 9862
rect 15304 9654 15608 9674
rect 14188 9648 14240 9654
rect 15304 9648 15620 9654
rect 15304 9646 15568 9648
rect 14188 9590 14240 9596
rect 15568 9590 15620 9596
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14108 9042 14136 9318
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14108 8566 14136 8978
rect 14200 8838 14228 9590
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14384 8906 14412 9318
rect 14844 9178 14872 9454
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 14372 8900 14424 8906
rect 14372 8842 14424 8848
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13832 8378 13860 8434
rect 13832 8350 13952 8378
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13464 7954 13492 8230
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13464 7818 13492 7890
rect 13452 7812 13504 7818
rect 13452 7754 13504 7760
rect 13464 7002 13492 7754
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13740 7274 13768 7686
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13372 5370 13400 6598
rect 13464 5778 13492 6938
rect 13924 6866 13952 8350
rect 14108 8022 14136 8502
rect 14200 8294 14228 8774
rect 14328 8732 14636 8752
rect 14328 8730 14334 8732
rect 14390 8730 14414 8732
rect 14470 8730 14494 8732
rect 14550 8730 14574 8732
rect 14630 8730 14636 8732
rect 14390 8678 14392 8730
rect 14572 8678 14574 8730
rect 14328 8676 14334 8678
rect 14390 8676 14414 8678
rect 14470 8676 14494 8678
rect 14550 8676 14574 8678
rect 14630 8676 14636 8678
rect 14328 8656 14636 8676
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 14096 8016 14148 8022
rect 14096 7958 14148 7964
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14016 7449 14044 7822
rect 14200 7546 14228 7822
rect 14328 7644 14636 7664
rect 14328 7642 14334 7644
rect 14390 7642 14414 7644
rect 14470 7642 14494 7644
rect 14550 7642 14574 7644
rect 14630 7642 14636 7644
rect 14390 7590 14392 7642
rect 14572 7590 14574 7642
rect 14328 7588 14334 7590
rect 14390 7588 14414 7590
rect 14470 7588 14494 7590
rect 14550 7588 14574 7590
rect 14630 7588 14636 7590
rect 14328 7568 14636 7588
rect 14752 7546 14780 7890
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14002 7440 14058 7449
rect 14002 7375 14058 7384
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 13924 6474 13952 6802
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 13832 6458 13952 6474
rect 14016 6458 14044 6734
rect 13820 6452 13952 6458
rect 13872 6446 13952 6452
rect 14004 6452 14056 6458
rect 13820 6394 13872 6400
rect 14004 6394 14056 6400
rect 14108 6322 14136 7142
rect 14292 6746 14320 7346
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14200 6718 14320 6746
rect 14384 6730 14412 7142
rect 14476 6866 14504 7346
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14372 6724 14424 6730
rect 14200 6390 14228 6718
rect 14372 6666 14424 6672
rect 14328 6556 14636 6576
rect 14328 6554 14334 6556
rect 14390 6554 14414 6556
rect 14470 6554 14494 6556
rect 14550 6554 14574 6556
rect 14630 6554 14636 6556
rect 14390 6502 14392 6554
rect 14572 6502 14574 6554
rect 14328 6500 14334 6502
rect 14390 6500 14414 6502
rect 14470 6500 14494 6502
rect 14550 6500 14574 6502
rect 14630 6500 14636 6502
rect 14328 6480 14636 6500
rect 14188 6384 14240 6390
rect 14188 6326 14240 6332
rect 14752 6322 14780 7482
rect 14844 7426 14872 9114
rect 15580 8566 15608 9590
rect 15568 8560 15620 8566
rect 15568 8502 15620 8508
rect 15384 8288 15436 8294
rect 15580 8276 15608 8502
rect 15436 8248 15608 8276
rect 15384 8230 15436 8236
rect 15106 7984 15162 7993
rect 14924 7948 14976 7954
rect 15106 7919 15162 7928
rect 14924 7890 14976 7896
rect 14936 7546 14964 7890
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 15120 7478 15148 7919
rect 15396 7886 15424 8230
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15108 7472 15160 7478
rect 14844 7410 14964 7426
rect 15108 7414 15160 7420
rect 14844 7404 14976 7410
rect 14844 7398 14924 7404
rect 14924 7346 14976 7352
rect 14832 7268 14884 7274
rect 14832 7210 14884 7216
rect 14844 6458 14872 7210
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14936 6254 14964 7346
rect 15212 6934 15240 7686
rect 15396 7478 15424 7822
rect 15384 7472 15436 7478
rect 15384 7414 15436 7420
rect 15396 7206 15424 7414
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15200 6928 15252 6934
rect 15200 6870 15252 6876
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 13452 5772 13504 5778
rect 13452 5714 13504 5720
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13464 5302 13492 5714
rect 14476 5710 14504 6122
rect 15028 6066 15056 6802
rect 15212 6322 15240 6870
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 14844 6038 15056 6066
rect 14844 5778 14872 6038
rect 15488 5846 15516 6190
rect 15672 5914 15700 11200
rect 17428 10908 17736 10928
rect 17428 10906 17434 10908
rect 17490 10906 17514 10908
rect 17570 10906 17594 10908
rect 17650 10906 17674 10908
rect 17730 10906 17736 10908
rect 17490 10854 17492 10906
rect 17672 10854 17674 10906
rect 17428 10852 17434 10854
rect 17490 10852 17514 10854
rect 17570 10852 17594 10854
rect 17650 10852 17674 10854
rect 17730 10852 17736 10854
rect 17428 10832 17736 10852
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 15878 10364 16186 10384
rect 15878 10362 15884 10364
rect 15940 10362 15964 10364
rect 16020 10362 16044 10364
rect 16100 10362 16124 10364
rect 16180 10362 16186 10364
rect 15940 10310 15942 10362
rect 16122 10310 16124 10362
rect 15878 10308 15884 10310
rect 15940 10308 15964 10310
rect 16020 10308 16044 10310
rect 16100 10308 16124 10310
rect 16180 10308 16186 10310
rect 15878 10288 16186 10308
rect 18064 10266 18092 10610
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17428 9820 17736 9840
rect 17428 9818 17434 9820
rect 17490 9818 17514 9820
rect 17570 9818 17594 9820
rect 17650 9818 17674 9820
rect 17730 9818 17736 9820
rect 17490 9766 17492 9818
rect 17672 9766 17674 9818
rect 17428 9764 17434 9766
rect 17490 9764 17514 9766
rect 17570 9764 17594 9766
rect 17650 9764 17674 9766
rect 17730 9764 17736 9766
rect 17428 9744 17736 9764
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 15878 9276 16186 9296
rect 15878 9274 15884 9276
rect 15940 9274 15964 9276
rect 16020 9274 16044 9276
rect 16100 9274 16124 9276
rect 16180 9274 16186 9276
rect 15940 9222 15942 9274
rect 16122 9222 16124 9274
rect 15878 9220 15884 9222
rect 15940 9220 15964 9222
rect 16020 9220 16044 9222
rect 16100 9220 16124 9222
rect 16180 9220 16186 9222
rect 15878 9200 16186 9220
rect 16592 9178 16620 9454
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16868 9042 16896 9454
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16408 8634 16436 8910
rect 17132 8900 17184 8906
rect 17132 8842 17184 8848
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 17144 8362 17172 8842
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 17428 8732 17736 8752
rect 17428 8730 17434 8732
rect 17490 8730 17514 8732
rect 17570 8730 17594 8732
rect 17650 8730 17674 8732
rect 17730 8730 17736 8732
rect 17490 8678 17492 8730
rect 17672 8678 17674 8730
rect 17428 8676 17434 8678
rect 17490 8676 17514 8678
rect 17570 8676 17594 8678
rect 17650 8676 17674 8678
rect 17730 8676 17736 8678
rect 17428 8656 17736 8676
rect 18156 8566 18184 8774
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 15878 8188 16186 8208
rect 15878 8186 15884 8188
rect 15940 8186 15964 8188
rect 16020 8186 16044 8188
rect 16100 8186 16124 8188
rect 16180 8186 16186 8188
rect 15940 8134 15942 8186
rect 16122 8134 16124 8186
rect 15878 8132 15884 8134
rect 15940 8132 15964 8134
rect 16020 8132 16044 8134
rect 16100 8132 16124 8134
rect 16180 8132 16186 8134
rect 15878 8112 16186 8132
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 16120 7744 16172 7750
rect 16120 7686 16172 7692
rect 16132 7546 16160 7686
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 15878 7100 16186 7120
rect 15878 7098 15884 7100
rect 15940 7098 15964 7100
rect 16020 7098 16044 7100
rect 16100 7098 16124 7100
rect 16180 7098 16186 7100
rect 15940 7046 15942 7098
rect 16122 7046 16124 7098
rect 15878 7044 15884 7046
rect 15940 7044 15964 7046
rect 16020 7044 16044 7046
rect 16100 7044 16124 7046
rect 16180 7044 16186 7046
rect 15878 7024 16186 7044
rect 16408 7002 16436 7754
rect 16672 7336 16724 7342
rect 16868 7324 16896 8230
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 17052 7410 17080 7890
rect 17144 7818 17172 8298
rect 18524 8090 18552 11200
rect 18786 11183 18842 11192
rect 18800 10810 18828 11183
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18694 9752 18750 9761
rect 18694 9687 18750 9696
rect 18708 9586 18736 9687
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18616 8265 18644 8298
rect 18602 8256 18658 8265
rect 18602 8191 18658 8200
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 17132 7812 17184 7818
rect 17132 7754 17184 7760
rect 17868 7812 17920 7818
rect 17868 7754 17920 7760
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16724 7296 16896 7324
rect 16672 7278 16724 7284
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 15764 6254 15792 6598
rect 16224 6458 16252 6598
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16316 6390 16344 6802
rect 16408 6798 16436 6938
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16304 6384 16356 6390
rect 16304 6326 16356 6332
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 14832 5772 14884 5778
rect 14832 5714 14884 5720
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14740 5636 14792 5642
rect 14740 5578 14792 5584
rect 14328 5468 14636 5488
rect 14328 5466 14334 5468
rect 14390 5466 14414 5468
rect 14470 5466 14494 5468
rect 14550 5466 14574 5468
rect 14630 5466 14636 5468
rect 14390 5414 14392 5466
rect 14572 5414 14574 5466
rect 14328 5412 14334 5414
rect 14390 5412 14414 5414
rect 14470 5412 14494 5414
rect 14550 5412 14574 5414
rect 14630 5412 14636 5414
rect 14328 5392 14636 5412
rect 14752 5370 14780 5578
rect 14844 5574 14872 5714
rect 15764 5574 15792 6054
rect 15878 6012 16186 6032
rect 15878 6010 15884 6012
rect 15940 6010 15964 6012
rect 16020 6010 16044 6012
rect 16100 6010 16124 6012
rect 16180 6010 16186 6012
rect 15940 5958 15942 6010
rect 16122 5958 16124 6010
rect 15878 5956 15884 5958
rect 15940 5956 15964 5958
rect 16020 5956 16044 5958
rect 16100 5956 16124 5958
rect 16180 5956 16186 5958
rect 15878 5936 16186 5956
rect 16212 5636 16264 5642
rect 16212 5578 16264 5584
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 15752 5568 15804 5574
rect 15752 5510 15804 5516
rect 15844 5568 15896 5574
rect 15844 5510 15896 5516
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 13452 5296 13504 5302
rect 13452 5238 13504 5244
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 11228 4380 11536 4400
rect 11228 4378 11234 4380
rect 11290 4378 11314 4380
rect 11370 4378 11394 4380
rect 11450 4378 11474 4380
rect 11530 4378 11536 4380
rect 11290 4326 11292 4378
rect 11472 4326 11474 4378
rect 11228 4324 11234 4326
rect 11290 4324 11314 4326
rect 11370 4324 11394 4326
rect 11450 4324 11474 4326
rect 11530 4324 11536 4326
rect 11228 4304 11536 4324
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 7576 3534 7604 3674
rect 7555 3528 7607 3534
rect 7392 3488 7555 3516
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7392 3126 7420 3488
rect 7555 3470 7607 3476
rect 7944 3466 7972 3674
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7932 3052 7984 3058
rect 8036 3040 8064 3878
rect 8220 3738 8248 4014
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8128 3292 8436 3312
rect 8128 3290 8134 3292
rect 8190 3290 8214 3292
rect 8270 3290 8294 3292
rect 8350 3290 8374 3292
rect 8430 3290 8436 3292
rect 8190 3238 8192 3290
rect 8372 3238 8374 3290
rect 8128 3236 8134 3238
rect 8190 3236 8214 3238
rect 8270 3236 8294 3238
rect 8350 3236 8374 3238
rect 8430 3236 8436 3238
rect 8128 3216 8436 3236
rect 7984 3012 8064 3040
rect 7932 2994 7984 3000
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5828 2446 5856 2790
rect 6578 2748 6886 2768
rect 6578 2746 6584 2748
rect 6640 2746 6664 2748
rect 6720 2746 6744 2748
rect 6800 2746 6824 2748
rect 6880 2746 6886 2748
rect 6640 2694 6642 2746
rect 6822 2694 6824 2746
rect 6578 2692 6584 2694
rect 6640 2692 6664 2694
rect 6720 2692 6744 2694
rect 6800 2692 6824 2694
rect 6880 2692 6886 2694
rect 6578 2672 6886 2692
rect 5908 2576 5960 2582
rect 5908 2518 5960 2524
rect 6920 2576 6972 2582
rect 6920 2518 6972 2524
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 5632 2032 5684 2038
rect 5632 1974 5684 1980
rect 5540 1964 5592 1970
rect 5540 1906 5592 1912
rect 5448 1556 5500 1562
rect 5448 1498 5500 1504
rect 5356 1420 5408 1426
rect 5356 1362 5408 1368
rect 4804 1352 4856 1358
rect 4804 1294 4856 1300
rect 4816 1222 4844 1294
rect 4804 1216 4856 1222
rect 4804 1158 4856 1164
rect 4712 876 4764 882
rect 4712 818 4764 824
rect 4620 400 4672 406
rect 4620 342 4672 348
rect 4816 202 4844 1158
rect 5028 1116 5336 1136
rect 5028 1114 5034 1116
rect 5090 1114 5114 1116
rect 5170 1114 5194 1116
rect 5250 1114 5274 1116
rect 5330 1114 5336 1116
rect 5090 1062 5092 1114
rect 5272 1062 5274 1114
rect 5028 1060 5034 1062
rect 5090 1060 5114 1062
rect 5170 1060 5194 1062
rect 5250 1060 5274 1062
rect 5330 1060 5336 1062
rect 5028 1040 5336 1060
rect 5644 950 5672 1974
rect 5736 1426 5764 2314
rect 5920 2310 5948 2518
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 6012 1970 6040 2382
rect 6000 1964 6052 1970
rect 6000 1906 6052 1912
rect 6368 1896 6420 1902
rect 6368 1838 6420 1844
rect 5724 1420 5776 1426
rect 5724 1362 5776 1368
rect 6380 1358 6408 1838
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 6092 1216 6144 1222
rect 6092 1158 6144 1164
rect 5632 944 5684 950
rect 5908 944 5960 950
rect 5632 886 5684 892
rect 5906 912 5908 921
rect 5960 912 5962 921
rect 5906 847 5962 856
rect 4988 808 5040 814
rect 4988 750 5040 756
rect 5816 808 5868 814
rect 5816 750 5868 756
rect 5000 474 5028 750
rect 5172 672 5224 678
rect 5172 614 5224 620
rect 5448 672 5500 678
rect 5448 614 5500 620
rect 4988 468 5040 474
rect 4988 410 5040 416
rect 5184 406 5212 614
rect 5172 400 5224 406
rect 5078 368 5134 377
rect 5172 342 5224 348
rect 5078 303 5134 312
rect 5092 270 5120 303
rect 5080 264 5132 270
rect 5080 206 5132 212
rect 4804 196 4856 202
rect 4804 138 4856 144
rect 5460 134 5488 614
rect 5828 474 5856 750
rect 5816 468 5868 474
rect 5816 410 5868 416
rect 5920 270 5948 847
rect 6104 338 6132 1158
rect 6380 474 6408 1294
rect 6472 474 6500 2382
rect 6932 2038 6960 2518
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 6920 2032 6972 2038
rect 6920 1974 6972 1980
rect 7024 1766 7052 2382
rect 7116 2310 7144 2858
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7012 1760 7064 1766
rect 7012 1702 7064 1708
rect 6578 1660 6886 1680
rect 6578 1658 6584 1660
rect 6640 1658 6664 1660
rect 6720 1658 6744 1660
rect 6800 1658 6824 1660
rect 6880 1658 6886 1660
rect 6640 1606 6642 1658
rect 6822 1606 6824 1658
rect 6578 1604 6584 1606
rect 6640 1604 6664 1606
rect 6720 1604 6744 1606
rect 6800 1604 6824 1606
rect 6880 1604 6886 1606
rect 6578 1584 6886 1604
rect 7208 1222 7236 2994
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 7288 2916 7340 2922
rect 7288 2858 7340 2864
rect 7300 2582 7328 2858
rect 7288 2576 7340 2582
rect 7288 2518 7340 2524
rect 7484 2446 7512 2926
rect 7656 2848 7708 2854
rect 7656 2790 7708 2796
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7300 2106 7328 2382
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 7668 1970 7696 2790
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 7656 1964 7708 1970
rect 7656 1906 7708 1912
rect 7944 1562 7972 2382
rect 8128 2204 8436 2224
rect 8128 2202 8134 2204
rect 8190 2202 8214 2204
rect 8270 2202 8294 2204
rect 8350 2202 8374 2204
rect 8430 2202 8436 2204
rect 8190 2150 8192 2202
rect 8372 2150 8374 2202
rect 8128 2148 8134 2150
rect 8190 2148 8214 2150
rect 8270 2148 8294 2150
rect 8350 2148 8374 2150
rect 8430 2148 8436 2150
rect 8128 2128 8436 2148
rect 8588 2122 8616 2926
rect 8864 2514 8892 3470
rect 9416 3210 9444 4150
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10060 3942 10088 4082
rect 10704 4078 10732 4218
rect 12268 4214 12296 4490
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 9678 3836 9986 3856
rect 9678 3834 9684 3836
rect 9740 3834 9764 3836
rect 9820 3834 9844 3836
rect 9900 3834 9924 3836
rect 9980 3834 9986 3836
rect 9740 3782 9742 3834
rect 9922 3782 9924 3834
rect 9678 3780 9684 3782
rect 9740 3780 9764 3782
rect 9820 3780 9844 3782
rect 9900 3780 9924 3782
rect 9980 3780 9986 3782
rect 9678 3760 9986 3780
rect 10060 3602 10088 3878
rect 10244 3670 10272 3878
rect 10232 3664 10284 3670
rect 10232 3606 10284 3612
rect 10704 3602 10732 4014
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 9232 3182 9444 3210
rect 10232 3188 10284 3194
rect 9232 3126 9260 3182
rect 10284 3148 10364 3176
rect 10232 3130 10284 3136
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 9678 2748 9986 2768
rect 9678 2746 9684 2748
rect 9740 2746 9764 2748
rect 9820 2746 9844 2748
rect 9900 2746 9924 2748
rect 9980 2746 9986 2748
rect 9740 2694 9742 2746
rect 9922 2694 9924 2746
rect 9678 2692 9684 2694
rect 9740 2692 9764 2694
rect 9820 2692 9844 2694
rect 9900 2692 9924 2694
rect 9980 2692 9986 2694
rect 9678 2672 9986 2692
rect 10060 2514 10088 2994
rect 8852 2508 8904 2514
rect 8852 2450 8904 2456
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 8496 2106 8616 2122
rect 8484 2100 8616 2106
rect 8536 2094 8616 2100
rect 8484 2042 8536 2048
rect 8864 2038 8892 2450
rect 10244 2378 10272 2994
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 8852 2032 8904 2038
rect 8852 1974 8904 1980
rect 8116 1964 8168 1970
rect 8168 1924 8340 1952
rect 8116 1906 8168 1912
rect 7932 1556 7984 1562
rect 7932 1498 7984 1504
rect 7944 1426 7972 1498
rect 8312 1494 8340 1924
rect 10244 1902 10272 2314
rect 10336 2310 10364 3148
rect 10428 3058 10456 3334
rect 10520 3194 10548 3470
rect 10600 3460 10652 3466
rect 10600 3402 10652 3408
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 10336 2106 10364 2246
rect 10324 2100 10376 2106
rect 10324 2042 10376 2048
rect 10232 1896 10284 1902
rect 10232 1838 10284 1844
rect 9220 1760 9272 1766
rect 9220 1702 9272 1708
rect 9496 1760 9548 1766
rect 9496 1702 9548 1708
rect 9588 1760 9640 1766
rect 9588 1702 9640 1708
rect 9232 1562 9260 1702
rect 9220 1556 9272 1562
rect 9220 1498 9272 1504
rect 8300 1488 8352 1494
rect 8300 1430 8352 1436
rect 9312 1488 9364 1494
rect 9312 1430 9364 1436
rect 7932 1420 7984 1426
rect 7932 1362 7984 1368
rect 8668 1420 8720 1426
rect 8668 1362 8720 1368
rect 7288 1352 7340 1358
rect 8208 1352 8260 1358
rect 7288 1294 7340 1300
rect 8206 1320 8208 1329
rect 8260 1320 8262 1329
rect 6920 1216 6972 1222
rect 6920 1158 6972 1164
rect 7196 1216 7248 1222
rect 7196 1158 7248 1164
rect 6578 572 6886 592
rect 6578 570 6584 572
rect 6640 570 6664 572
rect 6720 570 6744 572
rect 6800 570 6824 572
rect 6880 570 6886 572
rect 6640 518 6642 570
rect 6822 518 6824 570
rect 6578 516 6584 518
rect 6640 516 6664 518
rect 6720 516 6744 518
rect 6800 516 6824 518
rect 6880 516 6886 518
rect 6578 496 6886 516
rect 6368 468 6420 474
rect 6368 410 6420 416
rect 6460 468 6512 474
rect 6460 410 6512 416
rect 6092 332 6144 338
rect 6092 274 6144 280
rect 6460 332 6512 338
rect 6460 274 6512 280
rect 5908 264 5960 270
rect 5908 206 5960 212
rect 6472 202 6500 274
rect 6828 264 6880 270
rect 6932 252 6960 1158
rect 7300 1018 7328 1294
rect 8206 1255 8262 1264
rect 8484 1284 8536 1290
rect 8484 1226 8536 1232
rect 8128 1116 8436 1136
rect 8128 1114 8134 1116
rect 8190 1114 8214 1116
rect 8270 1114 8294 1116
rect 8350 1114 8374 1116
rect 8430 1114 8436 1116
rect 8190 1062 8192 1114
rect 8372 1062 8374 1114
rect 8128 1060 8134 1062
rect 8190 1060 8214 1062
rect 8270 1060 8294 1062
rect 8350 1060 8374 1062
rect 8430 1060 8436 1062
rect 8128 1040 8436 1060
rect 7288 1012 7340 1018
rect 7288 954 7340 960
rect 8024 1012 8076 1018
rect 8024 954 8076 960
rect 7932 876 7984 882
rect 7932 818 7984 824
rect 7944 746 7972 818
rect 7932 740 7984 746
rect 7932 682 7984 688
rect 7944 338 7972 682
rect 7932 332 7984 338
rect 7932 274 7984 280
rect 8036 270 8064 954
rect 8116 672 8168 678
rect 8116 614 8168 620
rect 8128 338 8156 614
rect 8496 474 8524 1226
rect 8680 1018 8708 1362
rect 8668 1012 8720 1018
rect 8668 954 8720 960
rect 9324 814 9352 1430
rect 9404 1216 9456 1222
rect 9404 1158 9456 1164
rect 9416 1018 9444 1158
rect 9508 1018 9536 1702
rect 9600 1494 9628 1702
rect 9678 1660 9986 1680
rect 9678 1658 9684 1660
rect 9740 1658 9764 1660
rect 9820 1658 9844 1660
rect 9900 1658 9924 1660
rect 9980 1658 9986 1660
rect 9740 1606 9742 1658
rect 9922 1606 9924 1658
rect 9678 1604 9684 1606
rect 9740 1604 9764 1606
rect 9820 1604 9844 1606
rect 9900 1604 9924 1606
rect 9980 1604 9986 1606
rect 9678 1584 9986 1604
rect 10336 1494 10364 2042
rect 10520 1970 10548 3130
rect 10508 1964 10560 1970
rect 10508 1906 10560 1912
rect 9588 1488 9640 1494
rect 9588 1430 9640 1436
rect 10324 1488 10376 1494
rect 10324 1430 10376 1436
rect 10612 1358 10640 3402
rect 10600 1352 10652 1358
rect 10600 1294 10652 1300
rect 10704 1306 10732 3538
rect 11256 3534 11284 4082
rect 12268 3942 12296 4150
rect 12728 4078 12756 4422
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 13280 3942 13308 4558
rect 13372 4078 13400 4558
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 11228 3292 11536 3312
rect 11228 3290 11234 3292
rect 11290 3290 11314 3292
rect 11370 3290 11394 3292
rect 11450 3290 11474 3292
rect 11530 3290 11536 3292
rect 11290 3238 11292 3290
rect 11472 3238 11474 3290
rect 11228 3236 11234 3238
rect 11290 3236 11314 3238
rect 11370 3236 11394 3238
rect 11450 3236 11474 3238
rect 11530 3236 11536 3238
rect 11228 3216 11536 3236
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 10796 2582 10824 2994
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 11072 2514 11100 2858
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 11072 1970 11100 2450
rect 11060 1964 11112 1970
rect 11164 1952 11192 2994
rect 11808 2650 11836 2994
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 11716 2378 11744 2518
rect 11704 2372 11756 2378
rect 11704 2314 11756 2320
rect 11228 2204 11536 2224
rect 11228 2202 11234 2204
rect 11290 2202 11314 2204
rect 11370 2202 11394 2204
rect 11450 2202 11474 2204
rect 11530 2202 11536 2204
rect 11290 2150 11292 2202
rect 11472 2150 11474 2202
rect 11228 2148 11234 2150
rect 11290 2148 11314 2150
rect 11370 2148 11394 2150
rect 11450 2148 11474 2150
rect 11530 2148 11536 2150
rect 11228 2128 11536 2148
rect 11244 1964 11296 1970
rect 11164 1924 11244 1952
rect 11060 1906 11112 1912
rect 11244 1906 11296 1912
rect 10968 1896 11020 1902
rect 10968 1838 11020 1844
rect 10980 1329 11008 1838
rect 11152 1760 11204 1766
rect 11152 1702 11204 1708
rect 10966 1320 11022 1329
rect 9588 1216 9640 1222
rect 9588 1158 9640 1164
rect 9404 1012 9456 1018
rect 9404 954 9456 960
rect 9496 1012 9548 1018
rect 9496 954 9548 960
rect 8852 808 8904 814
rect 8852 750 8904 756
rect 9312 808 9364 814
rect 9312 750 9364 756
rect 8484 468 8536 474
rect 8484 410 8536 416
rect 8116 332 8168 338
rect 8116 274 8168 280
rect 8864 270 8892 750
rect 8944 740 8996 746
rect 8944 682 8996 688
rect 8956 338 8984 682
rect 9036 672 9088 678
rect 9036 614 9088 620
rect 9048 377 9076 614
rect 9600 406 9628 1158
rect 10612 921 10640 1294
rect 10704 1278 10824 1306
rect 10692 1216 10744 1222
rect 10692 1158 10744 1164
rect 10704 950 10732 1158
rect 10692 944 10744 950
rect 10598 912 10654 921
rect 10692 886 10744 892
rect 10598 847 10654 856
rect 10796 814 10824 1278
rect 10966 1255 11022 1264
rect 11164 950 11192 1702
rect 11256 1358 11284 1906
rect 11716 1766 11744 2314
rect 11704 1760 11756 1766
rect 11704 1702 11756 1708
rect 12084 1358 12112 3470
rect 12268 2650 12296 3878
rect 12452 2990 12480 3878
rect 12778 3836 13086 3856
rect 12778 3834 12784 3836
rect 12840 3834 12864 3836
rect 12920 3834 12944 3836
rect 13000 3834 13024 3836
rect 13080 3834 13086 3836
rect 12840 3782 12842 3834
rect 13022 3782 13024 3834
rect 12778 3780 12784 3782
rect 12840 3780 12864 3782
rect 12920 3780 12944 3782
rect 13000 3780 13024 3782
rect 13080 3780 13086 3782
rect 12778 3760 13086 3780
rect 13280 3738 13308 3878
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13372 3618 13400 4014
rect 13280 3590 13400 3618
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12256 1760 12308 1766
rect 12256 1702 12308 1708
rect 12268 1426 12296 1702
rect 12452 1562 12480 2246
rect 12636 1970 12664 2790
rect 12778 2748 13086 2768
rect 12778 2746 12784 2748
rect 12840 2746 12864 2748
rect 12920 2746 12944 2748
rect 13000 2746 13024 2748
rect 13080 2746 13086 2748
rect 12840 2694 12842 2746
rect 13022 2694 13024 2746
rect 12778 2692 12784 2694
rect 12840 2692 12864 2694
rect 12920 2692 12944 2694
rect 13000 2692 13024 2694
rect 13080 2692 13086 2694
rect 12778 2672 13086 2692
rect 13084 2576 13136 2582
rect 13004 2524 13084 2530
rect 13004 2518 13136 2524
rect 13004 2502 13124 2518
rect 13004 2446 13032 2502
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 13188 2360 13216 3130
rect 13096 2332 13216 2360
rect 13096 1970 13124 2332
rect 12624 1964 12676 1970
rect 12624 1906 12676 1912
rect 13084 1964 13136 1970
rect 13084 1906 13136 1912
rect 12778 1660 13086 1680
rect 12778 1658 12784 1660
rect 12840 1658 12864 1660
rect 12920 1658 12944 1660
rect 13000 1658 13024 1660
rect 13080 1658 13086 1660
rect 12840 1606 12842 1658
rect 13022 1606 13024 1658
rect 12778 1604 12784 1606
rect 12840 1604 12864 1606
rect 12920 1604 12944 1606
rect 13000 1604 13024 1606
rect 13080 1604 13086 1606
rect 12778 1584 13086 1604
rect 12440 1556 12492 1562
rect 12440 1498 12492 1504
rect 12256 1420 12308 1426
rect 12256 1362 12308 1368
rect 13084 1420 13136 1426
rect 13280 1408 13308 3590
rect 13464 3534 13492 4490
rect 14108 3602 14136 4626
rect 15764 4554 15792 5510
rect 15856 5166 15884 5510
rect 16224 5234 16252 5578
rect 16316 5370 16344 6326
rect 16408 5846 16436 6734
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 16684 5658 16712 6598
rect 16868 6458 16896 7296
rect 17144 6730 17172 7754
rect 17428 7644 17736 7664
rect 17428 7642 17434 7644
rect 17490 7642 17514 7644
rect 17570 7642 17594 7644
rect 17650 7642 17674 7644
rect 17730 7642 17736 7644
rect 17490 7590 17492 7642
rect 17672 7590 17674 7642
rect 17428 7588 17434 7590
rect 17490 7588 17514 7590
rect 17570 7588 17594 7590
rect 17650 7588 17674 7590
rect 17730 7588 17736 7590
rect 17428 7568 17736 7588
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17236 6866 17264 7142
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17132 6724 17184 6730
rect 17132 6666 17184 6672
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16592 5630 16712 5658
rect 16764 5636 16816 5642
rect 16592 5574 16620 5630
rect 16764 5578 16816 5584
rect 16856 5636 16908 5642
rect 17144 5624 17172 6666
rect 17328 6186 17356 7346
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 17428 6556 17736 6576
rect 17428 6554 17434 6556
rect 17490 6554 17514 6556
rect 17570 6554 17594 6556
rect 17650 6554 17674 6556
rect 17730 6554 17736 6556
rect 17490 6502 17492 6554
rect 17672 6502 17674 6554
rect 17428 6500 17434 6502
rect 17490 6500 17514 6502
rect 17570 6500 17594 6502
rect 17650 6500 17674 6502
rect 17730 6500 17736 6502
rect 17428 6480 17736 6500
rect 17788 6458 17816 6802
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17880 6254 17908 7754
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18340 6458 18368 7278
rect 18510 6760 18566 6769
rect 18510 6695 18566 6704
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18524 6322 18552 6695
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17316 6180 17368 6186
rect 17316 6122 17368 6128
rect 17880 5914 17908 6190
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17224 5636 17276 5642
rect 17144 5596 17224 5624
rect 16856 5578 16908 5584
rect 17224 5578 17276 5584
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16592 5370 16620 5510
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16684 5234 16712 5510
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16776 5166 16804 5578
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 15878 4924 16186 4944
rect 15878 4922 15884 4924
rect 15940 4922 15964 4924
rect 16020 4922 16044 4924
rect 16100 4922 16124 4924
rect 16180 4922 16186 4924
rect 15940 4870 15942 4922
rect 16122 4870 16124 4922
rect 15878 4868 15884 4870
rect 15940 4868 15964 4870
rect 16020 4868 16044 4870
rect 16100 4868 16124 4870
rect 16180 4868 16186 4870
rect 15878 4848 16186 4868
rect 16868 4554 16896 5578
rect 17428 5468 17736 5488
rect 17428 5466 17434 5468
rect 17490 5466 17514 5468
rect 17570 5466 17594 5468
rect 17650 5466 17674 5468
rect 17730 5466 17736 5468
rect 17490 5414 17492 5466
rect 17672 5414 17674 5466
rect 17428 5412 17434 5414
rect 17490 5412 17514 5414
rect 17570 5412 17594 5414
rect 17650 5412 17674 5414
rect 17730 5412 17736 5414
rect 17428 5392 17736 5412
rect 18510 5264 18566 5273
rect 18510 5199 18512 5208
rect 18564 5199 18566 5208
rect 18512 5170 18564 5176
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 14188 4548 14240 4554
rect 14188 4490 14240 4496
rect 15752 4548 15804 4554
rect 15752 4490 15804 4496
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 14200 4282 14228 4490
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 14328 4380 14636 4400
rect 14328 4378 14334 4380
rect 14390 4378 14414 4380
rect 14470 4378 14494 4380
rect 14550 4378 14574 4380
rect 14630 4378 14636 4380
rect 14390 4326 14392 4378
rect 14572 4326 14574 4378
rect 14328 4324 14334 4326
rect 14390 4324 14414 4326
rect 14470 4324 14494 4326
rect 14550 4324 14574 4326
rect 14630 4324 14636 4326
rect 14328 4304 14636 4324
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 15488 4146 15516 4422
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13464 3058 13492 3470
rect 13740 3194 13768 3470
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13372 2106 13400 2382
rect 13360 2100 13412 2106
rect 13360 2042 13412 2048
rect 13136 1380 13308 1408
rect 13084 1362 13136 1368
rect 11244 1352 11296 1358
rect 12072 1352 12124 1358
rect 11244 1294 11296 1300
rect 11440 1290 11652 1306
rect 12072 1294 12124 1300
rect 12624 1352 12676 1358
rect 13096 1329 13124 1362
rect 12624 1294 12676 1300
rect 13082 1320 13138 1329
rect 11428 1284 11652 1290
rect 11480 1278 11652 1284
rect 11428 1226 11480 1232
rect 11228 1116 11536 1136
rect 11228 1114 11234 1116
rect 11290 1114 11314 1116
rect 11370 1114 11394 1116
rect 11450 1114 11474 1116
rect 11530 1114 11536 1116
rect 11290 1062 11292 1114
rect 11472 1062 11474 1114
rect 11228 1060 11234 1062
rect 11290 1060 11314 1062
rect 11370 1060 11394 1062
rect 11450 1060 11474 1062
rect 11530 1060 11536 1062
rect 11228 1040 11536 1060
rect 11624 1018 11652 1278
rect 12636 1018 12664 1294
rect 13082 1255 13138 1264
rect 13176 1284 13228 1290
rect 13176 1226 13228 1232
rect 13360 1284 13412 1290
rect 13360 1226 13412 1232
rect 11612 1012 11664 1018
rect 11612 954 11664 960
rect 12624 1012 12676 1018
rect 12624 954 12676 960
rect 11152 944 11204 950
rect 11152 886 11204 892
rect 12532 876 12584 882
rect 12532 818 12584 824
rect 10784 808 10836 814
rect 10784 750 10836 756
rect 9678 572 9986 592
rect 9678 570 9684 572
rect 9740 570 9764 572
rect 9820 570 9844 572
rect 9900 570 9924 572
rect 9980 570 9986 572
rect 9740 518 9742 570
rect 9922 518 9924 570
rect 9678 516 9684 518
rect 9740 516 9764 518
rect 9820 516 9844 518
rect 9900 516 9924 518
rect 9980 516 9986 518
rect 9678 496 9986 516
rect 9588 400 9640 406
rect 9034 368 9090 377
rect 8944 332 8996 338
rect 9588 342 9640 348
rect 9034 303 9090 312
rect 8944 274 8996 280
rect 12544 270 12572 818
rect 12778 572 13086 592
rect 12778 570 12784 572
rect 12840 570 12864 572
rect 12920 570 12944 572
rect 13000 570 13024 572
rect 13080 570 13086 572
rect 12840 518 12842 570
rect 13022 518 13024 570
rect 12778 516 12784 518
rect 12840 516 12864 518
rect 12920 516 12944 518
rect 13000 516 13024 518
rect 13080 516 13086 518
rect 12778 496 13086 516
rect 13188 474 13216 1226
rect 13372 1018 13400 1226
rect 13360 1012 13412 1018
rect 13360 954 13412 960
rect 13464 950 13492 2586
rect 14016 2530 14044 2994
rect 13832 2502 14044 2530
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 13556 2106 13584 2314
rect 13544 2100 13596 2106
rect 13544 2042 13596 2048
rect 13636 2100 13688 2106
rect 13636 2042 13688 2048
rect 13648 1986 13676 2042
rect 13556 1958 13676 1986
rect 13452 944 13504 950
rect 13452 886 13504 892
rect 13556 882 13584 1958
rect 13728 1896 13780 1902
rect 13648 1856 13728 1884
rect 13648 1222 13676 1856
rect 13728 1838 13780 1844
rect 13728 1556 13780 1562
rect 13728 1498 13780 1504
rect 13740 1426 13768 1498
rect 13728 1420 13780 1426
rect 13728 1362 13780 1368
rect 13636 1216 13688 1222
rect 13636 1158 13688 1164
rect 13648 882 13676 1158
rect 13740 1018 13768 1362
rect 13728 1012 13780 1018
rect 13728 954 13780 960
rect 13832 921 13860 2502
rect 14108 2378 14136 3538
rect 15212 3534 15240 3878
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15292 3460 15344 3466
rect 15292 3402 15344 3408
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 14328 3292 14636 3312
rect 14328 3290 14334 3292
rect 14390 3290 14414 3292
rect 14470 3290 14494 3292
rect 14550 3290 14574 3292
rect 14630 3290 14636 3292
rect 14390 3238 14392 3290
rect 14572 3238 14574 3290
rect 14328 3236 14334 3238
rect 14390 3236 14414 3238
rect 14470 3236 14494 3238
rect 14550 3236 14574 3238
rect 14630 3236 14636 3238
rect 14328 3216 14636 3236
rect 15212 3058 15240 3334
rect 15304 3194 15332 3402
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 14200 2514 14228 2790
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14568 2378 14596 2586
rect 14096 2372 14148 2378
rect 14016 2332 14096 2360
rect 14016 1426 14044 2332
rect 14096 2314 14148 2320
rect 14556 2372 14608 2378
rect 14556 2314 14608 2320
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14328 2204 14636 2224
rect 14328 2202 14334 2204
rect 14390 2202 14414 2204
rect 14470 2202 14494 2204
rect 14550 2202 14574 2204
rect 14630 2202 14636 2204
rect 14390 2150 14392 2202
rect 14572 2150 14574 2202
rect 14328 2148 14334 2150
rect 14390 2148 14414 2150
rect 14470 2148 14494 2150
rect 14550 2148 14574 2150
rect 14630 2148 14636 2150
rect 14328 2128 14636 2148
rect 14752 2038 14780 2246
rect 14740 2032 14792 2038
rect 14792 1992 14872 2020
rect 14740 1974 14792 1980
rect 14188 1964 14240 1970
rect 14188 1906 14240 1912
rect 14004 1420 14056 1426
rect 14004 1362 14056 1368
rect 14096 1352 14148 1358
rect 14096 1294 14148 1300
rect 13912 1284 13964 1290
rect 13912 1226 13964 1232
rect 13818 912 13874 921
rect 13544 876 13596 882
rect 13544 818 13596 824
rect 13636 876 13688 882
rect 13818 847 13820 856
rect 13636 818 13688 824
rect 13872 847 13874 856
rect 13820 818 13872 824
rect 13176 468 13228 474
rect 13176 410 13228 416
rect 6880 224 6960 252
rect 8024 264 8076 270
rect 6828 206 6880 212
rect 8024 206 8076 212
rect 8852 264 8904 270
rect 8852 206 8904 212
rect 12532 264 12584 270
rect 12532 206 12584 212
rect 13556 202 13584 818
rect 13832 787 13860 818
rect 13924 406 13952 1226
rect 14108 678 14136 1294
rect 14200 1000 14228 1906
rect 14740 1760 14792 1766
rect 14740 1702 14792 1708
rect 14328 1116 14636 1136
rect 14328 1114 14334 1116
rect 14390 1114 14414 1116
rect 14470 1114 14494 1116
rect 14550 1114 14574 1116
rect 14630 1114 14636 1116
rect 14390 1062 14392 1114
rect 14572 1062 14574 1114
rect 14328 1060 14334 1062
rect 14390 1060 14414 1062
rect 14470 1060 14494 1062
rect 14550 1060 14574 1062
rect 14630 1060 14636 1062
rect 14328 1040 14636 1060
rect 14752 1018 14780 1702
rect 14740 1012 14792 1018
rect 14200 972 14412 1000
rect 14384 882 14412 972
rect 14740 954 14792 960
rect 14844 950 14872 1992
rect 14924 1828 14976 1834
rect 14924 1770 14976 1776
rect 14832 944 14884 950
rect 14832 886 14884 892
rect 14372 876 14424 882
rect 14372 818 14424 824
rect 14188 808 14240 814
rect 14188 750 14240 756
rect 14740 808 14792 814
rect 14936 762 14964 1770
rect 15120 1290 15148 2586
rect 15304 2514 15332 3130
rect 15396 3058 15424 3946
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15488 3126 15516 3878
rect 15878 3836 16186 3856
rect 15878 3834 15884 3836
rect 15940 3834 15964 3836
rect 16020 3834 16044 3836
rect 16100 3834 16124 3836
rect 16180 3834 16186 3836
rect 15940 3782 15942 3834
rect 16122 3782 16124 3834
rect 15878 3780 15884 3782
rect 15940 3780 15964 3782
rect 16020 3780 16044 3782
rect 16100 3780 16124 3782
rect 16180 3780 16186 3782
rect 15878 3760 16186 3780
rect 16224 3466 16252 4422
rect 17428 4380 17736 4400
rect 17428 4378 17434 4380
rect 17490 4378 17514 4380
rect 17570 4378 17594 4380
rect 17650 4378 17674 4380
rect 17730 4378 17736 4380
rect 17490 4326 17492 4378
rect 17672 4326 17674 4378
rect 17428 4324 17434 4326
rect 17490 4324 17514 4326
rect 17570 4324 17594 4326
rect 17650 4324 17674 4326
rect 17730 4324 17736 4326
rect 17428 4304 17736 4324
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16316 3602 16344 3674
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 15672 3126 15700 3334
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 15660 3120 15712 3126
rect 15660 3062 15712 3068
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15764 2650 15792 3334
rect 16132 2990 16160 3334
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 15878 2748 16186 2768
rect 15878 2746 15884 2748
rect 15940 2746 15964 2748
rect 16020 2746 16044 2748
rect 16100 2746 16124 2748
rect 16180 2746 16186 2748
rect 15940 2694 15942 2746
rect 16122 2694 16124 2746
rect 15878 2692 15884 2694
rect 15940 2692 15964 2694
rect 16020 2692 16044 2694
rect 16100 2692 16124 2694
rect 16180 2692 16186 2694
rect 15878 2672 16186 2692
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15304 2038 15332 2450
rect 15844 2372 15896 2378
rect 15844 2314 15896 2320
rect 15568 2100 15620 2106
rect 15568 2042 15620 2048
rect 15292 2032 15344 2038
rect 15292 1974 15344 1980
rect 15292 1760 15344 1766
rect 15292 1702 15344 1708
rect 15108 1284 15160 1290
rect 15160 1244 15240 1272
rect 15108 1226 15160 1232
rect 15108 1012 15160 1018
rect 15108 954 15160 960
rect 15016 944 15068 950
rect 15016 886 15068 892
rect 14792 756 14964 762
rect 14740 750 14964 756
rect 14096 672 14148 678
rect 14096 614 14148 620
rect 13912 400 13964 406
rect 13912 342 13964 348
rect 13924 270 13952 342
rect 14200 270 14228 750
rect 14752 734 14964 750
rect 14924 400 14976 406
rect 15028 388 15056 886
rect 14976 360 15056 388
rect 14924 342 14976 348
rect 15120 338 15148 954
rect 15212 474 15240 1244
rect 15200 468 15252 474
rect 15200 410 15252 416
rect 15304 338 15332 1702
rect 15580 1290 15608 2042
rect 15856 1902 15884 2314
rect 15844 1896 15896 1902
rect 15844 1838 15896 1844
rect 15878 1660 16186 1680
rect 15878 1658 15884 1660
rect 15940 1658 15964 1660
rect 16020 1658 16044 1660
rect 16100 1658 16124 1660
rect 16180 1658 16186 1660
rect 15940 1606 15942 1658
rect 16122 1606 16124 1658
rect 15878 1604 15884 1606
rect 15940 1604 15964 1606
rect 16020 1604 16044 1606
rect 16100 1604 16124 1606
rect 16180 1604 16186 1606
rect 15878 1584 16186 1604
rect 15660 1420 15712 1426
rect 15660 1362 15712 1368
rect 15568 1284 15620 1290
rect 15568 1226 15620 1232
rect 15476 808 15528 814
rect 15476 750 15528 756
rect 15488 474 15516 750
rect 15672 678 15700 1362
rect 16316 1358 16344 3538
rect 16408 3398 16436 4082
rect 17880 3534 17908 4422
rect 17972 4282 18000 4558
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16500 3194 16528 3470
rect 17428 3292 17736 3312
rect 17428 3290 17434 3292
rect 17490 3290 17514 3292
rect 17570 3290 17594 3292
rect 17650 3290 17674 3292
rect 17730 3290 17736 3292
rect 17490 3238 17492 3290
rect 17672 3238 17674 3290
rect 17428 3236 17434 3238
rect 17490 3236 17514 3238
rect 17570 3236 17594 3238
rect 17650 3236 17674 3238
rect 17730 3236 17736 3238
rect 17428 3216 17736 3236
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16500 2774 16528 3130
rect 16500 2746 16620 2774
rect 16592 1902 16620 2746
rect 17960 2372 18012 2378
rect 17960 2314 18012 2320
rect 17428 2204 17736 2224
rect 17428 2202 17434 2204
rect 17490 2202 17514 2204
rect 17570 2202 17594 2204
rect 17650 2202 17674 2204
rect 17730 2202 17736 2204
rect 17490 2150 17492 2202
rect 17672 2150 17674 2202
rect 17428 2148 17434 2150
rect 17490 2148 17514 2150
rect 17570 2148 17594 2150
rect 17650 2148 17674 2150
rect 17730 2148 17736 2150
rect 17428 2128 17736 2148
rect 17224 1964 17276 1970
rect 17224 1906 17276 1912
rect 16580 1896 16632 1902
rect 16632 1844 16712 1850
rect 16580 1838 16712 1844
rect 16592 1822 16712 1838
rect 16304 1352 16356 1358
rect 16304 1294 16356 1300
rect 16212 1284 16264 1290
rect 16212 1226 16264 1232
rect 15936 1216 15988 1222
rect 15936 1158 15988 1164
rect 15948 950 15976 1158
rect 15936 944 15988 950
rect 15936 886 15988 892
rect 15660 672 15712 678
rect 15660 614 15712 620
rect 15878 572 16186 592
rect 15878 570 15884 572
rect 15940 570 15964 572
rect 16020 570 16044 572
rect 16100 570 16124 572
rect 16180 570 16186 572
rect 15940 518 15942 570
rect 16122 518 16124 570
rect 15878 516 15884 518
rect 15940 516 15964 518
rect 16020 516 16044 518
rect 16100 516 16124 518
rect 16180 516 16186 518
rect 15878 496 16186 516
rect 15476 468 15528 474
rect 15476 410 15528 416
rect 15108 332 15160 338
rect 15108 274 15160 280
rect 15292 332 15344 338
rect 15292 274 15344 280
rect 16224 270 16252 1226
rect 16684 814 16712 1822
rect 17236 1018 17264 1906
rect 17868 1896 17920 1902
rect 17868 1838 17920 1844
rect 17880 1562 17908 1838
rect 17972 1562 18000 2314
rect 18156 2106 18184 4966
rect 18340 4826 18368 4966
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 18248 3602 18276 4558
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18524 3777 18552 4082
rect 18510 3768 18566 3777
rect 18510 3703 18566 3712
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 18248 2514 18276 3538
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 18510 2272 18566 2281
rect 18510 2207 18566 2216
rect 18144 2100 18196 2106
rect 18144 2042 18196 2048
rect 18236 2032 18288 2038
rect 18236 1974 18288 1980
rect 18052 1964 18104 1970
rect 18052 1906 18104 1912
rect 17868 1556 17920 1562
rect 17868 1498 17920 1504
rect 17960 1556 18012 1562
rect 17960 1498 18012 1504
rect 17428 1116 17736 1136
rect 17428 1114 17434 1116
rect 17490 1114 17514 1116
rect 17570 1114 17594 1116
rect 17650 1114 17674 1116
rect 17730 1114 17736 1116
rect 17490 1062 17492 1114
rect 17672 1062 17674 1114
rect 17428 1060 17434 1062
rect 17490 1060 17514 1062
rect 17570 1060 17594 1062
rect 17650 1060 17674 1062
rect 17730 1060 17736 1062
rect 17428 1040 17736 1060
rect 17224 1012 17276 1018
rect 17224 954 17276 960
rect 17880 950 17908 1498
rect 17868 944 17920 950
rect 17868 886 17920 892
rect 17592 876 17644 882
rect 17592 818 17644 824
rect 16672 808 16724 814
rect 16672 750 16724 756
rect 16948 740 17000 746
rect 16948 682 17000 688
rect 16960 406 16988 682
rect 17604 474 17632 818
rect 18064 474 18092 1906
rect 18248 1018 18276 1974
rect 18524 1970 18552 2207
rect 18512 1964 18564 1970
rect 18512 1906 18564 1912
rect 18328 1760 18380 1766
rect 18328 1702 18380 1708
rect 18340 1426 18368 1702
rect 18524 1562 18552 1906
rect 18512 1556 18564 1562
rect 18512 1498 18564 1504
rect 18328 1420 18380 1426
rect 18328 1362 18380 1368
rect 18236 1012 18288 1018
rect 18236 954 18288 960
rect 18510 776 18566 785
rect 18510 711 18566 720
rect 18524 474 18552 711
rect 17592 468 17644 474
rect 17592 410 17644 416
rect 18052 468 18104 474
rect 18052 410 18104 416
rect 18512 468 18564 474
rect 18512 410 18564 416
rect 16948 400 17000 406
rect 16948 342 17000 348
rect 18524 270 18552 410
rect 13912 264 13964 270
rect 13912 206 13964 212
rect 14188 264 14240 270
rect 14188 206 14240 212
rect 16212 264 16264 270
rect 16212 206 16264 212
rect 18512 264 18564 270
rect 18512 206 18564 212
rect 6460 196 6512 202
rect 6460 138 6512 144
rect 13544 196 13596 202
rect 13544 138 13596 144
rect 5448 128 5500 134
rect 5448 70 5500 76
rect 5028 28 5336 48
rect 5028 26 5034 28
rect 5090 26 5114 28
rect 5170 26 5194 28
rect 5250 26 5274 28
rect 5330 26 5336 28
rect 5090 -26 5092 26
rect 5272 -26 5274 26
rect 5028 -28 5034 -26
rect 5090 -28 5114 -26
rect 5170 -28 5194 -26
rect 5250 -28 5274 -26
rect 5330 -28 5336 -26
rect 5028 -48 5336 -28
rect 8128 28 8436 48
rect 8128 26 8134 28
rect 8190 26 8214 28
rect 8270 26 8294 28
rect 8350 26 8374 28
rect 8430 26 8436 28
rect 8190 -26 8192 26
rect 8372 -26 8374 26
rect 8128 -28 8134 -26
rect 8190 -28 8214 -26
rect 8270 -28 8294 -26
rect 8350 -28 8374 -26
rect 8430 -28 8436 -26
rect 8128 -48 8436 -28
rect 11228 28 11536 48
rect 11228 26 11234 28
rect 11290 26 11314 28
rect 11370 26 11394 28
rect 11450 26 11474 28
rect 11530 26 11536 28
rect 11290 -26 11292 26
rect 11472 -26 11474 26
rect 11228 -28 11234 -26
rect 11290 -28 11314 -26
rect 11370 -28 11394 -26
rect 11450 -28 11474 -26
rect 11530 -28 11536 -26
rect 11228 -48 11536 -28
rect 14328 28 14636 48
rect 14328 26 14334 28
rect 14390 26 14414 28
rect 14470 26 14494 28
rect 14550 26 14574 28
rect 14630 26 14636 28
rect 14390 -26 14392 26
rect 14572 -26 14574 26
rect 14328 -28 14334 -26
rect 14390 -28 14414 -26
rect 14470 -28 14494 -26
rect 14550 -28 14574 -26
rect 14630 -28 14636 -26
rect 14328 -48 14636 -28
rect 17428 28 17736 48
rect 17428 26 17434 28
rect 17490 26 17514 28
rect 17570 26 17594 28
rect 17650 26 17674 28
rect 17730 26 17736 28
rect 17490 -26 17492 26
rect 17672 -26 17674 26
rect 17428 -28 17434 -26
rect 17490 -28 17514 -26
rect 17570 -28 17594 -26
rect 17650 -28 17674 -26
rect 17730 -28 17736 -26
rect 17428 -48 17736 -28
<< via2 >>
rect 3484 10362 3540 10364
rect 3564 10362 3620 10364
rect 3644 10362 3700 10364
rect 3724 10362 3780 10364
rect 3484 10310 3530 10362
rect 3530 10310 3540 10362
rect 3564 10310 3594 10362
rect 3594 10310 3606 10362
rect 3606 10310 3620 10362
rect 3644 10310 3658 10362
rect 3658 10310 3670 10362
rect 3670 10310 3700 10362
rect 3724 10310 3734 10362
rect 3734 10310 3780 10362
rect 3484 10308 3540 10310
rect 3564 10308 3620 10310
rect 3644 10308 3700 10310
rect 3724 10308 3780 10310
rect 5034 10906 5090 10908
rect 5114 10906 5170 10908
rect 5194 10906 5250 10908
rect 5274 10906 5330 10908
rect 5034 10854 5080 10906
rect 5080 10854 5090 10906
rect 5114 10854 5144 10906
rect 5144 10854 5156 10906
rect 5156 10854 5170 10906
rect 5194 10854 5208 10906
rect 5208 10854 5220 10906
rect 5220 10854 5250 10906
rect 5274 10854 5284 10906
rect 5284 10854 5330 10906
rect 5034 10852 5090 10854
rect 5114 10852 5170 10854
rect 5194 10852 5250 10854
rect 5274 10852 5330 10854
rect 8134 10906 8190 10908
rect 8214 10906 8270 10908
rect 8294 10906 8350 10908
rect 8374 10906 8430 10908
rect 8134 10854 8180 10906
rect 8180 10854 8190 10906
rect 8214 10854 8244 10906
rect 8244 10854 8256 10906
rect 8256 10854 8270 10906
rect 8294 10854 8308 10906
rect 8308 10854 8320 10906
rect 8320 10854 8350 10906
rect 8374 10854 8384 10906
rect 8384 10854 8430 10906
rect 8134 10852 8190 10854
rect 8214 10852 8270 10854
rect 8294 10852 8350 10854
rect 8374 10852 8430 10854
rect 11234 10906 11290 10908
rect 11314 10906 11370 10908
rect 11394 10906 11450 10908
rect 11474 10906 11530 10908
rect 11234 10854 11280 10906
rect 11280 10854 11290 10906
rect 11314 10854 11344 10906
rect 11344 10854 11356 10906
rect 11356 10854 11370 10906
rect 11394 10854 11408 10906
rect 11408 10854 11420 10906
rect 11420 10854 11450 10906
rect 11474 10854 11484 10906
rect 11484 10854 11530 10906
rect 11234 10852 11290 10854
rect 11314 10852 11370 10854
rect 11394 10852 11450 10854
rect 11474 10852 11530 10854
rect 14334 10906 14390 10908
rect 14414 10906 14470 10908
rect 14494 10906 14550 10908
rect 14574 10906 14630 10908
rect 14334 10854 14380 10906
rect 14380 10854 14390 10906
rect 14414 10854 14444 10906
rect 14444 10854 14456 10906
rect 14456 10854 14470 10906
rect 14494 10854 14508 10906
rect 14508 10854 14520 10906
rect 14520 10854 14550 10906
rect 14574 10854 14584 10906
rect 14584 10854 14630 10906
rect 14334 10852 14390 10854
rect 14414 10852 14470 10854
rect 14494 10852 14550 10854
rect 14574 10852 14630 10854
rect 6584 10362 6640 10364
rect 6664 10362 6720 10364
rect 6744 10362 6800 10364
rect 6824 10362 6880 10364
rect 6584 10310 6630 10362
rect 6630 10310 6640 10362
rect 6664 10310 6694 10362
rect 6694 10310 6706 10362
rect 6706 10310 6720 10362
rect 6744 10310 6758 10362
rect 6758 10310 6770 10362
rect 6770 10310 6800 10362
rect 6824 10310 6834 10362
rect 6834 10310 6880 10362
rect 6584 10308 6640 10310
rect 6664 10308 6720 10310
rect 6744 10308 6800 10310
rect 6824 10308 6880 10310
rect 5034 9818 5090 9820
rect 5114 9818 5170 9820
rect 5194 9818 5250 9820
rect 5274 9818 5330 9820
rect 5034 9766 5080 9818
rect 5080 9766 5090 9818
rect 5114 9766 5144 9818
rect 5144 9766 5156 9818
rect 5156 9766 5170 9818
rect 5194 9766 5208 9818
rect 5208 9766 5220 9818
rect 5220 9766 5250 9818
rect 5274 9766 5284 9818
rect 5284 9766 5330 9818
rect 5034 9764 5090 9766
rect 5114 9764 5170 9766
rect 5194 9764 5250 9766
rect 5274 9764 5330 9766
rect 3484 9274 3540 9276
rect 3564 9274 3620 9276
rect 3644 9274 3700 9276
rect 3724 9274 3780 9276
rect 3484 9222 3530 9274
rect 3530 9222 3540 9274
rect 3564 9222 3594 9274
rect 3594 9222 3606 9274
rect 3606 9222 3620 9274
rect 3644 9222 3658 9274
rect 3658 9222 3670 9274
rect 3670 9222 3700 9274
rect 3724 9222 3734 9274
rect 3734 9222 3780 9274
rect 3484 9220 3540 9222
rect 3564 9220 3620 9222
rect 3644 9220 3700 9222
rect 3724 9220 3780 9222
rect 3484 8186 3540 8188
rect 3564 8186 3620 8188
rect 3644 8186 3700 8188
rect 3724 8186 3780 8188
rect 3484 8134 3530 8186
rect 3530 8134 3540 8186
rect 3564 8134 3594 8186
rect 3594 8134 3606 8186
rect 3606 8134 3620 8186
rect 3644 8134 3658 8186
rect 3658 8134 3670 8186
rect 3670 8134 3700 8186
rect 3724 8134 3734 8186
rect 3734 8134 3780 8186
rect 3484 8132 3540 8134
rect 3564 8132 3620 8134
rect 3644 8132 3700 8134
rect 3724 8132 3780 8134
rect 5034 8730 5090 8732
rect 5114 8730 5170 8732
rect 5194 8730 5250 8732
rect 5274 8730 5330 8732
rect 5034 8678 5080 8730
rect 5080 8678 5090 8730
rect 5114 8678 5144 8730
rect 5144 8678 5156 8730
rect 5156 8678 5170 8730
rect 5194 8678 5208 8730
rect 5208 8678 5220 8730
rect 5220 8678 5250 8730
rect 5274 8678 5284 8730
rect 5284 8678 5330 8730
rect 5034 8676 5090 8678
rect 5114 8676 5170 8678
rect 5194 8676 5250 8678
rect 5274 8676 5330 8678
rect 3484 7098 3540 7100
rect 3564 7098 3620 7100
rect 3644 7098 3700 7100
rect 3724 7098 3780 7100
rect 3484 7046 3530 7098
rect 3530 7046 3540 7098
rect 3564 7046 3594 7098
rect 3594 7046 3606 7098
rect 3606 7046 3620 7098
rect 3644 7046 3658 7098
rect 3658 7046 3670 7098
rect 3670 7046 3700 7098
rect 3724 7046 3734 7098
rect 3734 7046 3780 7098
rect 3484 7044 3540 7046
rect 3564 7044 3620 7046
rect 3644 7044 3700 7046
rect 3724 7044 3780 7046
rect 3484 6010 3540 6012
rect 3564 6010 3620 6012
rect 3644 6010 3700 6012
rect 3724 6010 3780 6012
rect 3484 5958 3530 6010
rect 3530 5958 3540 6010
rect 3564 5958 3594 6010
rect 3594 5958 3606 6010
rect 3606 5958 3620 6010
rect 3644 5958 3658 6010
rect 3658 5958 3670 6010
rect 3670 5958 3700 6010
rect 3724 5958 3734 6010
rect 3734 5958 3780 6010
rect 3484 5956 3540 5958
rect 3564 5956 3620 5958
rect 3644 5956 3700 5958
rect 3724 5956 3780 5958
rect 5034 7642 5090 7644
rect 5114 7642 5170 7644
rect 5194 7642 5250 7644
rect 5274 7642 5330 7644
rect 5034 7590 5080 7642
rect 5080 7590 5090 7642
rect 5114 7590 5144 7642
rect 5144 7590 5156 7642
rect 5156 7590 5170 7642
rect 5194 7590 5208 7642
rect 5208 7590 5220 7642
rect 5220 7590 5250 7642
rect 5274 7590 5284 7642
rect 5284 7590 5330 7642
rect 5034 7588 5090 7590
rect 5114 7588 5170 7590
rect 5194 7588 5250 7590
rect 5274 7588 5330 7590
rect 5034 6554 5090 6556
rect 5114 6554 5170 6556
rect 5194 6554 5250 6556
rect 5274 6554 5330 6556
rect 5034 6502 5080 6554
rect 5080 6502 5090 6554
rect 5114 6502 5144 6554
rect 5144 6502 5156 6554
rect 5156 6502 5170 6554
rect 5194 6502 5208 6554
rect 5208 6502 5220 6554
rect 5220 6502 5250 6554
rect 5274 6502 5284 6554
rect 5284 6502 5330 6554
rect 5034 6500 5090 6502
rect 5114 6500 5170 6502
rect 5194 6500 5250 6502
rect 5274 6500 5330 6502
rect 6584 9274 6640 9276
rect 6664 9274 6720 9276
rect 6744 9274 6800 9276
rect 6824 9274 6880 9276
rect 6584 9222 6630 9274
rect 6630 9222 6640 9274
rect 6664 9222 6694 9274
rect 6694 9222 6706 9274
rect 6706 9222 6720 9274
rect 6744 9222 6758 9274
rect 6758 9222 6770 9274
rect 6770 9222 6800 9274
rect 6824 9222 6834 9274
rect 6834 9222 6880 9274
rect 6584 9220 6640 9222
rect 6664 9220 6720 9222
rect 6744 9220 6800 9222
rect 6824 9220 6880 9222
rect 6584 8186 6640 8188
rect 6664 8186 6720 8188
rect 6744 8186 6800 8188
rect 6824 8186 6880 8188
rect 6584 8134 6630 8186
rect 6630 8134 6640 8186
rect 6664 8134 6694 8186
rect 6694 8134 6706 8186
rect 6706 8134 6720 8186
rect 6744 8134 6758 8186
rect 6758 8134 6770 8186
rect 6770 8134 6800 8186
rect 6824 8134 6834 8186
rect 6834 8134 6880 8186
rect 6584 8132 6640 8134
rect 6664 8132 6720 8134
rect 6744 8132 6800 8134
rect 6824 8132 6880 8134
rect 5034 5466 5090 5468
rect 5114 5466 5170 5468
rect 5194 5466 5250 5468
rect 5274 5466 5330 5468
rect 5034 5414 5080 5466
rect 5080 5414 5090 5466
rect 5114 5414 5144 5466
rect 5144 5414 5156 5466
rect 5156 5414 5170 5466
rect 5194 5414 5208 5466
rect 5208 5414 5220 5466
rect 5220 5414 5250 5466
rect 5274 5414 5284 5466
rect 5284 5414 5330 5466
rect 5034 5412 5090 5414
rect 5114 5412 5170 5414
rect 5194 5412 5250 5414
rect 5274 5412 5330 5414
rect 3484 4922 3540 4924
rect 3564 4922 3620 4924
rect 3644 4922 3700 4924
rect 3724 4922 3780 4924
rect 3484 4870 3530 4922
rect 3530 4870 3540 4922
rect 3564 4870 3594 4922
rect 3594 4870 3606 4922
rect 3606 4870 3620 4922
rect 3644 4870 3658 4922
rect 3658 4870 3670 4922
rect 3670 4870 3700 4922
rect 3724 4870 3734 4922
rect 3734 4870 3780 4922
rect 3484 4868 3540 4870
rect 3564 4868 3620 4870
rect 3644 4868 3700 4870
rect 3724 4868 3780 4870
rect 6584 7098 6640 7100
rect 6664 7098 6720 7100
rect 6744 7098 6800 7100
rect 6824 7098 6880 7100
rect 6584 7046 6630 7098
rect 6630 7046 6640 7098
rect 6664 7046 6694 7098
rect 6694 7046 6706 7098
rect 6706 7046 6720 7098
rect 6744 7046 6758 7098
rect 6758 7046 6770 7098
rect 6770 7046 6800 7098
rect 6824 7046 6834 7098
rect 6834 7046 6880 7098
rect 6584 7044 6640 7046
rect 6664 7044 6720 7046
rect 6744 7044 6800 7046
rect 6824 7044 6880 7046
rect 6584 6010 6640 6012
rect 6664 6010 6720 6012
rect 6744 6010 6800 6012
rect 6824 6010 6880 6012
rect 6584 5958 6630 6010
rect 6630 5958 6640 6010
rect 6664 5958 6694 6010
rect 6694 5958 6706 6010
rect 6706 5958 6720 6010
rect 6744 5958 6758 6010
rect 6758 5958 6770 6010
rect 6770 5958 6800 6010
rect 6824 5958 6834 6010
rect 6834 5958 6880 6010
rect 6584 5956 6640 5958
rect 6664 5956 6720 5958
rect 6744 5956 6800 5958
rect 6824 5956 6880 5958
rect 8134 9818 8190 9820
rect 8214 9818 8270 9820
rect 8294 9818 8350 9820
rect 8374 9818 8430 9820
rect 8134 9766 8180 9818
rect 8180 9766 8190 9818
rect 8214 9766 8244 9818
rect 8244 9766 8256 9818
rect 8256 9766 8270 9818
rect 8294 9766 8308 9818
rect 8308 9766 8320 9818
rect 8320 9766 8350 9818
rect 8374 9766 8384 9818
rect 8384 9766 8430 9818
rect 8134 9764 8190 9766
rect 8214 9764 8270 9766
rect 8294 9764 8350 9766
rect 8374 9764 8430 9766
rect 8134 8730 8190 8732
rect 8214 8730 8270 8732
rect 8294 8730 8350 8732
rect 8374 8730 8430 8732
rect 8134 8678 8180 8730
rect 8180 8678 8190 8730
rect 8214 8678 8244 8730
rect 8244 8678 8256 8730
rect 8256 8678 8270 8730
rect 8294 8678 8308 8730
rect 8308 8678 8320 8730
rect 8320 8678 8350 8730
rect 8374 8678 8384 8730
rect 8384 8678 8430 8730
rect 8134 8676 8190 8678
rect 8214 8676 8270 8678
rect 8294 8676 8350 8678
rect 8374 8676 8430 8678
rect 8134 7642 8190 7644
rect 8214 7642 8270 7644
rect 8294 7642 8350 7644
rect 8374 7642 8430 7644
rect 8134 7590 8180 7642
rect 8180 7590 8190 7642
rect 8214 7590 8244 7642
rect 8244 7590 8256 7642
rect 8256 7590 8270 7642
rect 8294 7590 8308 7642
rect 8308 7590 8320 7642
rect 8320 7590 8350 7642
rect 8374 7590 8384 7642
rect 8384 7590 8430 7642
rect 8134 7588 8190 7590
rect 8214 7588 8270 7590
rect 8294 7588 8350 7590
rect 8374 7588 8430 7590
rect 9684 10362 9740 10364
rect 9764 10362 9820 10364
rect 9844 10362 9900 10364
rect 9924 10362 9980 10364
rect 9684 10310 9730 10362
rect 9730 10310 9740 10362
rect 9764 10310 9794 10362
rect 9794 10310 9806 10362
rect 9806 10310 9820 10362
rect 9844 10310 9858 10362
rect 9858 10310 9870 10362
rect 9870 10310 9900 10362
rect 9924 10310 9934 10362
rect 9934 10310 9980 10362
rect 9684 10308 9740 10310
rect 9764 10308 9820 10310
rect 9844 10308 9900 10310
rect 9924 10308 9980 10310
rect 9684 9274 9740 9276
rect 9764 9274 9820 9276
rect 9844 9274 9900 9276
rect 9924 9274 9980 9276
rect 9684 9222 9730 9274
rect 9730 9222 9740 9274
rect 9764 9222 9794 9274
rect 9794 9222 9806 9274
rect 9806 9222 9820 9274
rect 9844 9222 9858 9274
rect 9858 9222 9870 9274
rect 9870 9222 9900 9274
rect 9924 9222 9934 9274
rect 9934 9222 9980 9274
rect 9684 9220 9740 9222
rect 9764 9220 9820 9222
rect 9844 9220 9900 9222
rect 9924 9220 9980 9222
rect 6584 4922 6640 4924
rect 6664 4922 6720 4924
rect 6744 4922 6800 4924
rect 6824 4922 6880 4924
rect 6584 4870 6630 4922
rect 6630 4870 6640 4922
rect 6664 4870 6694 4922
rect 6694 4870 6706 4922
rect 6706 4870 6720 4922
rect 6744 4870 6758 4922
rect 6758 4870 6770 4922
rect 6770 4870 6800 4922
rect 6824 4870 6834 4922
rect 6834 4870 6880 4922
rect 6584 4868 6640 4870
rect 6664 4868 6720 4870
rect 6744 4868 6800 4870
rect 6824 4868 6880 4870
rect 3484 3834 3540 3836
rect 3564 3834 3620 3836
rect 3644 3834 3700 3836
rect 3724 3834 3780 3836
rect 3484 3782 3530 3834
rect 3530 3782 3540 3834
rect 3564 3782 3594 3834
rect 3594 3782 3606 3834
rect 3606 3782 3620 3834
rect 3644 3782 3658 3834
rect 3658 3782 3670 3834
rect 3670 3782 3700 3834
rect 3724 3782 3734 3834
rect 3734 3782 3780 3834
rect 3484 3780 3540 3782
rect 3564 3780 3620 3782
rect 3644 3780 3700 3782
rect 3724 3780 3780 3782
rect 5034 4378 5090 4380
rect 5114 4378 5170 4380
rect 5194 4378 5250 4380
rect 5274 4378 5330 4380
rect 5034 4326 5080 4378
rect 5080 4326 5090 4378
rect 5114 4326 5144 4378
rect 5144 4326 5156 4378
rect 5156 4326 5170 4378
rect 5194 4326 5208 4378
rect 5208 4326 5220 4378
rect 5220 4326 5250 4378
rect 5274 4326 5284 4378
rect 5284 4326 5330 4378
rect 5034 4324 5090 4326
rect 5114 4324 5170 4326
rect 5194 4324 5250 4326
rect 5274 4324 5330 4326
rect 5034 3290 5090 3292
rect 5114 3290 5170 3292
rect 5194 3290 5250 3292
rect 5274 3290 5330 3292
rect 5034 3238 5080 3290
rect 5080 3238 5090 3290
rect 5114 3238 5144 3290
rect 5144 3238 5156 3290
rect 5156 3238 5170 3290
rect 5194 3238 5208 3290
rect 5208 3238 5220 3290
rect 5220 3238 5250 3290
rect 5274 3238 5284 3290
rect 5284 3238 5330 3290
rect 5034 3236 5090 3238
rect 5114 3236 5170 3238
rect 5194 3236 5250 3238
rect 5274 3236 5330 3238
rect 2502 1964 2558 2000
rect 2502 1944 2504 1964
rect 2504 1944 2556 1964
rect 2556 1944 2558 1964
rect 3484 2746 3540 2748
rect 3564 2746 3620 2748
rect 3644 2746 3700 2748
rect 3724 2746 3780 2748
rect 3484 2694 3530 2746
rect 3530 2694 3540 2746
rect 3564 2694 3594 2746
rect 3594 2694 3606 2746
rect 3606 2694 3620 2746
rect 3644 2694 3658 2746
rect 3658 2694 3670 2746
rect 3670 2694 3700 2746
rect 3724 2694 3734 2746
rect 3734 2694 3780 2746
rect 3484 2692 3540 2694
rect 3564 2692 3620 2694
rect 3644 2692 3700 2694
rect 3724 2692 3780 2694
rect 4710 1944 4766 2000
rect 5034 2202 5090 2204
rect 5114 2202 5170 2204
rect 5194 2202 5250 2204
rect 5274 2202 5330 2204
rect 5034 2150 5080 2202
rect 5080 2150 5090 2202
rect 5114 2150 5144 2202
rect 5144 2150 5156 2202
rect 5156 2150 5170 2202
rect 5194 2150 5208 2202
rect 5208 2150 5220 2202
rect 5220 2150 5250 2202
rect 5274 2150 5284 2202
rect 5284 2150 5330 2202
rect 5034 2148 5090 2150
rect 5114 2148 5170 2150
rect 5194 2148 5250 2150
rect 5274 2148 5330 2150
rect 3484 1658 3540 1660
rect 3564 1658 3620 1660
rect 3644 1658 3700 1660
rect 3724 1658 3780 1660
rect 3484 1606 3530 1658
rect 3530 1606 3540 1658
rect 3564 1606 3594 1658
rect 3594 1606 3606 1658
rect 3606 1606 3620 1658
rect 3644 1606 3658 1658
rect 3658 1606 3670 1658
rect 3670 1606 3700 1658
rect 3724 1606 3734 1658
rect 3734 1606 3780 1658
rect 3484 1604 3540 1606
rect 3564 1604 3620 1606
rect 3644 1604 3700 1606
rect 3724 1604 3780 1606
rect 3974 892 3976 912
rect 3976 892 4028 912
rect 4028 892 4030 912
rect 3974 856 4030 892
rect 3484 570 3540 572
rect 3564 570 3620 572
rect 3644 570 3700 572
rect 3724 570 3780 572
rect 3484 518 3530 570
rect 3530 518 3540 570
rect 3564 518 3594 570
rect 3594 518 3606 570
rect 3606 518 3620 570
rect 3644 518 3658 570
rect 3658 518 3670 570
rect 3670 518 3700 570
rect 3724 518 3734 570
rect 3734 518 3780 570
rect 3484 516 3540 518
rect 3564 516 3620 518
rect 3644 516 3700 518
rect 3724 516 3780 518
rect 6584 3834 6640 3836
rect 6664 3834 6720 3836
rect 6744 3834 6800 3836
rect 6824 3834 6880 3836
rect 6584 3782 6630 3834
rect 6630 3782 6640 3834
rect 6664 3782 6694 3834
rect 6694 3782 6706 3834
rect 6706 3782 6720 3834
rect 6744 3782 6758 3834
rect 6758 3782 6770 3834
rect 6770 3782 6800 3834
rect 6824 3782 6834 3834
rect 6834 3782 6880 3834
rect 6584 3780 6640 3782
rect 6664 3780 6720 3782
rect 6744 3780 6800 3782
rect 6824 3780 6880 3782
rect 9684 8186 9740 8188
rect 9764 8186 9820 8188
rect 9844 8186 9900 8188
rect 9924 8186 9980 8188
rect 9684 8134 9730 8186
rect 9730 8134 9740 8186
rect 9764 8134 9794 8186
rect 9794 8134 9806 8186
rect 9806 8134 9820 8186
rect 9844 8134 9858 8186
rect 9858 8134 9870 8186
rect 9870 8134 9900 8186
rect 9924 8134 9934 8186
rect 9934 8134 9980 8186
rect 9684 8132 9740 8134
rect 9764 8132 9820 8134
rect 9844 8132 9900 8134
rect 9924 8132 9980 8134
rect 8134 6554 8190 6556
rect 8214 6554 8270 6556
rect 8294 6554 8350 6556
rect 8374 6554 8430 6556
rect 8134 6502 8180 6554
rect 8180 6502 8190 6554
rect 8214 6502 8244 6554
rect 8244 6502 8256 6554
rect 8256 6502 8270 6554
rect 8294 6502 8308 6554
rect 8308 6502 8320 6554
rect 8320 6502 8350 6554
rect 8374 6502 8384 6554
rect 8384 6502 8430 6554
rect 8134 6500 8190 6502
rect 8214 6500 8270 6502
rect 8294 6500 8350 6502
rect 8374 6500 8430 6502
rect 8134 5466 8190 5468
rect 8214 5466 8270 5468
rect 8294 5466 8350 5468
rect 8374 5466 8430 5468
rect 8134 5414 8180 5466
rect 8180 5414 8190 5466
rect 8214 5414 8244 5466
rect 8244 5414 8256 5466
rect 8256 5414 8270 5466
rect 8294 5414 8308 5466
rect 8308 5414 8320 5466
rect 8320 5414 8350 5466
rect 8374 5414 8384 5466
rect 8384 5414 8430 5466
rect 8134 5412 8190 5414
rect 8214 5412 8270 5414
rect 8294 5412 8350 5414
rect 8374 5412 8430 5414
rect 10046 7404 10102 7440
rect 10046 7384 10048 7404
rect 10048 7384 10100 7404
rect 10100 7384 10102 7404
rect 9684 7098 9740 7100
rect 9764 7098 9820 7100
rect 9844 7098 9900 7100
rect 9924 7098 9980 7100
rect 9684 7046 9730 7098
rect 9730 7046 9740 7098
rect 9764 7046 9794 7098
rect 9794 7046 9806 7098
rect 9806 7046 9820 7098
rect 9844 7046 9858 7098
rect 9858 7046 9870 7098
rect 9870 7046 9900 7098
rect 9924 7046 9934 7098
rect 9934 7046 9980 7098
rect 9684 7044 9740 7046
rect 9764 7044 9820 7046
rect 9844 7044 9900 7046
rect 9924 7044 9980 7046
rect 9684 6010 9740 6012
rect 9764 6010 9820 6012
rect 9844 6010 9900 6012
rect 9924 6010 9980 6012
rect 9684 5958 9730 6010
rect 9730 5958 9740 6010
rect 9764 5958 9794 6010
rect 9794 5958 9806 6010
rect 9806 5958 9820 6010
rect 9844 5958 9858 6010
rect 9858 5958 9870 6010
rect 9870 5958 9900 6010
rect 9924 5958 9934 6010
rect 9934 5958 9980 6010
rect 9684 5956 9740 5958
rect 9764 5956 9820 5958
rect 9844 5956 9900 5958
rect 9924 5956 9980 5958
rect 10230 6840 10286 6896
rect 11234 9818 11290 9820
rect 11314 9818 11370 9820
rect 11394 9818 11450 9820
rect 11474 9818 11530 9820
rect 11234 9766 11280 9818
rect 11280 9766 11290 9818
rect 11314 9766 11344 9818
rect 11344 9766 11356 9818
rect 11356 9766 11370 9818
rect 11394 9766 11408 9818
rect 11408 9766 11420 9818
rect 11420 9766 11450 9818
rect 11474 9766 11484 9818
rect 11484 9766 11530 9818
rect 11234 9764 11290 9766
rect 11314 9764 11370 9766
rect 11394 9764 11450 9766
rect 11474 9764 11530 9766
rect 12784 10362 12840 10364
rect 12864 10362 12920 10364
rect 12944 10362 13000 10364
rect 13024 10362 13080 10364
rect 12784 10310 12830 10362
rect 12830 10310 12840 10362
rect 12864 10310 12894 10362
rect 12894 10310 12906 10362
rect 12906 10310 12920 10362
rect 12944 10310 12958 10362
rect 12958 10310 12970 10362
rect 12970 10310 13000 10362
rect 13024 10310 13034 10362
rect 13034 10310 13080 10362
rect 12784 10308 12840 10310
rect 12864 10308 12920 10310
rect 12944 10308 13000 10310
rect 13024 10308 13080 10310
rect 12784 9274 12840 9276
rect 12864 9274 12920 9276
rect 12944 9274 13000 9276
rect 13024 9274 13080 9276
rect 12784 9222 12830 9274
rect 12830 9222 12840 9274
rect 12864 9222 12894 9274
rect 12894 9222 12906 9274
rect 12906 9222 12920 9274
rect 12944 9222 12958 9274
rect 12958 9222 12970 9274
rect 12970 9222 13000 9274
rect 13024 9222 13034 9274
rect 13034 9222 13080 9274
rect 12784 9220 12840 9222
rect 12864 9220 12920 9222
rect 12944 9220 13000 9222
rect 13024 9220 13080 9222
rect 11234 8730 11290 8732
rect 11314 8730 11370 8732
rect 11394 8730 11450 8732
rect 11474 8730 11530 8732
rect 11234 8678 11280 8730
rect 11280 8678 11290 8730
rect 11314 8678 11344 8730
rect 11344 8678 11356 8730
rect 11356 8678 11370 8730
rect 11394 8678 11408 8730
rect 11408 8678 11420 8730
rect 11420 8678 11450 8730
rect 11474 8678 11484 8730
rect 11484 8678 11530 8730
rect 11234 8676 11290 8678
rect 11314 8676 11370 8678
rect 11394 8676 11450 8678
rect 11474 8676 11530 8678
rect 10414 7420 10416 7440
rect 10416 7420 10468 7440
rect 10468 7420 10470 7440
rect 10414 7384 10470 7420
rect 10598 7404 10654 7440
rect 10598 7384 10600 7404
rect 10600 7384 10652 7404
rect 10652 7384 10654 7404
rect 10414 7248 10470 7304
rect 10690 6876 10692 6896
rect 10692 6876 10744 6896
rect 10744 6876 10746 6896
rect 10690 6840 10746 6876
rect 11334 7928 11390 7984
rect 10414 6724 10470 6760
rect 11058 6740 11060 6760
rect 11060 6740 11112 6760
rect 11112 6740 11114 6760
rect 10414 6704 10416 6724
rect 10416 6704 10468 6724
rect 10468 6704 10470 6724
rect 11058 6704 11114 6740
rect 11234 7642 11290 7644
rect 11314 7642 11370 7644
rect 11394 7642 11450 7644
rect 11474 7642 11530 7644
rect 11234 7590 11280 7642
rect 11280 7590 11290 7642
rect 11314 7590 11344 7642
rect 11344 7590 11356 7642
rect 11356 7590 11370 7642
rect 11394 7590 11408 7642
rect 11408 7590 11420 7642
rect 11420 7590 11450 7642
rect 11474 7590 11484 7642
rect 11484 7590 11530 7642
rect 11234 7588 11290 7590
rect 11314 7588 11370 7590
rect 11394 7588 11450 7590
rect 11474 7588 11530 7590
rect 11234 6554 11290 6556
rect 11314 6554 11370 6556
rect 11394 6554 11450 6556
rect 11474 6554 11530 6556
rect 11234 6502 11280 6554
rect 11280 6502 11290 6554
rect 11314 6502 11344 6554
rect 11344 6502 11356 6554
rect 11356 6502 11370 6554
rect 11394 6502 11408 6554
rect 11408 6502 11420 6554
rect 11420 6502 11450 6554
rect 11474 6502 11484 6554
rect 11484 6502 11530 6554
rect 11234 6500 11290 6502
rect 11314 6500 11370 6502
rect 11394 6500 11450 6502
rect 11474 6500 11530 6502
rect 12784 8186 12840 8188
rect 12864 8186 12920 8188
rect 12944 8186 13000 8188
rect 13024 8186 13080 8188
rect 12784 8134 12830 8186
rect 12830 8134 12840 8186
rect 12864 8134 12894 8186
rect 12894 8134 12906 8186
rect 12906 8134 12920 8186
rect 12944 8134 12958 8186
rect 12958 8134 12970 8186
rect 12970 8134 13000 8186
rect 13024 8134 13034 8186
rect 13034 8134 13080 8186
rect 12784 8132 12840 8134
rect 12864 8132 12920 8134
rect 12944 8132 13000 8134
rect 13024 8132 13080 8134
rect 12714 7284 12716 7304
rect 12716 7284 12768 7304
rect 12768 7284 12770 7304
rect 12714 7248 12770 7284
rect 12784 7098 12840 7100
rect 12864 7098 12920 7100
rect 12944 7098 13000 7100
rect 13024 7098 13080 7100
rect 12784 7046 12830 7098
rect 12830 7046 12840 7098
rect 12864 7046 12894 7098
rect 12894 7046 12906 7098
rect 12906 7046 12920 7098
rect 12944 7046 12958 7098
rect 12958 7046 12970 7098
rect 12970 7046 13000 7098
rect 13024 7046 13034 7098
rect 13034 7046 13080 7098
rect 12784 7044 12840 7046
rect 12864 7044 12920 7046
rect 12944 7044 13000 7046
rect 13024 7044 13080 7046
rect 12784 6010 12840 6012
rect 12864 6010 12920 6012
rect 12944 6010 13000 6012
rect 13024 6010 13080 6012
rect 12784 5958 12830 6010
rect 12830 5958 12840 6010
rect 12864 5958 12894 6010
rect 12894 5958 12906 6010
rect 12906 5958 12920 6010
rect 12944 5958 12958 6010
rect 12958 5958 12970 6010
rect 12970 5958 13000 6010
rect 13024 5958 13034 6010
rect 13034 5958 13080 6010
rect 12784 5956 12840 5958
rect 12864 5956 12920 5958
rect 12944 5956 13000 5958
rect 13024 5956 13080 5958
rect 11234 5466 11290 5468
rect 11314 5466 11370 5468
rect 11394 5466 11450 5468
rect 11474 5466 11530 5468
rect 11234 5414 11280 5466
rect 11280 5414 11290 5466
rect 11314 5414 11344 5466
rect 11344 5414 11356 5466
rect 11356 5414 11370 5466
rect 11394 5414 11408 5466
rect 11408 5414 11420 5466
rect 11420 5414 11450 5466
rect 11474 5414 11484 5466
rect 11484 5414 11530 5466
rect 11234 5412 11290 5414
rect 11314 5412 11370 5414
rect 11394 5412 11450 5414
rect 11474 5412 11530 5414
rect 9684 4922 9740 4924
rect 9764 4922 9820 4924
rect 9844 4922 9900 4924
rect 9924 4922 9980 4924
rect 9684 4870 9730 4922
rect 9730 4870 9740 4922
rect 9764 4870 9794 4922
rect 9794 4870 9806 4922
rect 9806 4870 9820 4922
rect 9844 4870 9858 4922
rect 9858 4870 9870 4922
rect 9870 4870 9900 4922
rect 9924 4870 9934 4922
rect 9934 4870 9980 4922
rect 9684 4868 9740 4870
rect 9764 4868 9820 4870
rect 9844 4868 9900 4870
rect 9924 4868 9980 4870
rect 8134 4378 8190 4380
rect 8214 4378 8270 4380
rect 8294 4378 8350 4380
rect 8374 4378 8430 4380
rect 8134 4326 8180 4378
rect 8180 4326 8190 4378
rect 8214 4326 8244 4378
rect 8244 4326 8256 4378
rect 8256 4326 8270 4378
rect 8294 4326 8308 4378
rect 8308 4326 8320 4378
rect 8320 4326 8350 4378
rect 8374 4326 8384 4378
rect 8384 4326 8430 4378
rect 8134 4324 8190 4326
rect 8214 4324 8270 4326
rect 8294 4324 8350 4326
rect 8374 4324 8430 4326
rect 12784 4922 12840 4924
rect 12864 4922 12920 4924
rect 12944 4922 13000 4924
rect 13024 4922 13080 4924
rect 12784 4870 12830 4922
rect 12830 4870 12840 4922
rect 12864 4870 12894 4922
rect 12894 4870 12906 4922
rect 12906 4870 12920 4922
rect 12944 4870 12958 4922
rect 12958 4870 12970 4922
rect 12970 4870 13000 4922
rect 13024 4870 13034 4922
rect 13034 4870 13080 4922
rect 12784 4868 12840 4870
rect 12864 4868 12920 4870
rect 12944 4868 13000 4870
rect 13024 4868 13080 4870
rect 14334 9818 14390 9820
rect 14414 9818 14470 9820
rect 14494 9818 14550 9820
rect 14574 9818 14630 9820
rect 14334 9766 14380 9818
rect 14380 9766 14390 9818
rect 14414 9766 14444 9818
rect 14444 9766 14456 9818
rect 14456 9766 14470 9818
rect 14494 9766 14508 9818
rect 14508 9766 14520 9818
rect 14520 9766 14550 9818
rect 14574 9766 14584 9818
rect 14584 9766 14630 9818
rect 14334 9764 14390 9766
rect 14414 9764 14470 9766
rect 14494 9764 14550 9766
rect 14574 9764 14630 9766
rect 14334 8730 14390 8732
rect 14414 8730 14470 8732
rect 14494 8730 14550 8732
rect 14574 8730 14630 8732
rect 14334 8678 14380 8730
rect 14380 8678 14390 8730
rect 14414 8678 14444 8730
rect 14444 8678 14456 8730
rect 14456 8678 14470 8730
rect 14494 8678 14508 8730
rect 14508 8678 14520 8730
rect 14520 8678 14550 8730
rect 14574 8678 14584 8730
rect 14584 8678 14630 8730
rect 14334 8676 14390 8678
rect 14414 8676 14470 8678
rect 14494 8676 14550 8678
rect 14574 8676 14630 8678
rect 14334 7642 14390 7644
rect 14414 7642 14470 7644
rect 14494 7642 14550 7644
rect 14574 7642 14630 7644
rect 14334 7590 14380 7642
rect 14380 7590 14390 7642
rect 14414 7590 14444 7642
rect 14444 7590 14456 7642
rect 14456 7590 14470 7642
rect 14494 7590 14508 7642
rect 14508 7590 14520 7642
rect 14520 7590 14550 7642
rect 14574 7590 14584 7642
rect 14584 7590 14630 7642
rect 14334 7588 14390 7590
rect 14414 7588 14470 7590
rect 14494 7588 14550 7590
rect 14574 7588 14630 7590
rect 14002 7384 14058 7440
rect 14334 6554 14390 6556
rect 14414 6554 14470 6556
rect 14494 6554 14550 6556
rect 14574 6554 14630 6556
rect 14334 6502 14380 6554
rect 14380 6502 14390 6554
rect 14414 6502 14444 6554
rect 14444 6502 14456 6554
rect 14456 6502 14470 6554
rect 14494 6502 14508 6554
rect 14508 6502 14520 6554
rect 14520 6502 14550 6554
rect 14574 6502 14584 6554
rect 14584 6502 14630 6554
rect 14334 6500 14390 6502
rect 14414 6500 14470 6502
rect 14494 6500 14550 6502
rect 14574 6500 14630 6502
rect 15106 7928 15162 7984
rect 17434 10906 17490 10908
rect 17514 10906 17570 10908
rect 17594 10906 17650 10908
rect 17674 10906 17730 10908
rect 17434 10854 17480 10906
rect 17480 10854 17490 10906
rect 17514 10854 17544 10906
rect 17544 10854 17556 10906
rect 17556 10854 17570 10906
rect 17594 10854 17608 10906
rect 17608 10854 17620 10906
rect 17620 10854 17650 10906
rect 17674 10854 17684 10906
rect 17684 10854 17730 10906
rect 17434 10852 17490 10854
rect 17514 10852 17570 10854
rect 17594 10852 17650 10854
rect 17674 10852 17730 10854
rect 15884 10362 15940 10364
rect 15964 10362 16020 10364
rect 16044 10362 16100 10364
rect 16124 10362 16180 10364
rect 15884 10310 15930 10362
rect 15930 10310 15940 10362
rect 15964 10310 15994 10362
rect 15994 10310 16006 10362
rect 16006 10310 16020 10362
rect 16044 10310 16058 10362
rect 16058 10310 16070 10362
rect 16070 10310 16100 10362
rect 16124 10310 16134 10362
rect 16134 10310 16180 10362
rect 15884 10308 15940 10310
rect 15964 10308 16020 10310
rect 16044 10308 16100 10310
rect 16124 10308 16180 10310
rect 17434 9818 17490 9820
rect 17514 9818 17570 9820
rect 17594 9818 17650 9820
rect 17674 9818 17730 9820
rect 17434 9766 17480 9818
rect 17480 9766 17490 9818
rect 17514 9766 17544 9818
rect 17544 9766 17556 9818
rect 17556 9766 17570 9818
rect 17594 9766 17608 9818
rect 17608 9766 17620 9818
rect 17620 9766 17650 9818
rect 17674 9766 17684 9818
rect 17684 9766 17730 9818
rect 17434 9764 17490 9766
rect 17514 9764 17570 9766
rect 17594 9764 17650 9766
rect 17674 9764 17730 9766
rect 15884 9274 15940 9276
rect 15964 9274 16020 9276
rect 16044 9274 16100 9276
rect 16124 9274 16180 9276
rect 15884 9222 15930 9274
rect 15930 9222 15940 9274
rect 15964 9222 15994 9274
rect 15994 9222 16006 9274
rect 16006 9222 16020 9274
rect 16044 9222 16058 9274
rect 16058 9222 16070 9274
rect 16070 9222 16100 9274
rect 16124 9222 16134 9274
rect 16134 9222 16180 9274
rect 15884 9220 15940 9222
rect 15964 9220 16020 9222
rect 16044 9220 16100 9222
rect 16124 9220 16180 9222
rect 17434 8730 17490 8732
rect 17514 8730 17570 8732
rect 17594 8730 17650 8732
rect 17674 8730 17730 8732
rect 17434 8678 17480 8730
rect 17480 8678 17490 8730
rect 17514 8678 17544 8730
rect 17544 8678 17556 8730
rect 17556 8678 17570 8730
rect 17594 8678 17608 8730
rect 17608 8678 17620 8730
rect 17620 8678 17650 8730
rect 17674 8678 17684 8730
rect 17684 8678 17730 8730
rect 17434 8676 17490 8678
rect 17514 8676 17570 8678
rect 17594 8676 17650 8678
rect 17674 8676 17730 8678
rect 15884 8186 15940 8188
rect 15964 8186 16020 8188
rect 16044 8186 16100 8188
rect 16124 8186 16180 8188
rect 15884 8134 15930 8186
rect 15930 8134 15940 8186
rect 15964 8134 15994 8186
rect 15994 8134 16006 8186
rect 16006 8134 16020 8186
rect 16044 8134 16058 8186
rect 16058 8134 16070 8186
rect 16070 8134 16100 8186
rect 16124 8134 16134 8186
rect 16134 8134 16180 8186
rect 15884 8132 15940 8134
rect 15964 8132 16020 8134
rect 16044 8132 16100 8134
rect 16124 8132 16180 8134
rect 15884 7098 15940 7100
rect 15964 7098 16020 7100
rect 16044 7098 16100 7100
rect 16124 7098 16180 7100
rect 15884 7046 15930 7098
rect 15930 7046 15940 7098
rect 15964 7046 15994 7098
rect 15994 7046 16006 7098
rect 16006 7046 16020 7098
rect 16044 7046 16058 7098
rect 16058 7046 16070 7098
rect 16070 7046 16100 7098
rect 16124 7046 16134 7098
rect 16134 7046 16180 7098
rect 15884 7044 15940 7046
rect 15964 7044 16020 7046
rect 16044 7044 16100 7046
rect 16124 7044 16180 7046
rect 18786 11192 18842 11248
rect 18694 9696 18750 9752
rect 18602 8200 18658 8256
rect 14334 5466 14390 5468
rect 14414 5466 14470 5468
rect 14494 5466 14550 5468
rect 14574 5466 14630 5468
rect 14334 5414 14380 5466
rect 14380 5414 14390 5466
rect 14414 5414 14444 5466
rect 14444 5414 14456 5466
rect 14456 5414 14470 5466
rect 14494 5414 14508 5466
rect 14508 5414 14520 5466
rect 14520 5414 14550 5466
rect 14574 5414 14584 5466
rect 14584 5414 14630 5466
rect 14334 5412 14390 5414
rect 14414 5412 14470 5414
rect 14494 5412 14550 5414
rect 14574 5412 14630 5414
rect 15884 6010 15940 6012
rect 15964 6010 16020 6012
rect 16044 6010 16100 6012
rect 16124 6010 16180 6012
rect 15884 5958 15930 6010
rect 15930 5958 15940 6010
rect 15964 5958 15994 6010
rect 15994 5958 16006 6010
rect 16006 5958 16020 6010
rect 16044 5958 16058 6010
rect 16058 5958 16070 6010
rect 16070 5958 16100 6010
rect 16124 5958 16134 6010
rect 16134 5958 16180 6010
rect 15884 5956 15940 5958
rect 15964 5956 16020 5958
rect 16044 5956 16100 5958
rect 16124 5956 16180 5958
rect 11234 4378 11290 4380
rect 11314 4378 11370 4380
rect 11394 4378 11450 4380
rect 11474 4378 11530 4380
rect 11234 4326 11280 4378
rect 11280 4326 11290 4378
rect 11314 4326 11344 4378
rect 11344 4326 11356 4378
rect 11356 4326 11370 4378
rect 11394 4326 11408 4378
rect 11408 4326 11420 4378
rect 11420 4326 11450 4378
rect 11474 4326 11484 4378
rect 11484 4326 11530 4378
rect 11234 4324 11290 4326
rect 11314 4324 11370 4326
rect 11394 4324 11450 4326
rect 11474 4324 11530 4326
rect 8134 3290 8190 3292
rect 8214 3290 8270 3292
rect 8294 3290 8350 3292
rect 8374 3290 8430 3292
rect 8134 3238 8180 3290
rect 8180 3238 8190 3290
rect 8214 3238 8244 3290
rect 8244 3238 8256 3290
rect 8256 3238 8270 3290
rect 8294 3238 8308 3290
rect 8308 3238 8320 3290
rect 8320 3238 8350 3290
rect 8374 3238 8384 3290
rect 8384 3238 8430 3290
rect 8134 3236 8190 3238
rect 8214 3236 8270 3238
rect 8294 3236 8350 3238
rect 8374 3236 8430 3238
rect 6584 2746 6640 2748
rect 6664 2746 6720 2748
rect 6744 2746 6800 2748
rect 6824 2746 6880 2748
rect 6584 2694 6630 2746
rect 6630 2694 6640 2746
rect 6664 2694 6694 2746
rect 6694 2694 6706 2746
rect 6706 2694 6720 2746
rect 6744 2694 6758 2746
rect 6758 2694 6770 2746
rect 6770 2694 6800 2746
rect 6824 2694 6834 2746
rect 6834 2694 6880 2746
rect 6584 2692 6640 2694
rect 6664 2692 6720 2694
rect 6744 2692 6800 2694
rect 6824 2692 6880 2694
rect 5034 1114 5090 1116
rect 5114 1114 5170 1116
rect 5194 1114 5250 1116
rect 5274 1114 5330 1116
rect 5034 1062 5080 1114
rect 5080 1062 5090 1114
rect 5114 1062 5144 1114
rect 5144 1062 5156 1114
rect 5156 1062 5170 1114
rect 5194 1062 5208 1114
rect 5208 1062 5220 1114
rect 5220 1062 5250 1114
rect 5274 1062 5284 1114
rect 5284 1062 5330 1114
rect 5034 1060 5090 1062
rect 5114 1060 5170 1062
rect 5194 1060 5250 1062
rect 5274 1060 5330 1062
rect 5906 892 5908 912
rect 5908 892 5960 912
rect 5960 892 5962 912
rect 5906 856 5962 892
rect 5078 312 5134 368
rect 6584 1658 6640 1660
rect 6664 1658 6720 1660
rect 6744 1658 6800 1660
rect 6824 1658 6880 1660
rect 6584 1606 6630 1658
rect 6630 1606 6640 1658
rect 6664 1606 6694 1658
rect 6694 1606 6706 1658
rect 6706 1606 6720 1658
rect 6744 1606 6758 1658
rect 6758 1606 6770 1658
rect 6770 1606 6800 1658
rect 6824 1606 6834 1658
rect 6834 1606 6880 1658
rect 6584 1604 6640 1606
rect 6664 1604 6720 1606
rect 6744 1604 6800 1606
rect 6824 1604 6880 1606
rect 8134 2202 8190 2204
rect 8214 2202 8270 2204
rect 8294 2202 8350 2204
rect 8374 2202 8430 2204
rect 8134 2150 8180 2202
rect 8180 2150 8190 2202
rect 8214 2150 8244 2202
rect 8244 2150 8256 2202
rect 8256 2150 8270 2202
rect 8294 2150 8308 2202
rect 8308 2150 8320 2202
rect 8320 2150 8350 2202
rect 8374 2150 8384 2202
rect 8384 2150 8430 2202
rect 8134 2148 8190 2150
rect 8214 2148 8270 2150
rect 8294 2148 8350 2150
rect 8374 2148 8430 2150
rect 9684 3834 9740 3836
rect 9764 3834 9820 3836
rect 9844 3834 9900 3836
rect 9924 3834 9980 3836
rect 9684 3782 9730 3834
rect 9730 3782 9740 3834
rect 9764 3782 9794 3834
rect 9794 3782 9806 3834
rect 9806 3782 9820 3834
rect 9844 3782 9858 3834
rect 9858 3782 9870 3834
rect 9870 3782 9900 3834
rect 9924 3782 9934 3834
rect 9934 3782 9980 3834
rect 9684 3780 9740 3782
rect 9764 3780 9820 3782
rect 9844 3780 9900 3782
rect 9924 3780 9980 3782
rect 9684 2746 9740 2748
rect 9764 2746 9820 2748
rect 9844 2746 9900 2748
rect 9924 2746 9980 2748
rect 9684 2694 9730 2746
rect 9730 2694 9740 2746
rect 9764 2694 9794 2746
rect 9794 2694 9806 2746
rect 9806 2694 9820 2746
rect 9844 2694 9858 2746
rect 9858 2694 9870 2746
rect 9870 2694 9900 2746
rect 9924 2694 9934 2746
rect 9934 2694 9980 2746
rect 9684 2692 9740 2694
rect 9764 2692 9820 2694
rect 9844 2692 9900 2694
rect 9924 2692 9980 2694
rect 8206 1300 8208 1320
rect 8208 1300 8260 1320
rect 8260 1300 8262 1320
rect 6584 570 6640 572
rect 6664 570 6720 572
rect 6744 570 6800 572
rect 6824 570 6880 572
rect 6584 518 6630 570
rect 6630 518 6640 570
rect 6664 518 6694 570
rect 6694 518 6706 570
rect 6706 518 6720 570
rect 6744 518 6758 570
rect 6758 518 6770 570
rect 6770 518 6800 570
rect 6824 518 6834 570
rect 6834 518 6880 570
rect 6584 516 6640 518
rect 6664 516 6720 518
rect 6744 516 6800 518
rect 6824 516 6880 518
rect 8206 1264 8262 1300
rect 8134 1114 8190 1116
rect 8214 1114 8270 1116
rect 8294 1114 8350 1116
rect 8374 1114 8430 1116
rect 8134 1062 8180 1114
rect 8180 1062 8190 1114
rect 8214 1062 8244 1114
rect 8244 1062 8256 1114
rect 8256 1062 8270 1114
rect 8294 1062 8308 1114
rect 8308 1062 8320 1114
rect 8320 1062 8350 1114
rect 8374 1062 8384 1114
rect 8384 1062 8430 1114
rect 8134 1060 8190 1062
rect 8214 1060 8270 1062
rect 8294 1060 8350 1062
rect 8374 1060 8430 1062
rect 9684 1658 9740 1660
rect 9764 1658 9820 1660
rect 9844 1658 9900 1660
rect 9924 1658 9980 1660
rect 9684 1606 9730 1658
rect 9730 1606 9740 1658
rect 9764 1606 9794 1658
rect 9794 1606 9806 1658
rect 9806 1606 9820 1658
rect 9844 1606 9858 1658
rect 9858 1606 9870 1658
rect 9870 1606 9900 1658
rect 9924 1606 9934 1658
rect 9934 1606 9980 1658
rect 9684 1604 9740 1606
rect 9764 1604 9820 1606
rect 9844 1604 9900 1606
rect 9924 1604 9980 1606
rect 11234 3290 11290 3292
rect 11314 3290 11370 3292
rect 11394 3290 11450 3292
rect 11474 3290 11530 3292
rect 11234 3238 11280 3290
rect 11280 3238 11290 3290
rect 11314 3238 11344 3290
rect 11344 3238 11356 3290
rect 11356 3238 11370 3290
rect 11394 3238 11408 3290
rect 11408 3238 11420 3290
rect 11420 3238 11450 3290
rect 11474 3238 11484 3290
rect 11484 3238 11530 3290
rect 11234 3236 11290 3238
rect 11314 3236 11370 3238
rect 11394 3236 11450 3238
rect 11474 3236 11530 3238
rect 11234 2202 11290 2204
rect 11314 2202 11370 2204
rect 11394 2202 11450 2204
rect 11474 2202 11530 2204
rect 11234 2150 11280 2202
rect 11280 2150 11290 2202
rect 11314 2150 11344 2202
rect 11344 2150 11356 2202
rect 11356 2150 11370 2202
rect 11394 2150 11408 2202
rect 11408 2150 11420 2202
rect 11420 2150 11450 2202
rect 11474 2150 11484 2202
rect 11484 2150 11530 2202
rect 11234 2148 11290 2150
rect 11314 2148 11370 2150
rect 11394 2148 11450 2150
rect 11474 2148 11530 2150
rect 10598 856 10654 912
rect 10966 1264 11022 1320
rect 12784 3834 12840 3836
rect 12864 3834 12920 3836
rect 12944 3834 13000 3836
rect 13024 3834 13080 3836
rect 12784 3782 12830 3834
rect 12830 3782 12840 3834
rect 12864 3782 12894 3834
rect 12894 3782 12906 3834
rect 12906 3782 12920 3834
rect 12944 3782 12958 3834
rect 12958 3782 12970 3834
rect 12970 3782 13000 3834
rect 13024 3782 13034 3834
rect 13034 3782 13080 3834
rect 12784 3780 12840 3782
rect 12864 3780 12920 3782
rect 12944 3780 13000 3782
rect 13024 3780 13080 3782
rect 12784 2746 12840 2748
rect 12864 2746 12920 2748
rect 12944 2746 13000 2748
rect 13024 2746 13080 2748
rect 12784 2694 12830 2746
rect 12830 2694 12840 2746
rect 12864 2694 12894 2746
rect 12894 2694 12906 2746
rect 12906 2694 12920 2746
rect 12944 2694 12958 2746
rect 12958 2694 12970 2746
rect 12970 2694 13000 2746
rect 13024 2694 13034 2746
rect 13034 2694 13080 2746
rect 12784 2692 12840 2694
rect 12864 2692 12920 2694
rect 12944 2692 13000 2694
rect 13024 2692 13080 2694
rect 12784 1658 12840 1660
rect 12864 1658 12920 1660
rect 12944 1658 13000 1660
rect 13024 1658 13080 1660
rect 12784 1606 12830 1658
rect 12830 1606 12840 1658
rect 12864 1606 12894 1658
rect 12894 1606 12906 1658
rect 12906 1606 12920 1658
rect 12944 1606 12958 1658
rect 12958 1606 12970 1658
rect 12970 1606 13000 1658
rect 13024 1606 13034 1658
rect 13034 1606 13080 1658
rect 12784 1604 12840 1606
rect 12864 1604 12920 1606
rect 12944 1604 13000 1606
rect 13024 1604 13080 1606
rect 17434 7642 17490 7644
rect 17514 7642 17570 7644
rect 17594 7642 17650 7644
rect 17674 7642 17730 7644
rect 17434 7590 17480 7642
rect 17480 7590 17490 7642
rect 17514 7590 17544 7642
rect 17544 7590 17556 7642
rect 17556 7590 17570 7642
rect 17594 7590 17608 7642
rect 17608 7590 17620 7642
rect 17620 7590 17650 7642
rect 17674 7590 17684 7642
rect 17684 7590 17730 7642
rect 17434 7588 17490 7590
rect 17514 7588 17570 7590
rect 17594 7588 17650 7590
rect 17674 7588 17730 7590
rect 17434 6554 17490 6556
rect 17514 6554 17570 6556
rect 17594 6554 17650 6556
rect 17674 6554 17730 6556
rect 17434 6502 17480 6554
rect 17480 6502 17490 6554
rect 17514 6502 17544 6554
rect 17544 6502 17556 6554
rect 17556 6502 17570 6554
rect 17594 6502 17608 6554
rect 17608 6502 17620 6554
rect 17620 6502 17650 6554
rect 17674 6502 17684 6554
rect 17684 6502 17730 6554
rect 17434 6500 17490 6502
rect 17514 6500 17570 6502
rect 17594 6500 17650 6502
rect 17674 6500 17730 6502
rect 18510 6704 18566 6760
rect 15884 4922 15940 4924
rect 15964 4922 16020 4924
rect 16044 4922 16100 4924
rect 16124 4922 16180 4924
rect 15884 4870 15930 4922
rect 15930 4870 15940 4922
rect 15964 4870 15994 4922
rect 15994 4870 16006 4922
rect 16006 4870 16020 4922
rect 16044 4870 16058 4922
rect 16058 4870 16070 4922
rect 16070 4870 16100 4922
rect 16124 4870 16134 4922
rect 16134 4870 16180 4922
rect 15884 4868 15940 4870
rect 15964 4868 16020 4870
rect 16044 4868 16100 4870
rect 16124 4868 16180 4870
rect 17434 5466 17490 5468
rect 17514 5466 17570 5468
rect 17594 5466 17650 5468
rect 17674 5466 17730 5468
rect 17434 5414 17480 5466
rect 17480 5414 17490 5466
rect 17514 5414 17544 5466
rect 17544 5414 17556 5466
rect 17556 5414 17570 5466
rect 17594 5414 17608 5466
rect 17608 5414 17620 5466
rect 17620 5414 17650 5466
rect 17674 5414 17684 5466
rect 17684 5414 17730 5466
rect 17434 5412 17490 5414
rect 17514 5412 17570 5414
rect 17594 5412 17650 5414
rect 17674 5412 17730 5414
rect 18510 5228 18566 5264
rect 18510 5208 18512 5228
rect 18512 5208 18564 5228
rect 18564 5208 18566 5228
rect 14334 4378 14390 4380
rect 14414 4378 14470 4380
rect 14494 4378 14550 4380
rect 14574 4378 14630 4380
rect 14334 4326 14380 4378
rect 14380 4326 14390 4378
rect 14414 4326 14444 4378
rect 14444 4326 14456 4378
rect 14456 4326 14470 4378
rect 14494 4326 14508 4378
rect 14508 4326 14520 4378
rect 14520 4326 14550 4378
rect 14574 4326 14584 4378
rect 14584 4326 14630 4378
rect 14334 4324 14390 4326
rect 14414 4324 14470 4326
rect 14494 4324 14550 4326
rect 14574 4324 14630 4326
rect 11234 1114 11290 1116
rect 11314 1114 11370 1116
rect 11394 1114 11450 1116
rect 11474 1114 11530 1116
rect 11234 1062 11280 1114
rect 11280 1062 11290 1114
rect 11314 1062 11344 1114
rect 11344 1062 11356 1114
rect 11356 1062 11370 1114
rect 11394 1062 11408 1114
rect 11408 1062 11420 1114
rect 11420 1062 11450 1114
rect 11474 1062 11484 1114
rect 11484 1062 11530 1114
rect 11234 1060 11290 1062
rect 11314 1060 11370 1062
rect 11394 1060 11450 1062
rect 11474 1060 11530 1062
rect 13082 1264 13138 1320
rect 9684 570 9740 572
rect 9764 570 9820 572
rect 9844 570 9900 572
rect 9924 570 9980 572
rect 9684 518 9730 570
rect 9730 518 9740 570
rect 9764 518 9794 570
rect 9794 518 9806 570
rect 9806 518 9820 570
rect 9844 518 9858 570
rect 9858 518 9870 570
rect 9870 518 9900 570
rect 9924 518 9934 570
rect 9934 518 9980 570
rect 9684 516 9740 518
rect 9764 516 9820 518
rect 9844 516 9900 518
rect 9924 516 9980 518
rect 9034 312 9090 368
rect 12784 570 12840 572
rect 12864 570 12920 572
rect 12944 570 13000 572
rect 13024 570 13080 572
rect 12784 518 12830 570
rect 12830 518 12840 570
rect 12864 518 12894 570
rect 12894 518 12906 570
rect 12906 518 12920 570
rect 12944 518 12958 570
rect 12958 518 12970 570
rect 12970 518 13000 570
rect 13024 518 13034 570
rect 13034 518 13080 570
rect 12784 516 12840 518
rect 12864 516 12920 518
rect 12944 516 13000 518
rect 13024 516 13080 518
rect 14334 3290 14390 3292
rect 14414 3290 14470 3292
rect 14494 3290 14550 3292
rect 14574 3290 14630 3292
rect 14334 3238 14380 3290
rect 14380 3238 14390 3290
rect 14414 3238 14444 3290
rect 14444 3238 14456 3290
rect 14456 3238 14470 3290
rect 14494 3238 14508 3290
rect 14508 3238 14520 3290
rect 14520 3238 14550 3290
rect 14574 3238 14584 3290
rect 14584 3238 14630 3290
rect 14334 3236 14390 3238
rect 14414 3236 14470 3238
rect 14494 3236 14550 3238
rect 14574 3236 14630 3238
rect 14334 2202 14390 2204
rect 14414 2202 14470 2204
rect 14494 2202 14550 2204
rect 14574 2202 14630 2204
rect 14334 2150 14380 2202
rect 14380 2150 14390 2202
rect 14414 2150 14444 2202
rect 14444 2150 14456 2202
rect 14456 2150 14470 2202
rect 14494 2150 14508 2202
rect 14508 2150 14520 2202
rect 14520 2150 14550 2202
rect 14574 2150 14584 2202
rect 14584 2150 14630 2202
rect 14334 2148 14390 2150
rect 14414 2148 14470 2150
rect 14494 2148 14550 2150
rect 14574 2148 14630 2150
rect 13818 876 13874 912
rect 13818 856 13820 876
rect 13820 856 13872 876
rect 13872 856 13874 876
rect 14334 1114 14390 1116
rect 14414 1114 14470 1116
rect 14494 1114 14550 1116
rect 14574 1114 14630 1116
rect 14334 1062 14380 1114
rect 14380 1062 14390 1114
rect 14414 1062 14444 1114
rect 14444 1062 14456 1114
rect 14456 1062 14470 1114
rect 14494 1062 14508 1114
rect 14508 1062 14520 1114
rect 14520 1062 14550 1114
rect 14574 1062 14584 1114
rect 14584 1062 14630 1114
rect 14334 1060 14390 1062
rect 14414 1060 14470 1062
rect 14494 1060 14550 1062
rect 14574 1060 14630 1062
rect 15884 3834 15940 3836
rect 15964 3834 16020 3836
rect 16044 3834 16100 3836
rect 16124 3834 16180 3836
rect 15884 3782 15930 3834
rect 15930 3782 15940 3834
rect 15964 3782 15994 3834
rect 15994 3782 16006 3834
rect 16006 3782 16020 3834
rect 16044 3782 16058 3834
rect 16058 3782 16070 3834
rect 16070 3782 16100 3834
rect 16124 3782 16134 3834
rect 16134 3782 16180 3834
rect 15884 3780 15940 3782
rect 15964 3780 16020 3782
rect 16044 3780 16100 3782
rect 16124 3780 16180 3782
rect 17434 4378 17490 4380
rect 17514 4378 17570 4380
rect 17594 4378 17650 4380
rect 17674 4378 17730 4380
rect 17434 4326 17480 4378
rect 17480 4326 17490 4378
rect 17514 4326 17544 4378
rect 17544 4326 17556 4378
rect 17556 4326 17570 4378
rect 17594 4326 17608 4378
rect 17608 4326 17620 4378
rect 17620 4326 17650 4378
rect 17674 4326 17684 4378
rect 17684 4326 17730 4378
rect 17434 4324 17490 4326
rect 17514 4324 17570 4326
rect 17594 4324 17650 4326
rect 17674 4324 17730 4326
rect 15884 2746 15940 2748
rect 15964 2746 16020 2748
rect 16044 2746 16100 2748
rect 16124 2746 16180 2748
rect 15884 2694 15930 2746
rect 15930 2694 15940 2746
rect 15964 2694 15994 2746
rect 15994 2694 16006 2746
rect 16006 2694 16020 2746
rect 16044 2694 16058 2746
rect 16058 2694 16070 2746
rect 16070 2694 16100 2746
rect 16124 2694 16134 2746
rect 16134 2694 16180 2746
rect 15884 2692 15940 2694
rect 15964 2692 16020 2694
rect 16044 2692 16100 2694
rect 16124 2692 16180 2694
rect 15884 1658 15940 1660
rect 15964 1658 16020 1660
rect 16044 1658 16100 1660
rect 16124 1658 16180 1660
rect 15884 1606 15930 1658
rect 15930 1606 15940 1658
rect 15964 1606 15994 1658
rect 15994 1606 16006 1658
rect 16006 1606 16020 1658
rect 16044 1606 16058 1658
rect 16058 1606 16070 1658
rect 16070 1606 16100 1658
rect 16124 1606 16134 1658
rect 16134 1606 16180 1658
rect 15884 1604 15940 1606
rect 15964 1604 16020 1606
rect 16044 1604 16100 1606
rect 16124 1604 16180 1606
rect 17434 3290 17490 3292
rect 17514 3290 17570 3292
rect 17594 3290 17650 3292
rect 17674 3290 17730 3292
rect 17434 3238 17480 3290
rect 17480 3238 17490 3290
rect 17514 3238 17544 3290
rect 17544 3238 17556 3290
rect 17556 3238 17570 3290
rect 17594 3238 17608 3290
rect 17608 3238 17620 3290
rect 17620 3238 17650 3290
rect 17674 3238 17684 3290
rect 17684 3238 17730 3290
rect 17434 3236 17490 3238
rect 17514 3236 17570 3238
rect 17594 3236 17650 3238
rect 17674 3236 17730 3238
rect 17434 2202 17490 2204
rect 17514 2202 17570 2204
rect 17594 2202 17650 2204
rect 17674 2202 17730 2204
rect 17434 2150 17480 2202
rect 17480 2150 17490 2202
rect 17514 2150 17544 2202
rect 17544 2150 17556 2202
rect 17556 2150 17570 2202
rect 17594 2150 17608 2202
rect 17608 2150 17620 2202
rect 17620 2150 17650 2202
rect 17674 2150 17684 2202
rect 17684 2150 17730 2202
rect 17434 2148 17490 2150
rect 17514 2148 17570 2150
rect 17594 2148 17650 2150
rect 17674 2148 17730 2150
rect 15884 570 15940 572
rect 15964 570 16020 572
rect 16044 570 16100 572
rect 16124 570 16180 572
rect 15884 518 15930 570
rect 15930 518 15940 570
rect 15964 518 15994 570
rect 15994 518 16006 570
rect 16006 518 16020 570
rect 16044 518 16058 570
rect 16058 518 16070 570
rect 16070 518 16100 570
rect 16124 518 16134 570
rect 16134 518 16180 570
rect 15884 516 15940 518
rect 15964 516 16020 518
rect 16044 516 16100 518
rect 16124 516 16180 518
rect 18510 3712 18566 3768
rect 18510 2216 18566 2272
rect 17434 1114 17490 1116
rect 17514 1114 17570 1116
rect 17594 1114 17650 1116
rect 17674 1114 17730 1116
rect 17434 1062 17480 1114
rect 17480 1062 17490 1114
rect 17514 1062 17544 1114
rect 17544 1062 17556 1114
rect 17556 1062 17570 1114
rect 17594 1062 17608 1114
rect 17608 1062 17620 1114
rect 17620 1062 17650 1114
rect 17674 1062 17684 1114
rect 17684 1062 17730 1114
rect 17434 1060 17490 1062
rect 17514 1060 17570 1062
rect 17594 1060 17650 1062
rect 17674 1060 17730 1062
rect 18510 720 18566 776
rect 5034 26 5090 28
rect 5114 26 5170 28
rect 5194 26 5250 28
rect 5274 26 5330 28
rect 5034 -26 5080 26
rect 5080 -26 5090 26
rect 5114 -26 5144 26
rect 5144 -26 5156 26
rect 5156 -26 5170 26
rect 5194 -26 5208 26
rect 5208 -26 5220 26
rect 5220 -26 5250 26
rect 5274 -26 5284 26
rect 5284 -26 5330 26
rect 5034 -28 5090 -26
rect 5114 -28 5170 -26
rect 5194 -28 5250 -26
rect 5274 -28 5330 -26
rect 8134 26 8190 28
rect 8214 26 8270 28
rect 8294 26 8350 28
rect 8374 26 8430 28
rect 8134 -26 8180 26
rect 8180 -26 8190 26
rect 8214 -26 8244 26
rect 8244 -26 8256 26
rect 8256 -26 8270 26
rect 8294 -26 8308 26
rect 8308 -26 8320 26
rect 8320 -26 8350 26
rect 8374 -26 8384 26
rect 8384 -26 8430 26
rect 8134 -28 8190 -26
rect 8214 -28 8270 -26
rect 8294 -28 8350 -26
rect 8374 -28 8430 -26
rect 11234 26 11290 28
rect 11314 26 11370 28
rect 11394 26 11450 28
rect 11474 26 11530 28
rect 11234 -26 11280 26
rect 11280 -26 11290 26
rect 11314 -26 11344 26
rect 11344 -26 11356 26
rect 11356 -26 11370 26
rect 11394 -26 11408 26
rect 11408 -26 11420 26
rect 11420 -26 11450 26
rect 11474 -26 11484 26
rect 11484 -26 11530 26
rect 11234 -28 11290 -26
rect 11314 -28 11370 -26
rect 11394 -28 11450 -26
rect 11474 -28 11530 -26
rect 14334 26 14390 28
rect 14414 26 14470 28
rect 14494 26 14550 28
rect 14574 26 14630 28
rect 14334 -26 14380 26
rect 14380 -26 14390 26
rect 14414 -26 14444 26
rect 14444 -26 14456 26
rect 14456 -26 14470 26
rect 14494 -26 14508 26
rect 14508 -26 14520 26
rect 14520 -26 14550 26
rect 14574 -26 14584 26
rect 14584 -26 14630 26
rect 14334 -28 14390 -26
rect 14414 -28 14470 -26
rect 14494 -28 14550 -26
rect 14574 -28 14630 -26
rect 17434 26 17490 28
rect 17514 26 17570 28
rect 17594 26 17650 28
rect 17674 26 17730 28
rect 17434 -26 17480 26
rect 17480 -26 17490 26
rect 17514 -26 17544 26
rect 17544 -26 17556 26
rect 17556 -26 17570 26
rect 17594 -26 17608 26
rect 17608 -26 17620 26
rect 17620 -26 17650 26
rect 17674 -26 17684 26
rect 17684 -26 17730 26
rect 17434 -28 17490 -26
rect 17514 -28 17570 -26
rect 17594 -28 17650 -26
rect 17674 -28 17730 -26
<< metal3 >>
rect 18781 11250 18847 11253
rect 19200 11250 20000 11280
rect 18781 11248 20000 11250
rect 18781 11192 18786 11248
rect 18842 11192 20000 11248
rect 18781 11190 20000 11192
rect 18781 11187 18847 11190
rect 19200 11160 20000 11190
rect 5022 10912 5342 10913
rect 5022 10848 5030 10912
rect 5094 10848 5110 10912
rect 5174 10848 5190 10912
rect 5254 10848 5270 10912
rect 5334 10848 5342 10912
rect 5022 10847 5342 10848
rect 8122 10912 8442 10913
rect 8122 10848 8130 10912
rect 8194 10848 8210 10912
rect 8274 10848 8290 10912
rect 8354 10848 8370 10912
rect 8434 10848 8442 10912
rect 8122 10847 8442 10848
rect 11222 10912 11542 10913
rect 11222 10848 11230 10912
rect 11294 10848 11310 10912
rect 11374 10848 11390 10912
rect 11454 10848 11470 10912
rect 11534 10848 11542 10912
rect 11222 10847 11542 10848
rect 14322 10912 14642 10913
rect 14322 10848 14330 10912
rect 14394 10848 14410 10912
rect 14474 10848 14490 10912
rect 14554 10848 14570 10912
rect 14634 10848 14642 10912
rect 14322 10847 14642 10848
rect 17422 10912 17742 10913
rect 17422 10848 17430 10912
rect 17494 10848 17510 10912
rect 17574 10848 17590 10912
rect 17654 10848 17670 10912
rect 17734 10848 17742 10912
rect 17422 10847 17742 10848
rect 3472 10368 3792 10369
rect 3472 10304 3480 10368
rect 3544 10304 3560 10368
rect 3624 10304 3640 10368
rect 3704 10304 3720 10368
rect 3784 10304 3792 10368
rect 3472 10303 3792 10304
rect 6572 10368 6892 10369
rect 6572 10304 6580 10368
rect 6644 10304 6660 10368
rect 6724 10304 6740 10368
rect 6804 10304 6820 10368
rect 6884 10304 6892 10368
rect 6572 10303 6892 10304
rect 9672 10368 9992 10369
rect 9672 10304 9680 10368
rect 9744 10304 9760 10368
rect 9824 10304 9840 10368
rect 9904 10304 9920 10368
rect 9984 10304 9992 10368
rect 9672 10303 9992 10304
rect 12772 10368 13092 10369
rect 12772 10304 12780 10368
rect 12844 10304 12860 10368
rect 12924 10304 12940 10368
rect 13004 10304 13020 10368
rect 13084 10304 13092 10368
rect 12772 10303 13092 10304
rect 15872 10368 16192 10369
rect 15872 10304 15880 10368
rect 15944 10304 15960 10368
rect 16024 10304 16040 10368
rect 16104 10304 16120 10368
rect 16184 10304 16192 10368
rect 15872 10303 16192 10304
rect 5022 9824 5342 9825
rect 5022 9760 5030 9824
rect 5094 9760 5110 9824
rect 5174 9760 5190 9824
rect 5254 9760 5270 9824
rect 5334 9760 5342 9824
rect 5022 9759 5342 9760
rect 8122 9824 8442 9825
rect 8122 9760 8130 9824
rect 8194 9760 8210 9824
rect 8274 9760 8290 9824
rect 8354 9760 8370 9824
rect 8434 9760 8442 9824
rect 8122 9759 8442 9760
rect 11222 9824 11542 9825
rect 11222 9760 11230 9824
rect 11294 9760 11310 9824
rect 11374 9760 11390 9824
rect 11454 9760 11470 9824
rect 11534 9760 11542 9824
rect 11222 9759 11542 9760
rect 14322 9824 14642 9825
rect 14322 9760 14330 9824
rect 14394 9760 14410 9824
rect 14474 9760 14490 9824
rect 14554 9760 14570 9824
rect 14634 9760 14642 9824
rect 14322 9759 14642 9760
rect 17422 9824 17742 9825
rect 17422 9760 17430 9824
rect 17494 9760 17510 9824
rect 17574 9760 17590 9824
rect 17654 9760 17670 9824
rect 17734 9760 17742 9824
rect 17422 9759 17742 9760
rect 18689 9754 18755 9757
rect 19200 9754 20000 9784
rect 18689 9752 20000 9754
rect 18689 9696 18694 9752
rect 18750 9696 20000 9752
rect 18689 9694 20000 9696
rect 18689 9691 18755 9694
rect 19200 9664 20000 9694
rect 3472 9280 3792 9281
rect 3472 9216 3480 9280
rect 3544 9216 3560 9280
rect 3624 9216 3640 9280
rect 3704 9216 3720 9280
rect 3784 9216 3792 9280
rect 3472 9215 3792 9216
rect 6572 9280 6892 9281
rect 6572 9216 6580 9280
rect 6644 9216 6660 9280
rect 6724 9216 6740 9280
rect 6804 9216 6820 9280
rect 6884 9216 6892 9280
rect 6572 9215 6892 9216
rect 9672 9280 9992 9281
rect 9672 9216 9680 9280
rect 9744 9216 9760 9280
rect 9824 9216 9840 9280
rect 9904 9216 9920 9280
rect 9984 9216 9992 9280
rect 9672 9215 9992 9216
rect 12772 9280 13092 9281
rect 12772 9216 12780 9280
rect 12844 9216 12860 9280
rect 12924 9216 12940 9280
rect 13004 9216 13020 9280
rect 13084 9216 13092 9280
rect 12772 9215 13092 9216
rect 15872 9280 16192 9281
rect 15872 9216 15880 9280
rect 15944 9216 15960 9280
rect 16024 9216 16040 9280
rect 16104 9216 16120 9280
rect 16184 9216 16192 9280
rect 15872 9215 16192 9216
rect 5022 8736 5342 8737
rect 5022 8672 5030 8736
rect 5094 8672 5110 8736
rect 5174 8672 5190 8736
rect 5254 8672 5270 8736
rect 5334 8672 5342 8736
rect 5022 8671 5342 8672
rect 8122 8736 8442 8737
rect 8122 8672 8130 8736
rect 8194 8672 8210 8736
rect 8274 8672 8290 8736
rect 8354 8672 8370 8736
rect 8434 8672 8442 8736
rect 8122 8671 8442 8672
rect 11222 8736 11542 8737
rect 11222 8672 11230 8736
rect 11294 8672 11310 8736
rect 11374 8672 11390 8736
rect 11454 8672 11470 8736
rect 11534 8672 11542 8736
rect 11222 8671 11542 8672
rect 14322 8736 14642 8737
rect 14322 8672 14330 8736
rect 14394 8672 14410 8736
rect 14474 8672 14490 8736
rect 14554 8672 14570 8736
rect 14634 8672 14642 8736
rect 14322 8671 14642 8672
rect 17422 8736 17742 8737
rect 17422 8672 17430 8736
rect 17494 8672 17510 8736
rect 17574 8672 17590 8736
rect 17654 8672 17670 8736
rect 17734 8672 17742 8736
rect 17422 8671 17742 8672
rect 18597 8258 18663 8261
rect 19200 8258 20000 8288
rect 18597 8256 20000 8258
rect 18597 8200 18602 8256
rect 18658 8200 20000 8256
rect 18597 8198 20000 8200
rect 18597 8195 18663 8198
rect 3472 8192 3792 8193
rect 3472 8128 3480 8192
rect 3544 8128 3560 8192
rect 3624 8128 3640 8192
rect 3704 8128 3720 8192
rect 3784 8128 3792 8192
rect 3472 8127 3792 8128
rect 6572 8192 6892 8193
rect 6572 8128 6580 8192
rect 6644 8128 6660 8192
rect 6724 8128 6740 8192
rect 6804 8128 6820 8192
rect 6884 8128 6892 8192
rect 6572 8127 6892 8128
rect 9672 8192 9992 8193
rect 9672 8128 9680 8192
rect 9744 8128 9760 8192
rect 9824 8128 9840 8192
rect 9904 8128 9920 8192
rect 9984 8128 9992 8192
rect 9672 8127 9992 8128
rect 12772 8192 13092 8193
rect 12772 8128 12780 8192
rect 12844 8128 12860 8192
rect 12924 8128 12940 8192
rect 13004 8128 13020 8192
rect 13084 8128 13092 8192
rect 12772 8127 13092 8128
rect 15872 8192 16192 8193
rect 15872 8128 15880 8192
rect 15944 8128 15960 8192
rect 16024 8128 16040 8192
rect 16104 8128 16120 8192
rect 16184 8128 16192 8192
rect 19200 8168 20000 8198
rect 15872 8127 16192 8128
rect 11329 7986 11395 7989
rect 15101 7986 15167 7989
rect 11329 7984 15167 7986
rect 11329 7928 11334 7984
rect 11390 7928 15106 7984
rect 15162 7928 15167 7984
rect 11329 7926 15167 7928
rect 11329 7923 11395 7926
rect 15101 7923 15167 7926
rect 5022 7648 5342 7649
rect 5022 7584 5030 7648
rect 5094 7584 5110 7648
rect 5174 7584 5190 7648
rect 5254 7584 5270 7648
rect 5334 7584 5342 7648
rect 5022 7583 5342 7584
rect 8122 7648 8442 7649
rect 8122 7584 8130 7648
rect 8194 7584 8210 7648
rect 8274 7584 8290 7648
rect 8354 7584 8370 7648
rect 8434 7584 8442 7648
rect 8122 7583 8442 7584
rect 11222 7648 11542 7649
rect 11222 7584 11230 7648
rect 11294 7584 11310 7648
rect 11374 7584 11390 7648
rect 11454 7584 11470 7648
rect 11534 7584 11542 7648
rect 11222 7583 11542 7584
rect 14322 7648 14642 7649
rect 14322 7584 14330 7648
rect 14394 7584 14410 7648
rect 14474 7584 14490 7648
rect 14554 7584 14570 7648
rect 14634 7584 14642 7648
rect 14322 7583 14642 7584
rect 17422 7648 17742 7649
rect 17422 7584 17430 7648
rect 17494 7584 17510 7648
rect 17574 7584 17590 7648
rect 17654 7584 17670 7648
rect 17734 7584 17742 7648
rect 17422 7583 17742 7584
rect 10041 7442 10107 7445
rect 10409 7442 10475 7445
rect 10041 7440 10475 7442
rect 10041 7384 10046 7440
rect 10102 7384 10414 7440
rect 10470 7384 10475 7440
rect 10041 7382 10475 7384
rect 10041 7379 10107 7382
rect 10409 7379 10475 7382
rect 10593 7442 10659 7445
rect 13997 7442 14063 7445
rect 10593 7440 14063 7442
rect 10593 7384 10598 7440
rect 10654 7384 14002 7440
rect 14058 7384 14063 7440
rect 10593 7382 14063 7384
rect 10593 7379 10659 7382
rect 13997 7379 14063 7382
rect 10409 7306 10475 7309
rect 12709 7306 12775 7309
rect 10409 7304 12775 7306
rect 10409 7248 10414 7304
rect 10470 7248 12714 7304
rect 12770 7248 12775 7304
rect 10409 7246 12775 7248
rect 10409 7243 10475 7246
rect 12709 7243 12775 7246
rect 3472 7104 3792 7105
rect 3472 7040 3480 7104
rect 3544 7040 3560 7104
rect 3624 7040 3640 7104
rect 3704 7040 3720 7104
rect 3784 7040 3792 7104
rect 3472 7039 3792 7040
rect 6572 7104 6892 7105
rect 6572 7040 6580 7104
rect 6644 7040 6660 7104
rect 6724 7040 6740 7104
rect 6804 7040 6820 7104
rect 6884 7040 6892 7104
rect 6572 7039 6892 7040
rect 9672 7104 9992 7105
rect 9672 7040 9680 7104
rect 9744 7040 9760 7104
rect 9824 7040 9840 7104
rect 9904 7040 9920 7104
rect 9984 7040 9992 7104
rect 9672 7039 9992 7040
rect 12772 7104 13092 7105
rect 12772 7040 12780 7104
rect 12844 7040 12860 7104
rect 12924 7040 12940 7104
rect 13004 7040 13020 7104
rect 13084 7040 13092 7104
rect 12772 7039 13092 7040
rect 15872 7104 16192 7105
rect 15872 7040 15880 7104
rect 15944 7040 15960 7104
rect 16024 7040 16040 7104
rect 16104 7040 16120 7104
rect 16184 7040 16192 7104
rect 15872 7039 16192 7040
rect 10225 6898 10291 6901
rect 10685 6898 10751 6901
rect 10225 6896 10751 6898
rect 10225 6840 10230 6896
rect 10286 6840 10690 6896
rect 10746 6840 10751 6896
rect 10225 6838 10751 6840
rect 10225 6835 10291 6838
rect 10685 6835 10751 6838
rect 10409 6762 10475 6765
rect 11053 6762 11119 6765
rect 10409 6760 11119 6762
rect 10409 6704 10414 6760
rect 10470 6704 11058 6760
rect 11114 6704 11119 6760
rect 10409 6702 11119 6704
rect 10409 6699 10475 6702
rect 11053 6699 11119 6702
rect 18505 6762 18571 6765
rect 19200 6762 20000 6792
rect 18505 6760 20000 6762
rect 18505 6704 18510 6760
rect 18566 6704 20000 6760
rect 18505 6702 20000 6704
rect 18505 6699 18571 6702
rect 19200 6672 20000 6702
rect 5022 6560 5342 6561
rect 5022 6496 5030 6560
rect 5094 6496 5110 6560
rect 5174 6496 5190 6560
rect 5254 6496 5270 6560
rect 5334 6496 5342 6560
rect 5022 6495 5342 6496
rect 8122 6560 8442 6561
rect 8122 6496 8130 6560
rect 8194 6496 8210 6560
rect 8274 6496 8290 6560
rect 8354 6496 8370 6560
rect 8434 6496 8442 6560
rect 8122 6495 8442 6496
rect 11222 6560 11542 6561
rect 11222 6496 11230 6560
rect 11294 6496 11310 6560
rect 11374 6496 11390 6560
rect 11454 6496 11470 6560
rect 11534 6496 11542 6560
rect 11222 6495 11542 6496
rect 14322 6560 14642 6561
rect 14322 6496 14330 6560
rect 14394 6496 14410 6560
rect 14474 6496 14490 6560
rect 14554 6496 14570 6560
rect 14634 6496 14642 6560
rect 14322 6495 14642 6496
rect 17422 6560 17742 6561
rect 17422 6496 17430 6560
rect 17494 6496 17510 6560
rect 17574 6496 17590 6560
rect 17654 6496 17670 6560
rect 17734 6496 17742 6560
rect 17422 6495 17742 6496
rect 3472 6016 3792 6017
rect 3472 5952 3480 6016
rect 3544 5952 3560 6016
rect 3624 5952 3640 6016
rect 3704 5952 3720 6016
rect 3784 5952 3792 6016
rect 3472 5951 3792 5952
rect 6572 6016 6892 6017
rect 6572 5952 6580 6016
rect 6644 5952 6660 6016
rect 6724 5952 6740 6016
rect 6804 5952 6820 6016
rect 6884 5952 6892 6016
rect 6572 5951 6892 5952
rect 9672 6016 9992 6017
rect 9672 5952 9680 6016
rect 9744 5952 9760 6016
rect 9824 5952 9840 6016
rect 9904 5952 9920 6016
rect 9984 5952 9992 6016
rect 9672 5951 9992 5952
rect 12772 6016 13092 6017
rect 12772 5952 12780 6016
rect 12844 5952 12860 6016
rect 12924 5952 12940 6016
rect 13004 5952 13020 6016
rect 13084 5952 13092 6016
rect 12772 5951 13092 5952
rect 15872 6016 16192 6017
rect 15872 5952 15880 6016
rect 15944 5952 15960 6016
rect 16024 5952 16040 6016
rect 16104 5952 16120 6016
rect 16184 5952 16192 6016
rect 15872 5951 16192 5952
rect 5022 5472 5342 5473
rect 5022 5408 5030 5472
rect 5094 5408 5110 5472
rect 5174 5408 5190 5472
rect 5254 5408 5270 5472
rect 5334 5408 5342 5472
rect 5022 5407 5342 5408
rect 8122 5472 8442 5473
rect 8122 5408 8130 5472
rect 8194 5408 8210 5472
rect 8274 5408 8290 5472
rect 8354 5408 8370 5472
rect 8434 5408 8442 5472
rect 8122 5407 8442 5408
rect 11222 5472 11542 5473
rect 11222 5408 11230 5472
rect 11294 5408 11310 5472
rect 11374 5408 11390 5472
rect 11454 5408 11470 5472
rect 11534 5408 11542 5472
rect 11222 5407 11542 5408
rect 14322 5472 14642 5473
rect 14322 5408 14330 5472
rect 14394 5408 14410 5472
rect 14474 5408 14490 5472
rect 14554 5408 14570 5472
rect 14634 5408 14642 5472
rect 14322 5407 14642 5408
rect 17422 5472 17742 5473
rect 17422 5408 17430 5472
rect 17494 5408 17510 5472
rect 17574 5408 17590 5472
rect 17654 5408 17670 5472
rect 17734 5408 17742 5472
rect 17422 5407 17742 5408
rect 18505 5266 18571 5269
rect 19200 5266 20000 5296
rect 18505 5264 20000 5266
rect 18505 5208 18510 5264
rect 18566 5208 20000 5264
rect 18505 5206 20000 5208
rect 18505 5203 18571 5206
rect 19200 5176 20000 5206
rect 3472 4928 3792 4929
rect 3472 4864 3480 4928
rect 3544 4864 3560 4928
rect 3624 4864 3640 4928
rect 3704 4864 3720 4928
rect 3784 4864 3792 4928
rect 3472 4863 3792 4864
rect 6572 4928 6892 4929
rect 6572 4864 6580 4928
rect 6644 4864 6660 4928
rect 6724 4864 6740 4928
rect 6804 4864 6820 4928
rect 6884 4864 6892 4928
rect 6572 4863 6892 4864
rect 9672 4928 9992 4929
rect 9672 4864 9680 4928
rect 9744 4864 9760 4928
rect 9824 4864 9840 4928
rect 9904 4864 9920 4928
rect 9984 4864 9992 4928
rect 9672 4863 9992 4864
rect 12772 4928 13092 4929
rect 12772 4864 12780 4928
rect 12844 4864 12860 4928
rect 12924 4864 12940 4928
rect 13004 4864 13020 4928
rect 13084 4864 13092 4928
rect 12772 4863 13092 4864
rect 15872 4928 16192 4929
rect 15872 4864 15880 4928
rect 15944 4864 15960 4928
rect 16024 4864 16040 4928
rect 16104 4864 16120 4928
rect 16184 4864 16192 4928
rect 15872 4863 16192 4864
rect 5022 4384 5342 4385
rect 5022 4320 5030 4384
rect 5094 4320 5110 4384
rect 5174 4320 5190 4384
rect 5254 4320 5270 4384
rect 5334 4320 5342 4384
rect 5022 4319 5342 4320
rect 8122 4384 8442 4385
rect 8122 4320 8130 4384
rect 8194 4320 8210 4384
rect 8274 4320 8290 4384
rect 8354 4320 8370 4384
rect 8434 4320 8442 4384
rect 8122 4319 8442 4320
rect 11222 4384 11542 4385
rect 11222 4320 11230 4384
rect 11294 4320 11310 4384
rect 11374 4320 11390 4384
rect 11454 4320 11470 4384
rect 11534 4320 11542 4384
rect 11222 4319 11542 4320
rect 14322 4384 14642 4385
rect 14322 4320 14330 4384
rect 14394 4320 14410 4384
rect 14474 4320 14490 4384
rect 14554 4320 14570 4384
rect 14634 4320 14642 4384
rect 14322 4319 14642 4320
rect 17422 4384 17742 4385
rect 17422 4320 17430 4384
rect 17494 4320 17510 4384
rect 17574 4320 17590 4384
rect 17654 4320 17670 4384
rect 17734 4320 17742 4384
rect 17422 4319 17742 4320
rect 3472 3840 3792 3841
rect 3472 3776 3480 3840
rect 3544 3776 3560 3840
rect 3624 3776 3640 3840
rect 3704 3776 3720 3840
rect 3784 3776 3792 3840
rect 3472 3775 3792 3776
rect 6572 3840 6892 3841
rect 6572 3776 6580 3840
rect 6644 3776 6660 3840
rect 6724 3776 6740 3840
rect 6804 3776 6820 3840
rect 6884 3776 6892 3840
rect 6572 3775 6892 3776
rect 9672 3840 9992 3841
rect 9672 3776 9680 3840
rect 9744 3776 9760 3840
rect 9824 3776 9840 3840
rect 9904 3776 9920 3840
rect 9984 3776 9992 3840
rect 9672 3775 9992 3776
rect 12772 3840 13092 3841
rect 12772 3776 12780 3840
rect 12844 3776 12860 3840
rect 12924 3776 12940 3840
rect 13004 3776 13020 3840
rect 13084 3776 13092 3840
rect 12772 3775 13092 3776
rect 15872 3840 16192 3841
rect 15872 3776 15880 3840
rect 15944 3776 15960 3840
rect 16024 3776 16040 3840
rect 16104 3776 16120 3840
rect 16184 3776 16192 3840
rect 15872 3775 16192 3776
rect 18505 3770 18571 3773
rect 19200 3770 20000 3800
rect 18505 3768 20000 3770
rect 18505 3712 18510 3768
rect 18566 3712 20000 3768
rect 18505 3710 20000 3712
rect 18505 3707 18571 3710
rect 19200 3680 20000 3710
rect 5022 3296 5342 3297
rect 5022 3232 5030 3296
rect 5094 3232 5110 3296
rect 5174 3232 5190 3296
rect 5254 3232 5270 3296
rect 5334 3232 5342 3296
rect 5022 3231 5342 3232
rect 8122 3296 8442 3297
rect 8122 3232 8130 3296
rect 8194 3232 8210 3296
rect 8274 3232 8290 3296
rect 8354 3232 8370 3296
rect 8434 3232 8442 3296
rect 8122 3231 8442 3232
rect 11222 3296 11542 3297
rect 11222 3232 11230 3296
rect 11294 3232 11310 3296
rect 11374 3232 11390 3296
rect 11454 3232 11470 3296
rect 11534 3232 11542 3296
rect 11222 3231 11542 3232
rect 14322 3296 14642 3297
rect 14322 3232 14330 3296
rect 14394 3232 14410 3296
rect 14474 3232 14490 3296
rect 14554 3232 14570 3296
rect 14634 3232 14642 3296
rect 14322 3231 14642 3232
rect 17422 3296 17742 3297
rect 17422 3232 17430 3296
rect 17494 3232 17510 3296
rect 17574 3232 17590 3296
rect 17654 3232 17670 3296
rect 17734 3232 17742 3296
rect 17422 3231 17742 3232
rect 3472 2752 3792 2753
rect 3472 2688 3480 2752
rect 3544 2688 3560 2752
rect 3624 2688 3640 2752
rect 3704 2688 3720 2752
rect 3784 2688 3792 2752
rect 3472 2687 3792 2688
rect 6572 2752 6892 2753
rect 6572 2688 6580 2752
rect 6644 2688 6660 2752
rect 6724 2688 6740 2752
rect 6804 2688 6820 2752
rect 6884 2688 6892 2752
rect 6572 2687 6892 2688
rect 9672 2752 9992 2753
rect 9672 2688 9680 2752
rect 9744 2688 9760 2752
rect 9824 2688 9840 2752
rect 9904 2688 9920 2752
rect 9984 2688 9992 2752
rect 9672 2687 9992 2688
rect 12772 2752 13092 2753
rect 12772 2688 12780 2752
rect 12844 2688 12860 2752
rect 12924 2688 12940 2752
rect 13004 2688 13020 2752
rect 13084 2688 13092 2752
rect 12772 2687 13092 2688
rect 15872 2752 16192 2753
rect 15872 2688 15880 2752
rect 15944 2688 15960 2752
rect 16024 2688 16040 2752
rect 16104 2688 16120 2752
rect 16184 2688 16192 2752
rect 15872 2687 16192 2688
rect 18505 2274 18571 2277
rect 19200 2274 20000 2304
rect 18505 2272 20000 2274
rect 18505 2216 18510 2272
rect 18566 2216 20000 2272
rect 18505 2214 20000 2216
rect 18505 2211 18571 2214
rect 5022 2208 5342 2209
rect 5022 2144 5030 2208
rect 5094 2144 5110 2208
rect 5174 2144 5190 2208
rect 5254 2144 5270 2208
rect 5334 2144 5342 2208
rect 5022 2143 5342 2144
rect 8122 2208 8442 2209
rect 8122 2144 8130 2208
rect 8194 2144 8210 2208
rect 8274 2144 8290 2208
rect 8354 2144 8370 2208
rect 8434 2144 8442 2208
rect 8122 2143 8442 2144
rect 11222 2208 11542 2209
rect 11222 2144 11230 2208
rect 11294 2144 11310 2208
rect 11374 2144 11390 2208
rect 11454 2144 11470 2208
rect 11534 2144 11542 2208
rect 11222 2143 11542 2144
rect 14322 2208 14642 2209
rect 14322 2144 14330 2208
rect 14394 2144 14410 2208
rect 14474 2144 14490 2208
rect 14554 2144 14570 2208
rect 14634 2144 14642 2208
rect 14322 2143 14642 2144
rect 17422 2208 17742 2209
rect 17422 2144 17430 2208
rect 17494 2144 17510 2208
rect 17574 2144 17590 2208
rect 17654 2144 17670 2208
rect 17734 2144 17742 2208
rect 19200 2184 20000 2214
rect 17422 2143 17742 2144
rect 2497 2002 2563 2005
rect 4705 2002 4771 2005
rect 2497 2000 4771 2002
rect 2497 1944 2502 2000
rect 2558 1944 4710 2000
rect 4766 1944 4771 2000
rect 2497 1942 4771 1944
rect 2497 1939 2563 1942
rect 4705 1939 4771 1942
rect 3472 1664 3792 1665
rect 3472 1600 3480 1664
rect 3544 1600 3560 1664
rect 3624 1600 3640 1664
rect 3704 1600 3720 1664
rect 3784 1600 3792 1664
rect 3472 1599 3792 1600
rect 6572 1664 6892 1665
rect 6572 1600 6580 1664
rect 6644 1600 6660 1664
rect 6724 1600 6740 1664
rect 6804 1600 6820 1664
rect 6884 1600 6892 1664
rect 6572 1599 6892 1600
rect 9672 1664 9992 1665
rect 9672 1600 9680 1664
rect 9744 1600 9760 1664
rect 9824 1600 9840 1664
rect 9904 1600 9920 1664
rect 9984 1600 9992 1664
rect 9672 1599 9992 1600
rect 12772 1664 13092 1665
rect 12772 1600 12780 1664
rect 12844 1600 12860 1664
rect 12924 1600 12940 1664
rect 13004 1600 13020 1664
rect 13084 1600 13092 1664
rect 12772 1599 13092 1600
rect 15872 1664 16192 1665
rect 15872 1600 15880 1664
rect 15944 1600 15960 1664
rect 16024 1600 16040 1664
rect 16104 1600 16120 1664
rect 16184 1600 16192 1664
rect 15872 1599 16192 1600
rect 8201 1322 8267 1325
rect 10961 1322 11027 1325
rect 13077 1322 13143 1325
rect 8201 1320 13143 1322
rect 8201 1264 8206 1320
rect 8262 1264 10966 1320
rect 11022 1264 13082 1320
rect 13138 1264 13143 1320
rect 8201 1262 13143 1264
rect 8201 1259 8267 1262
rect 10961 1259 11027 1262
rect 13077 1259 13143 1262
rect 5022 1120 5342 1121
rect 5022 1056 5030 1120
rect 5094 1056 5110 1120
rect 5174 1056 5190 1120
rect 5254 1056 5270 1120
rect 5334 1056 5342 1120
rect 5022 1055 5342 1056
rect 8122 1120 8442 1121
rect 8122 1056 8130 1120
rect 8194 1056 8210 1120
rect 8274 1056 8290 1120
rect 8354 1056 8370 1120
rect 8434 1056 8442 1120
rect 8122 1055 8442 1056
rect 11222 1120 11542 1121
rect 11222 1056 11230 1120
rect 11294 1056 11310 1120
rect 11374 1056 11390 1120
rect 11454 1056 11470 1120
rect 11534 1056 11542 1120
rect 11222 1055 11542 1056
rect 14322 1120 14642 1121
rect 14322 1056 14330 1120
rect 14394 1056 14410 1120
rect 14474 1056 14490 1120
rect 14554 1056 14570 1120
rect 14634 1056 14642 1120
rect 14322 1055 14642 1056
rect 17422 1120 17742 1121
rect 17422 1056 17430 1120
rect 17494 1056 17510 1120
rect 17574 1056 17590 1120
rect 17654 1056 17670 1120
rect 17734 1056 17742 1120
rect 17422 1055 17742 1056
rect 3969 914 4035 917
rect 5901 914 5967 917
rect 3969 912 5967 914
rect 3969 856 3974 912
rect 4030 856 5906 912
rect 5962 856 5967 912
rect 3969 854 5967 856
rect 3969 851 4035 854
rect 5901 851 5967 854
rect 10593 914 10659 917
rect 13813 914 13879 917
rect 10593 912 13879 914
rect 10593 856 10598 912
rect 10654 856 13818 912
rect 13874 856 13879 912
rect 10593 854 13879 856
rect 10593 851 10659 854
rect 13813 851 13879 854
rect 18505 778 18571 781
rect 19200 778 20000 808
rect 18505 776 20000 778
rect 18505 720 18510 776
rect 18566 720 20000 776
rect 18505 718 20000 720
rect 18505 715 18571 718
rect 19200 688 20000 718
rect 3472 576 3792 577
rect 3472 512 3480 576
rect 3544 512 3560 576
rect 3624 512 3640 576
rect 3704 512 3720 576
rect 3784 512 3792 576
rect 3472 511 3792 512
rect 6572 576 6892 577
rect 6572 512 6580 576
rect 6644 512 6660 576
rect 6724 512 6740 576
rect 6804 512 6820 576
rect 6884 512 6892 576
rect 6572 511 6892 512
rect 9672 576 9992 577
rect 9672 512 9680 576
rect 9744 512 9760 576
rect 9824 512 9840 576
rect 9904 512 9920 576
rect 9984 512 9992 576
rect 9672 511 9992 512
rect 12772 576 13092 577
rect 12772 512 12780 576
rect 12844 512 12860 576
rect 12924 512 12940 576
rect 13004 512 13020 576
rect 13084 512 13092 576
rect 12772 511 13092 512
rect 15872 576 16192 577
rect 15872 512 15880 576
rect 15944 512 15960 576
rect 16024 512 16040 576
rect 16104 512 16120 576
rect 16184 512 16192 576
rect 15872 511 16192 512
rect 5073 370 5139 373
rect 9029 370 9095 373
rect 5073 368 9095 370
rect 5073 312 5078 368
rect 5134 312 9034 368
rect 9090 312 9095 368
rect 5073 310 9095 312
rect 5073 307 5139 310
rect 9029 307 9095 310
rect 5022 32 5342 33
rect 5022 -32 5030 32
rect 5094 -32 5110 32
rect 5174 -32 5190 32
rect 5254 -32 5270 32
rect 5334 -32 5342 32
rect 5022 -33 5342 -32
rect 8122 32 8442 33
rect 8122 -32 8130 32
rect 8194 -32 8210 32
rect 8274 -32 8290 32
rect 8354 -32 8370 32
rect 8434 -32 8442 32
rect 8122 -33 8442 -32
rect 11222 32 11542 33
rect 11222 -32 11230 32
rect 11294 -32 11310 32
rect 11374 -32 11390 32
rect 11454 -32 11470 32
rect 11534 -32 11542 32
rect 11222 -33 11542 -32
rect 14322 32 14642 33
rect 14322 -32 14330 32
rect 14394 -32 14410 32
rect 14474 -32 14490 32
rect 14554 -32 14570 32
rect 14634 -32 14642 32
rect 14322 -33 14642 -32
rect 17422 32 17742 33
rect 17422 -32 17430 32
rect 17494 -32 17510 32
rect 17574 -32 17590 32
rect 17654 -32 17670 32
rect 17734 -32 17742 32
rect 17422 -33 17742 -32
<< via3 >>
rect 5030 10908 5094 10912
rect 5030 10852 5034 10908
rect 5034 10852 5090 10908
rect 5090 10852 5094 10908
rect 5030 10848 5094 10852
rect 5110 10908 5174 10912
rect 5110 10852 5114 10908
rect 5114 10852 5170 10908
rect 5170 10852 5174 10908
rect 5110 10848 5174 10852
rect 5190 10908 5254 10912
rect 5190 10852 5194 10908
rect 5194 10852 5250 10908
rect 5250 10852 5254 10908
rect 5190 10848 5254 10852
rect 5270 10908 5334 10912
rect 5270 10852 5274 10908
rect 5274 10852 5330 10908
rect 5330 10852 5334 10908
rect 5270 10848 5334 10852
rect 8130 10908 8194 10912
rect 8130 10852 8134 10908
rect 8134 10852 8190 10908
rect 8190 10852 8194 10908
rect 8130 10848 8194 10852
rect 8210 10908 8274 10912
rect 8210 10852 8214 10908
rect 8214 10852 8270 10908
rect 8270 10852 8274 10908
rect 8210 10848 8274 10852
rect 8290 10908 8354 10912
rect 8290 10852 8294 10908
rect 8294 10852 8350 10908
rect 8350 10852 8354 10908
rect 8290 10848 8354 10852
rect 8370 10908 8434 10912
rect 8370 10852 8374 10908
rect 8374 10852 8430 10908
rect 8430 10852 8434 10908
rect 8370 10848 8434 10852
rect 11230 10908 11294 10912
rect 11230 10852 11234 10908
rect 11234 10852 11290 10908
rect 11290 10852 11294 10908
rect 11230 10848 11294 10852
rect 11310 10908 11374 10912
rect 11310 10852 11314 10908
rect 11314 10852 11370 10908
rect 11370 10852 11374 10908
rect 11310 10848 11374 10852
rect 11390 10908 11454 10912
rect 11390 10852 11394 10908
rect 11394 10852 11450 10908
rect 11450 10852 11454 10908
rect 11390 10848 11454 10852
rect 11470 10908 11534 10912
rect 11470 10852 11474 10908
rect 11474 10852 11530 10908
rect 11530 10852 11534 10908
rect 11470 10848 11534 10852
rect 14330 10908 14394 10912
rect 14330 10852 14334 10908
rect 14334 10852 14390 10908
rect 14390 10852 14394 10908
rect 14330 10848 14394 10852
rect 14410 10908 14474 10912
rect 14410 10852 14414 10908
rect 14414 10852 14470 10908
rect 14470 10852 14474 10908
rect 14410 10848 14474 10852
rect 14490 10908 14554 10912
rect 14490 10852 14494 10908
rect 14494 10852 14550 10908
rect 14550 10852 14554 10908
rect 14490 10848 14554 10852
rect 14570 10908 14634 10912
rect 14570 10852 14574 10908
rect 14574 10852 14630 10908
rect 14630 10852 14634 10908
rect 14570 10848 14634 10852
rect 17430 10908 17494 10912
rect 17430 10852 17434 10908
rect 17434 10852 17490 10908
rect 17490 10852 17494 10908
rect 17430 10848 17494 10852
rect 17510 10908 17574 10912
rect 17510 10852 17514 10908
rect 17514 10852 17570 10908
rect 17570 10852 17574 10908
rect 17510 10848 17574 10852
rect 17590 10908 17654 10912
rect 17590 10852 17594 10908
rect 17594 10852 17650 10908
rect 17650 10852 17654 10908
rect 17590 10848 17654 10852
rect 17670 10908 17734 10912
rect 17670 10852 17674 10908
rect 17674 10852 17730 10908
rect 17730 10852 17734 10908
rect 17670 10848 17734 10852
rect 3480 10364 3544 10368
rect 3480 10308 3484 10364
rect 3484 10308 3540 10364
rect 3540 10308 3544 10364
rect 3480 10304 3544 10308
rect 3560 10364 3624 10368
rect 3560 10308 3564 10364
rect 3564 10308 3620 10364
rect 3620 10308 3624 10364
rect 3560 10304 3624 10308
rect 3640 10364 3704 10368
rect 3640 10308 3644 10364
rect 3644 10308 3700 10364
rect 3700 10308 3704 10364
rect 3640 10304 3704 10308
rect 3720 10364 3784 10368
rect 3720 10308 3724 10364
rect 3724 10308 3780 10364
rect 3780 10308 3784 10364
rect 3720 10304 3784 10308
rect 6580 10364 6644 10368
rect 6580 10308 6584 10364
rect 6584 10308 6640 10364
rect 6640 10308 6644 10364
rect 6580 10304 6644 10308
rect 6660 10364 6724 10368
rect 6660 10308 6664 10364
rect 6664 10308 6720 10364
rect 6720 10308 6724 10364
rect 6660 10304 6724 10308
rect 6740 10364 6804 10368
rect 6740 10308 6744 10364
rect 6744 10308 6800 10364
rect 6800 10308 6804 10364
rect 6740 10304 6804 10308
rect 6820 10364 6884 10368
rect 6820 10308 6824 10364
rect 6824 10308 6880 10364
rect 6880 10308 6884 10364
rect 6820 10304 6884 10308
rect 9680 10364 9744 10368
rect 9680 10308 9684 10364
rect 9684 10308 9740 10364
rect 9740 10308 9744 10364
rect 9680 10304 9744 10308
rect 9760 10364 9824 10368
rect 9760 10308 9764 10364
rect 9764 10308 9820 10364
rect 9820 10308 9824 10364
rect 9760 10304 9824 10308
rect 9840 10364 9904 10368
rect 9840 10308 9844 10364
rect 9844 10308 9900 10364
rect 9900 10308 9904 10364
rect 9840 10304 9904 10308
rect 9920 10364 9984 10368
rect 9920 10308 9924 10364
rect 9924 10308 9980 10364
rect 9980 10308 9984 10364
rect 9920 10304 9984 10308
rect 12780 10364 12844 10368
rect 12780 10308 12784 10364
rect 12784 10308 12840 10364
rect 12840 10308 12844 10364
rect 12780 10304 12844 10308
rect 12860 10364 12924 10368
rect 12860 10308 12864 10364
rect 12864 10308 12920 10364
rect 12920 10308 12924 10364
rect 12860 10304 12924 10308
rect 12940 10364 13004 10368
rect 12940 10308 12944 10364
rect 12944 10308 13000 10364
rect 13000 10308 13004 10364
rect 12940 10304 13004 10308
rect 13020 10364 13084 10368
rect 13020 10308 13024 10364
rect 13024 10308 13080 10364
rect 13080 10308 13084 10364
rect 13020 10304 13084 10308
rect 15880 10364 15944 10368
rect 15880 10308 15884 10364
rect 15884 10308 15940 10364
rect 15940 10308 15944 10364
rect 15880 10304 15944 10308
rect 15960 10364 16024 10368
rect 15960 10308 15964 10364
rect 15964 10308 16020 10364
rect 16020 10308 16024 10364
rect 15960 10304 16024 10308
rect 16040 10364 16104 10368
rect 16040 10308 16044 10364
rect 16044 10308 16100 10364
rect 16100 10308 16104 10364
rect 16040 10304 16104 10308
rect 16120 10364 16184 10368
rect 16120 10308 16124 10364
rect 16124 10308 16180 10364
rect 16180 10308 16184 10364
rect 16120 10304 16184 10308
rect 5030 9820 5094 9824
rect 5030 9764 5034 9820
rect 5034 9764 5090 9820
rect 5090 9764 5094 9820
rect 5030 9760 5094 9764
rect 5110 9820 5174 9824
rect 5110 9764 5114 9820
rect 5114 9764 5170 9820
rect 5170 9764 5174 9820
rect 5110 9760 5174 9764
rect 5190 9820 5254 9824
rect 5190 9764 5194 9820
rect 5194 9764 5250 9820
rect 5250 9764 5254 9820
rect 5190 9760 5254 9764
rect 5270 9820 5334 9824
rect 5270 9764 5274 9820
rect 5274 9764 5330 9820
rect 5330 9764 5334 9820
rect 5270 9760 5334 9764
rect 8130 9820 8194 9824
rect 8130 9764 8134 9820
rect 8134 9764 8190 9820
rect 8190 9764 8194 9820
rect 8130 9760 8194 9764
rect 8210 9820 8274 9824
rect 8210 9764 8214 9820
rect 8214 9764 8270 9820
rect 8270 9764 8274 9820
rect 8210 9760 8274 9764
rect 8290 9820 8354 9824
rect 8290 9764 8294 9820
rect 8294 9764 8350 9820
rect 8350 9764 8354 9820
rect 8290 9760 8354 9764
rect 8370 9820 8434 9824
rect 8370 9764 8374 9820
rect 8374 9764 8430 9820
rect 8430 9764 8434 9820
rect 8370 9760 8434 9764
rect 11230 9820 11294 9824
rect 11230 9764 11234 9820
rect 11234 9764 11290 9820
rect 11290 9764 11294 9820
rect 11230 9760 11294 9764
rect 11310 9820 11374 9824
rect 11310 9764 11314 9820
rect 11314 9764 11370 9820
rect 11370 9764 11374 9820
rect 11310 9760 11374 9764
rect 11390 9820 11454 9824
rect 11390 9764 11394 9820
rect 11394 9764 11450 9820
rect 11450 9764 11454 9820
rect 11390 9760 11454 9764
rect 11470 9820 11534 9824
rect 11470 9764 11474 9820
rect 11474 9764 11530 9820
rect 11530 9764 11534 9820
rect 11470 9760 11534 9764
rect 14330 9820 14394 9824
rect 14330 9764 14334 9820
rect 14334 9764 14390 9820
rect 14390 9764 14394 9820
rect 14330 9760 14394 9764
rect 14410 9820 14474 9824
rect 14410 9764 14414 9820
rect 14414 9764 14470 9820
rect 14470 9764 14474 9820
rect 14410 9760 14474 9764
rect 14490 9820 14554 9824
rect 14490 9764 14494 9820
rect 14494 9764 14550 9820
rect 14550 9764 14554 9820
rect 14490 9760 14554 9764
rect 14570 9820 14634 9824
rect 14570 9764 14574 9820
rect 14574 9764 14630 9820
rect 14630 9764 14634 9820
rect 14570 9760 14634 9764
rect 17430 9820 17494 9824
rect 17430 9764 17434 9820
rect 17434 9764 17490 9820
rect 17490 9764 17494 9820
rect 17430 9760 17494 9764
rect 17510 9820 17574 9824
rect 17510 9764 17514 9820
rect 17514 9764 17570 9820
rect 17570 9764 17574 9820
rect 17510 9760 17574 9764
rect 17590 9820 17654 9824
rect 17590 9764 17594 9820
rect 17594 9764 17650 9820
rect 17650 9764 17654 9820
rect 17590 9760 17654 9764
rect 17670 9820 17734 9824
rect 17670 9764 17674 9820
rect 17674 9764 17730 9820
rect 17730 9764 17734 9820
rect 17670 9760 17734 9764
rect 3480 9276 3544 9280
rect 3480 9220 3484 9276
rect 3484 9220 3540 9276
rect 3540 9220 3544 9276
rect 3480 9216 3544 9220
rect 3560 9276 3624 9280
rect 3560 9220 3564 9276
rect 3564 9220 3620 9276
rect 3620 9220 3624 9276
rect 3560 9216 3624 9220
rect 3640 9276 3704 9280
rect 3640 9220 3644 9276
rect 3644 9220 3700 9276
rect 3700 9220 3704 9276
rect 3640 9216 3704 9220
rect 3720 9276 3784 9280
rect 3720 9220 3724 9276
rect 3724 9220 3780 9276
rect 3780 9220 3784 9276
rect 3720 9216 3784 9220
rect 6580 9276 6644 9280
rect 6580 9220 6584 9276
rect 6584 9220 6640 9276
rect 6640 9220 6644 9276
rect 6580 9216 6644 9220
rect 6660 9276 6724 9280
rect 6660 9220 6664 9276
rect 6664 9220 6720 9276
rect 6720 9220 6724 9276
rect 6660 9216 6724 9220
rect 6740 9276 6804 9280
rect 6740 9220 6744 9276
rect 6744 9220 6800 9276
rect 6800 9220 6804 9276
rect 6740 9216 6804 9220
rect 6820 9276 6884 9280
rect 6820 9220 6824 9276
rect 6824 9220 6880 9276
rect 6880 9220 6884 9276
rect 6820 9216 6884 9220
rect 9680 9276 9744 9280
rect 9680 9220 9684 9276
rect 9684 9220 9740 9276
rect 9740 9220 9744 9276
rect 9680 9216 9744 9220
rect 9760 9276 9824 9280
rect 9760 9220 9764 9276
rect 9764 9220 9820 9276
rect 9820 9220 9824 9276
rect 9760 9216 9824 9220
rect 9840 9276 9904 9280
rect 9840 9220 9844 9276
rect 9844 9220 9900 9276
rect 9900 9220 9904 9276
rect 9840 9216 9904 9220
rect 9920 9276 9984 9280
rect 9920 9220 9924 9276
rect 9924 9220 9980 9276
rect 9980 9220 9984 9276
rect 9920 9216 9984 9220
rect 12780 9276 12844 9280
rect 12780 9220 12784 9276
rect 12784 9220 12840 9276
rect 12840 9220 12844 9276
rect 12780 9216 12844 9220
rect 12860 9276 12924 9280
rect 12860 9220 12864 9276
rect 12864 9220 12920 9276
rect 12920 9220 12924 9276
rect 12860 9216 12924 9220
rect 12940 9276 13004 9280
rect 12940 9220 12944 9276
rect 12944 9220 13000 9276
rect 13000 9220 13004 9276
rect 12940 9216 13004 9220
rect 13020 9276 13084 9280
rect 13020 9220 13024 9276
rect 13024 9220 13080 9276
rect 13080 9220 13084 9276
rect 13020 9216 13084 9220
rect 15880 9276 15944 9280
rect 15880 9220 15884 9276
rect 15884 9220 15940 9276
rect 15940 9220 15944 9276
rect 15880 9216 15944 9220
rect 15960 9276 16024 9280
rect 15960 9220 15964 9276
rect 15964 9220 16020 9276
rect 16020 9220 16024 9276
rect 15960 9216 16024 9220
rect 16040 9276 16104 9280
rect 16040 9220 16044 9276
rect 16044 9220 16100 9276
rect 16100 9220 16104 9276
rect 16040 9216 16104 9220
rect 16120 9276 16184 9280
rect 16120 9220 16124 9276
rect 16124 9220 16180 9276
rect 16180 9220 16184 9276
rect 16120 9216 16184 9220
rect 5030 8732 5094 8736
rect 5030 8676 5034 8732
rect 5034 8676 5090 8732
rect 5090 8676 5094 8732
rect 5030 8672 5094 8676
rect 5110 8732 5174 8736
rect 5110 8676 5114 8732
rect 5114 8676 5170 8732
rect 5170 8676 5174 8732
rect 5110 8672 5174 8676
rect 5190 8732 5254 8736
rect 5190 8676 5194 8732
rect 5194 8676 5250 8732
rect 5250 8676 5254 8732
rect 5190 8672 5254 8676
rect 5270 8732 5334 8736
rect 5270 8676 5274 8732
rect 5274 8676 5330 8732
rect 5330 8676 5334 8732
rect 5270 8672 5334 8676
rect 8130 8732 8194 8736
rect 8130 8676 8134 8732
rect 8134 8676 8190 8732
rect 8190 8676 8194 8732
rect 8130 8672 8194 8676
rect 8210 8732 8274 8736
rect 8210 8676 8214 8732
rect 8214 8676 8270 8732
rect 8270 8676 8274 8732
rect 8210 8672 8274 8676
rect 8290 8732 8354 8736
rect 8290 8676 8294 8732
rect 8294 8676 8350 8732
rect 8350 8676 8354 8732
rect 8290 8672 8354 8676
rect 8370 8732 8434 8736
rect 8370 8676 8374 8732
rect 8374 8676 8430 8732
rect 8430 8676 8434 8732
rect 8370 8672 8434 8676
rect 11230 8732 11294 8736
rect 11230 8676 11234 8732
rect 11234 8676 11290 8732
rect 11290 8676 11294 8732
rect 11230 8672 11294 8676
rect 11310 8732 11374 8736
rect 11310 8676 11314 8732
rect 11314 8676 11370 8732
rect 11370 8676 11374 8732
rect 11310 8672 11374 8676
rect 11390 8732 11454 8736
rect 11390 8676 11394 8732
rect 11394 8676 11450 8732
rect 11450 8676 11454 8732
rect 11390 8672 11454 8676
rect 11470 8732 11534 8736
rect 11470 8676 11474 8732
rect 11474 8676 11530 8732
rect 11530 8676 11534 8732
rect 11470 8672 11534 8676
rect 14330 8732 14394 8736
rect 14330 8676 14334 8732
rect 14334 8676 14390 8732
rect 14390 8676 14394 8732
rect 14330 8672 14394 8676
rect 14410 8732 14474 8736
rect 14410 8676 14414 8732
rect 14414 8676 14470 8732
rect 14470 8676 14474 8732
rect 14410 8672 14474 8676
rect 14490 8732 14554 8736
rect 14490 8676 14494 8732
rect 14494 8676 14550 8732
rect 14550 8676 14554 8732
rect 14490 8672 14554 8676
rect 14570 8732 14634 8736
rect 14570 8676 14574 8732
rect 14574 8676 14630 8732
rect 14630 8676 14634 8732
rect 14570 8672 14634 8676
rect 17430 8732 17494 8736
rect 17430 8676 17434 8732
rect 17434 8676 17490 8732
rect 17490 8676 17494 8732
rect 17430 8672 17494 8676
rect 17510 8732 17574 8736
rect 17510 8676 17514 8732
rect 17514 8676 17570 8732
rect 17570 8676 17574 8732
rect 17510 8672 17574 8676
rect 17590 8732 17654 8736
rect 17590 8676 17594 8732
rect 17594 8676 17650 8732
rect 17650 8676 17654 8732
rect 17590 8672 17654 8676
rect 17670 8732 17734 8736
rect 17670 8676 17674 8732
rect 17674 8676 17730 8732
rect 17730 8676 17734 8732
rect 17670 8672 17734 8676
rect 3480 8188 3544 8192
rect 3480 8132 3484 8188
rect 3484 8132 3540 8188
rect 3540 8132 3544 8188
rect 3480 8128 3544 8132
rect 3560 8188 3624 8192
rect 3560 8132 3564 8188
rect 3564 8132 3620 8188
rect 3620 8132 3624 8188
rect 3560 8128 3624 8132
rect 3640 8188 3704 8192
rect 3640 8132 3644 8188
rect 3644 8132 3700 8188
rect 3700 8132 3704 8188
rect 3640 8128 3704 8132
rect 3720 8188 3784 8192
rect 3720 8132 3724 8188
rect 3724 8132 3780 8188
rect 3780 8132 3784 8188
rect 3720 8128 3784 8132
rect 6580 8188 6644 8192
rect 6580 8132 6584 8188
rect 6584 8132 6640 8188
rect 6640 8132 6644 8188
rect 6580 8128 6644 8132
rect 6660 8188 6724 8192
rect 6660 8132 6664 8188
rect 6664 8132 6720 8188
rect 6720 8132 6724 8188
rect 6660 8128 6724 8132
rect 6740 8188 6804 8192
rect 6740 8132 6744 8188
rect 6744 8132 6800 8188
rect 6800 8132 6804 8188
rect 6740 8128 6804 8132
rect 6820 8188 6884 8192
rect 6820 8132 6824 8188
rect 6824 8132 6880 8188
rect 6880 8132 6884 8188
rect 6820 8128 6884 8132
rect 9680 8188 9744 8192
rect 9680 8132 9684 8188
rect 9684 8132 9740 8188
rect 9740 8132 9744 8188
rect 9680 8128 9744 8132
rect 9760 8188 9824 8192
rect 9760 8132 9764 8188
rect 9764 8132 9820 8188
rect 9820 8132 9824 8188
rect 9760 8128 9824 8132
rect 9840 8188 9904 8192
rect 9840 8132 9844 8188
rect 9844 8132 9900 8188
rect 9900 8132 9904 8188
rect 9840 8128 9904 8132
rect 9920 8188 9984 8192
rect 9920 8132 9924 8188
rect 9924 8132 9980 8188
rect 9980 8132 9984 8188
rect 9920 8128 9984 8132
rect 12780 8188 12844 8192
rect 12780 8132 12784 8188
rect 12784 8132 12840 8188
rect 12840 8132 12844 8188
rect 12780 8128 12844 8132
rect 12860 8188 12924 8192
rect 12860 8132 12864 8188
rect 12864 8132 12920 8188
rect 12920 8132 12924 8188
rect 12860 8128 12924 8132
rect 12940 8188 13004 8192
rect 12940 8132 12944 8188
rect 12944 8132 13000 8188
rect 13000 8132 13004 8188
rect 12940 8128 13004 8132
rect 13020 8188 13084 8192
rect 13020 8132 13024 8188
rect 13024 8132 13080 8188
rect 13080 8132 13084 8188
rect 13020 8128 13084 8132
rect 15880 8188 15944 8192
rect 15880 8132 15884 8188
rect 15884 8132 15940 8188
rect 15940 8132 15944 8188
rect 15880 8128 15944 8132
rect 15960 8188 16024 8192
rect 15960 8132 15964 8188
rect 15964 8132 16020 8188
rect 16020 8132 16024 8188
rect 15960 8128 16024 8132
rect 16040 8188 16104 8192
rect 16040 8132 16044 8188
rect 16044 8132 16100 8188
rect 16100 8132 16104 8188
rect 16040 8128 16104 8132
rect 16120 8188 16184 8192
rect 16120 8132 16124 8188
rect 16124 8132 16180 8188
rect 16180 8132 16184 8188
rect 16120 8128 16184 8132
rect 5030 7644 5094 7648
rect 5030 7588 5034 7644
rect 5034 7588 5090 7644
rect 5090 7588 5094 7644
rect 5030 7584 5094 7588
rect 5110 7644 5174 7648
rect 5110 7588 5114 7644
rect 5114 7588 5170 7644
rect 5170 7588 5174 7644
rect 5110 7584 5174 7588
rect 5190 7644 5254 7648
rect 5190 7588 5194 7644
rect 5194 7588 5250 7644
rect 5250 7588 5254 7644
rect 5190 7584 5254 7588
rect 5270 7644 5334 7648
rect 5270 7588 5274 7644
rect 5274 7588 5330 7644
rect 5330 7588 5334 7644
rect 5270 7584 5334 7588
rect 8130 7644 8194 7648
rect 8130 7588 8134 7644
rect 8134 7588 8190 7644
rect 8190 7588 8194 7644
rect 8130 7584 8194 7588
rect 8210 7644 8274 7648
rect 8210 7588 8214 7644
rect 8214 7588 8270 7644
rect 8270 7588 8274 7644
rect 8210 7584 8274 7588
rect 8290 7644 8354 7648
rect 8290 7588 8294 7644
rect 8294 7588 8350 7644
rect 8350 7588 8354 7644
rect 8290 7584 8354 7588
rect 8370 7644 8434 7648
rect 8370 7588 8374 7644
rect 8374 7588 8430 7644
rect 8430 7588 8434 7644
rect 8370 7584 8434 7588
rect 11230 7644 11294 7648
rect 11230 7588 11234 7644
rect 11234 7588 11290 7644
rect 11290 7588 11294 7644
rect 11230 7584 11294 7588
rect 11310 7644 11374 7648
rect 11310 7588 11314 7644
rect 11314 7588 11370 7644
rect 11370 7588 11374 7644
rect 11310 7584 11374 7588
rect 11390 7644 11454 7648
rect 11390 7588 11394 7644
rect 11394 7588 11450 7644
rect 11450 7588 11454 7644
rect 11390 7584 11454 7588
rect 11470 7644 11534 7648
rect 11470 7588 11474 7644
rect 11474 7588 11530 7644
rect 11530 7588 11534 7644
rect 11470 7584 11534 7588
rect 14330 7644 14394 7648
rect 14330 7588 14334 7644
rect 14334 7588 14390 7644
rect 14390 7588 14394 7644
rect 14330 7584 14394 7588
rect 14410 7644 14474 7648
rect 14410 7588 14414 7644
rect 14414 7588 14470 7644
rect 14470 7588 14474 7644
rect 14410 7584 14474 7588
rect 14490 7644 14554 7648
rect 14490 7588 14494 7644
rect 14494 7588 14550 7644
rect 14550 7588 14554 7644
rect 14490 7584 14554 7588
rect 14570 7644 14634 7648
rect 14570 7588 14574 7644
rect 14574 7588 14630 7644
rect 14630 7588 14634 7644
rect 14570 7584 14634 7588
rect 17430 7644 17494 7648
rect 17430 7588 17434 7644
rect 17434 7588 17490 7644
rect 17490 7588 17494 7644
rect 17430 7584 17494 7588
rect 17510 7644 17574 7648
rect 17510 7588 17514 7644
rect 17514 7588 17570 7644
rect 17570 7588 17574 7644
rect 17510 7584 17574 7588
rect 17590 7644 17654 7648
rect 17590 7588 17594 7644
rect 17594 7588 17650 7644
rect 17650 7588 17654 7644
rect 17590 7584 17654 7588
rect 17670 7644 17734 7648
rect 17670 7588 17674 7644
rect 17674 7588 17730 7644
rect 17730 7588 17734 7644
rect 17670 7584 17734 7588
rect 3480 7100 3544 7104
rect 3480 7044 3484 7100
rect 3484 7044 3540 7100
rect 3540 7044 3544 7100
rect 3480 7040 3544 7044
rect 3560 7100 3624 7104
rect 3560 7044 3564 7100
rect 3564 7044 3620 7100
rect 3620 7044 3624 7100
rect 3560 7040 3624 7044
rect 3640 7100 3704 7104
rect 3640 7044 3644 7100
rect 3644 7044 3700 7100
rect 3700 7044 3704 7100
rect 3640 7040 3704 7044
rect 3720 7100 3784 7104
rect 3720 7044 3724 7100
rect 3724 7044 3780 7100
rect 3780 7044 3784 7100
rect 3720 7040 3784 7044
rect 6580 7100 6644 7104
rect 6580 7044 6584 7100
rect 6584 7044 6640 7100
rect 6640 7044 6644 7100
rect 6580 7040 6644 7044
rect 6660 7100 6724 7104
rect 6660 7044 6664 7100
rect 6664 7044 6720 7100
rect 6720 7044 6724 7100
rect 6660 7040 6724 7044
rect 6740 7100 6804 7104
rect 6740 7044 6744 7100
rect 6744 7044 6800 7100
rect 6800 7044 6804 7100
rect 6740 7040 6804 7044
rect 6820 7100 6884 7104
rect 6820 7044 6824 7100
rect 6824 7044 6880 7100
rect 6880 7044 6884 7100
rect 6820 7040 6884 7044
rect 9680 7100 9744 7104
rect 9680 7044 9684 7100
rect 9684 7044 9740 7100
rect 9740 7044 9744 7100
rect 9680 7040 9744 7044
rect 9760 7100 9824 7104
rect 9760 7044 9764 7100
rect 9764 7044 9820 7100
rect 9820 7044 9824 7100
rect 9760 7040 9824 7044
rect 9840 7100 9904 7104
rect 9840 7044 9844 7100
rect 9844 7044 9900 7100
rect 9900 7044 9904 7100
rect 9840 7040 9904 7044
rect 9920 7100 9984 7104
rect 9920 7044 9924 7100
rect 9924 7044 9980 7100
rect 9980 7044 9984 7100
rect 9920 7040 9984 7044
rect 12780 7100 12844 7104
rect 12780 7044 12784 7100
rect 12784 7044 12840 7100
rect 12840 7044 12844 7100
rect 12780 7040 12844 7044
rect 12860 7100 12924 7104
rect 12860 7044 12864 7100
rect 12864 7044 12920 7100
rect 12920 7044 12924 7100
rect 12860 7040 12924 7044
rect 12940 7100 13004 7104
rect 12940 7044 12944 7100
rect 12944 7044 13000 7100
rect 13000 7044 13004 7100
rect 12940 7040 13004 7044
rect 13020 7100 13084 7104
rect 13020 7044 13024 7100
rect 13024 7044 13080 7100
rect 13080 7044 13084 7100
rect 13020 7040 13084 7044
rect 15880 7100 15944 7104
rect 15880 7044 15884 7100
rect 15884 7044 15940 7100
rect 15940 7044 15944 7100
rect 15880 7040 15944 7044
rect 15960 7100 16024 7104
rect 15960 7044 15964 7100
rect 15964 7044 16020 7100
rect 16020 7044 16024 7100
rect 15960 7040 16024 7044
rect 16040 7100 16104 7104
rect 16040 7044 16044 7100
rect 16044 7044 16100 7100
rect 16100 7044 16104 7100
rect 16040 7040 16104 7044
rect 16120 7100 16184 7104
rect 16120 7044 16124 7100
rect 16124 7044 16180 7100
rect 16180 7044 16184 7100
rect 16120 7040 16184 7044
rect 5030 6556 5094 6560
rect 5030 6500 5034 6556
rect 5034 6500 5090 6556
rect 5090 6500 5094 6556
rect 5030 6496 5094 6500
rect 5110 6556 5174 6560
rect 5110 6500 5114 6556
rect 5114 6500 5170 6556
rect 5170 6500 5174 6556
rect 5110 6496 5174 6500
rect 5190 6556 5254 6560
rect 5190 6500 5194 6556
rect 5194 6500 5250 6556
rect 5250 6500 5254 6556
rect 5190 6496 5254 6500
rect 5270 6556 5334 6560
rect 5270 6500 5274 6556
rect 5274 6500 5330 6556
rect 5330 6500 5334 6556
rect 5270 6496 5334 6500
rect 8130 6556 8194 6560
rect 8130 6500 8134 6556
rect 8134 6500 8190 6556
rect 8190 6500 8194 6556
rect 8130 6496 8194 6500
rect 8210 6556 8274 6560
rect 8210 6500 8214 6556
rect 8214 6500 8270 6556
rect 8270 6500 8274 6556
rect 8210 6496 8274 6500
rect 8290 6556 8354 6560
rect 8290 6500 8294 6556
rect 8294 6500 8350 6556
rect 8350 6500 8354 6556
rect 8290 6496 8354 6500
rect 8370 6556 8434 6560
rect 8370 6500 8374 6556
rect 8374 6500 8430 6556
rect 8430 6500 8434 6556
rect 8370 6496 8434 6500
rect 11230 6556 11294 6560
rect 11230 6500 11234 6556
rect 11234 6500 11290 6556
rect 11290 6500 11294 6556
rect 11230 6496 11294 6500
rect 11310 6556 11374 6560
rect 11310 6500 11314 6556
rect 11314 6500 11370 6556
rect 11370 6500 11374 6556
rect 11310 6496 11374 6500
rect 11390 6556 11454 6560
rect 11390 6500 11394 6556
rect 11394 6500 11450 6556
rect 11450 6500 11454 6556
rect 11390 6496 11454 6500
rect 11470 6556 11534 6560
rect 11470 6500 11474 6556
rect 11474 6500 11530 6556
rect 11530 6500 11534 6556
rect 11470 6496 11534 6500
rect 14330 6556 14394 6560
rect 14330 6500 14334 6556
rect 14334 6500 14390 6556
rect 14390 6500 14394 6556
rect 14330 6496 14394 6500
rect 14410 6556 14474 6560
rect 14410 6500 14414 6556
rect 14414 6500 14470 6556
rect 14470 6500 14474 6556
rect 14410 6496 14474 6500
rect 14490 6556 14554 6560
rect 14490 6500 14494 6556
rect 14494 6500 14550 6556
rect 14550 6500 14554 6556
rect 14490 6496 14554 6500
rect 14570 6556 14634 6560
rect 14570 6500 14574 6556
rect 14574 6500 14630 6556
rect 14630 6500 14634 6556
rect 14570 6496 14634 6500
rect 17430 6556 17494 6560
rect 17430 6500 17434 6556
rect 17434 6500 17490 6556
rect 17490 6500 17494 6556
rect 17430 6496 17494 6500
rect 17510 6556 17574 6560
rect 17510 6500 17514 6556
rect 17514 6500 17570 6556
rect 17570 6500 17574 6556
rect 17510 6496 17574 6500
rect 17590 6556 17654 6560
rect 17590 6500 17594 6556
rect 17594 6500 17650 6556
rect 17650 6500 17654 6556
rect 17590 6496 17654 6500
rect 17670 6556 17734 6560
rect 17670 6500 17674 6556
rect 17674 6500 17730 6556
rect 17730 6500 17734 6556
rect 17670 6496 17734 6500
rect 3480 6012 3544 6016
rect 3480 5956 3484 6012
rect 3484 5956 3540 6012
rect 3540 5956 3544 6012
rect 3480 5952 3544 5956
rect 3560 6012 3624 6016
rect 3560 5956 3564 6012
rect 3564 5956 3620 6012
rect 3620 5956 3624 6012
rect 3560 5952 3624 5956
rect 3640 6012 3704 6016
rect 3640 5956 3644 6012
rect 3644 5956 3700 6012
rect 3700 5956 3704 6012
rect 3640 5952 3704 5956
rect 3720 6012 3784 6016
rect 3720 5956 3724 6012
rect 3724 5956 3780 6012
rect 3780 5956 3784 6012
rect 3720 5952 3784 5956
rect 6580 6012 6644 6016
rect 6580 5956 6584 6012
rect 6584 5956 6640 6012
rect 6640 5956 6644 6012
rect 6580 5952 6644 5956
rect 6660 6012 6724 6016
rect 6660 5956 6664 6012
rect 6664 5956 6720 6012
rect 6720 5956 6724 6012
rect 6660 5952 6724 5956
rect 6740 6012 6804 6016
rect 6740 5956 6744 6012
rect 6744 5956 6800 6012
rect 6800 5956 6804 6012
rect 6740 5952 6804 5956
rect 6820 6012 6884 6016
rect 6820 5956 6824 6012
rect 6824 5956 6880 6012
rect 6880 5956 6884 6012
rect 6820 5952 6884 5956
rect 9680 6012 9744 6016
rect 9680 5956 9684 6012
rect 9684 5956 9740 6012
rect 9740 5956 9744 6012
rect 9680 5952 9744 5956
rect 9760 6012 9824 6016
rect 9760 5956 9764 6012
rect 9764 5956 9820 6012
rect 9820 5956 9824 6012
rect 9760 5952 9824 5956
rect 9840 6012 9904 6016
rect 9840 5956 9844 6012
rect 9844 5956 9900 6012
rect 9900 5956 9904 6012
rect 9840 5952 9904 5956
rect 9920 6012 9984 6016
rect 9920 5956 9924 6012
rect 9924 5956 9980 6012
rect 9980 5956 9984 6012
rect 9920 5952 9984 5956
rect 12780 6012 12844 6016
rect 12780 5956 12784 6012
rect 12784 5956 12840 6012
rect 12840 5956 12844 6012
rect 12780 5952 12844 5956
rect 12860 6012 12924 6016
rect 12860 5956 12864 6012
rect 12864 5956 12920 6012
rect 12920 5956 12924 6012
rect 12860 5952 12924 5956
rect 12940 6012 13004 6016
rect 12940 5956 12944 6012
rect 12944 5956 13000 6012
rect 13000 5956 13004 6012
rect 12940 5952 13004 5956
rect 13020 6012 13084 6016
rect 13020 5956 13024 6012
rect 13024 5956 13080 6012
rect 13080 5956 13084 6012
rect 13020 5952 13084 5956
rect 15880 6012 15944 6016
rect 15880 5956 15884 6012
rect 15884 5956 15940 6012
rect 15940 5956 15944 6012
rect 15880 5952 15944 5956
rect 15960 6012 16024 6016
rect 15960 5956 15964 6012
rect 15964 5956 16020 6012
rect 16020 5956 16024 6012
rect 15960 5952 16024 5956
rect 16040 6012 16104 6016
rect 16040 5956 16044 6012
rect 16044 5956 16100 6012
rect 16100 5956 16104 6012
rect 16040 5952 16104 5956
rect 16120 6012 16184 6016
rect 16120 5956 16124 6012
rect 16124 5956 16180 6012
rect 16180 5956 16184 6012
rect 16120 5952 16184 5956
rect 5030 5468 5094 5472
rect 5030 5412 5034 5468
rect 5034 5412 5090 5468
rect 5090 5412 5094 5468
rect 5030 5408 5094 5412
rect 5110 5468 5174 5472
rect 5110 5412 5114 5468
rect 5114 5412 5170 5468
rect 5170 5412 5174 5468
rect 5110 5408 5174 5412
rect 5190 5468 5254 5472
rect 5190 5412 5194 5468
rect 5194 5412 5250 5468
rect 5250 5412 5254 5468
rect 5190 5408 5254 5412
rect 5270 5468 5334 5472
rect 5270 5412 5274 5468
rect 5274 5412 5330 5468
rect 5330 5412 5334 5468
rect 5270 5408 5334 5412
rect 8130 5468 8194 5472
rect 8130 5412 8134 5468
rect 8134 5412 8190 5468
rect 8190 5412 8194 5468
rect 8130 5408 8194 5412
rect 8210 5468 8274 5472
rect 8210 5412 8214 5468
rect 8214 5412 8270 5468
rect 8270 5412 8274 5468
rect 8210 5408 8274 5412
rect 8290 5468 8354 5472
rect 8290 5412 8294 5468
rect 8294 5412 8350 5468
rect 8350 5412 8354 5468
rect 8290 5408 8354 5412
rect 8370 5468 8434 5472
rect 8370 5412 8374 5468
rect 8374 5412 8430 5468
rect 8430 5412 8434 5468
rect 8370 5408 8434 5412
rect 11230 5468 11294 5472
rect 11230 5412 11234 5468
rect 11234 5412 11290 5468
rect 11290 5412 11294 5468
rect 11230 5408 11294 5412
rect 11310 5468 11374 5472
rect 11310 5412 11314 5468
rect 11314 5412 11370 5468
rect 11370 5412 11374 5468
rect 11310 5408 11374 5412
rect 11390 5468 11454 5472
rect 11390 5412 11394 5468
rect 11394 5412 11450 5468
rect 11450 5412 11454 5468
rect 11390 5408 11454 5412
rect 11470 5468 11534 5472
rect 11470 5412 11474 5468
rect 11474 5412 11530 5468
rect 11530 5412 11534 5468
rect 11470 5408 11534 5412
rect 14330 5468 14394 5472
rect 14330 5412 14334 5468
rect 14334 5412 14390 5468
rect 14390 5412 14394 5468
rect 14330 5408 14394 5412
rect 14410 5468 14474 5472
rect 14410 5412 14414 5468
rect 14414 5412 14470 5468
rect 14470 5412 14474 5468
rect 14410 5408 14474 5412
rect 14490 5468 14554 5472
rect 14490 5412 14494 5468
rect 14494 5412 14550 5468
rect 14550 5412 14554 5468
rect 14490 5408 14554 5412
rect 14570 5468 14634 5472
rect 14570 5412 14574 5468
rect 14574 5412 14630 5468
rect 14630 5412 14634 5468
rect 14570 5408 14634 5412
rect 17430 5468 17494 5472
rect 17430 5412 17434 5468
rect 17434 5412 17490 5468
rect 17490 5412 17494 5468
rect 17430 5408 17494 5412
rect 17510 5468 17574 5472
rect 17510 5412 17514 5468
rect 17514 5412 17570 5468
rect 17570 5412 17574 5468
rect 17510 5408 17574 5412
rect 17590 5468 17654 5472
rect 17590 5412 17594 5468
rect 17594 5412 17650 5468
rect 17650 5412 17654 5468
rect 17590 5408 17654 5412
rect 17670 5468 17734 5472
rect 17670 5412 17674 5468
rect 17674 5412 17730 5468
rect 17730 5412 17734 5468
rect 17670 5408 17734 5412
rect 3480 4924 3544 4928
rect 3480 4868 3484 4924
rect 3484 4868 3540 4924
rect 3540 4868 3544 4924
rect 3480 4864 3544 4868
rect 3560 4924 3624 4928
rect 3560 4868 3564 4924
rect 3564 4868 3620 4924
rect 3620 4868 3624 4924
rect 3560 4864 3624 4868
rect 3640 4924 3704 4928
rect 3640 4868 3644 4924
rect 3644 4868 3700 4924
rect 3700 4868 3704 4924
rect 3640 4864 3704 4868
rect 3720 4924 3784 4928
rect 3720 4868 3724 4924
rect 3724 4868 3780 4924
rect 3780 4868 3784 4924
rect 3720 4864 3784 4868
rect 6580 4924 6644 4928
rect 6580 4868 6584 4924
rect 6584 4868 6640 4924
rect 6640 4868 6644 4924
rect 6580 4864 6644 4868
rect 6660 4924 6724 4928
rect 6660 4868 6664 4924
rect 6664 4868 6720 4924
rect 6720 4868 6724 4924
rect 6660 4864 6724 4868
rect 6740 4924 6804 4928
rect 6740 4868 6744 4924
rect 6744 4868 6800 4924
rect 6800 4868 6804 4924
rect 6740 4864 6804 4868
rect 6820 4924 6884 4928
rect 6820 4868 6824 4924
rect 6824 4868 6880 4924
rect 6880 4868 6884 4924
rect 6820 4864 6884 4868
rect 9680 4924 9744 4928
rect 9680 4868 9684 4924
rect 9684 4868 9740 4924
rect 9740 4868 9744 4924
rect 9680 4864 9744 4868
rect 9760 4924 9824 4928
rect 9760 4868 9764 4924
rect 9764 4868 9820 4924
rect 9820 4868 9824 4924
rect 9760 4864 9824 4868
rect 9840 4924 9904 4928
rect 9840 4868 9844 4924
rect 9844 4868 9900 4924
rect 9900 4868 9904 4924
rect 9840 4864 9904 4868
rect 9920 4924 9984 4928
rect 9920 4868 9924 4924
rect 9924 4868 9980 4924
rect 9980 4868 9984 4924
rect 9920 4864 9984 4868
rect 12780 4924 12844 4928
rect 12780 4868 12784 4924
rect 12784 4868 12840 4924
rect 12840 4868 12844 4924
rect 12780 4864 12844 4868
rect 12860 4924 12924 4928
rect 12860 4868 12864 4924
rect 12864 4868 12920 4924
rect 12920 4868 12924 4924
rect 12860 4864 12924 4868
rect 12940 4924 13004 4928
rect 12940 4868 12944 4924
rect 12944 4868 13000 4924
rect 13000 4868 13004 4924
rect 12940 4864 13004 4868
rect 13020 4924 13084 4928
rect 13020 4868 13024 4924
rect 13024 4868 13080 4924
rect 13080 4868 13084 4924
rect 13020 4864 13084 4868
rect 15880 4924 15944 4928
rect 15880 4868 15884 4924
rect 15884 4868 15940 4924
rect 15940 4868 15944 4924
rect 15880 4864 15944 4868
rect 15960 4924 16024 4928
rect 15960 4868 15964 4924
rect 15964 4868 16020 4924
rect 16020 4868 16024 4924
rect 15960 4864 16024 4868
rect 16040 4924 16104 4928
rect 16040 4868 16044 4924
rect 16044 4868 16100 4924
rect 16100 4868 16104 4924
rect 16040 4864 16104 4868
rect 16120 4924 16184 4928
rect 16120 4868 16124 4924
rect 16124 4868 16180 4924
rect 16180 4868 16184 4924
rect 16120 4864 16184 4868
rect 5030 4380 5094 4384
rect 5030 4324 5034 4380
rect 5034 4324 5090 4380
rect 5090 4324 5094 4380
rect 5030 4320 5094 4324
rect 5110 4380 5174 4384
rect 5110 4324 5114 4380
rect 5114 4324 5170 4380
rect 5170 4324 5174 4380
rect 5110 4320 5174 4324
rect 5190 4380 5254 4384
rect 5190 4324 5194 4380
rect 5194 4324 5250 4380
rect 5250 4324 5254 4380
rect 5190 4320 5254 4324
rect 5270 4380 5334 4384
rect 5270 4324 5274 4380
rect 5274 4324 5330 4380
rect 5330 4324 5334 4380
rect 5270 4320 5334 4324
rect 8130 4380 8194 4384
rect 8130 4324 8134 4380
rect 8134 4324 8190 4380
rect 8190 4324 8194 4380
rect 8130 4320 8194 4324
rect 8210 4380 8274 4384
rect 8210 4324 8214 4380
rect 8214 4324 8270 4380
rect 8270 4324 8274 4380
rect 8210 4320 8274 4324
rect 8290 4380 8354 4384
rect 8290 4324 8294 4380
rect 8294 4324 8350 4380
rect 8350 4324 8354 4380
rect 8290 4320 8354 4324
rect 8370 4380 8434 4384
rect 8370 4324 8374 4380
rect 8374 4324 8430 4380
rect 8430 4324 8434 4380
rect 8370 4320 8434 4324
rect 11230 4380 11294 4384
rect 11230 4324 11234 4380
rect 11234 4324 11290 4380
rect 11290 4324 11294 4380
rect 11230 4320 11294 4324
rect 11310 4380 11374 4384
rect 11310 4324 11314 4380
rect 11314 4324 11370 4380
rect 11370 4324 11374 4380
rect 11310 4320 11374 4324
rect 11390 4380 11454 4384
rect 11390 4324 11394 4380
rect 11394 4324 11450 4380
rect 11450 4324 11454 4380
rect 11390 4320 11454 4324
rect 11470 4380 11534 4384
rect 11470 4324 11474 4380
rect 11474 4324 11530 4380
rect 11530 4324 11534 4380
rect 11470 4320 11534 4324
rect 14330 4380 14394 4384
rect 14330 4324 14334 4380
rect 14334 4324 14390 4380
rect 14390 4324 14394 4380
rect 14330 4320 14394 4324
rect 14410 4380 14474 4384
rect 14410 4324 14414 4380
rect 14414 4324 14470 4380
rect 14470 4324 14474 4380
rect 14410 4320 14474 4324
rect 14490 4380 14554 4384
rect 14490 4324 14494 4380
rect 14494 4324 14550 4380
rect 14550 4324 14554 4380
rect 14490 4320 14554 4324
rect 14570 4380 14634 4384
rect 14570 4324 14574 4380
rect 14574 4324 14630 4380
rect 14630 4324 14634 4380
rect 14570 4320 14634 4324
rect 17430 4380 17494 4384
rect 17430 4324 17434 4380
rect 17434 4324 17490 4380
rect 17490 4324 17494 4380
rect 17430 4320 17494 4324
rect 17510 4380 17574 4384
rect 17510 4324 17514 4380
rect 17514 4324 17570 4380
rect 17570 4324 17574 4380
rect 17510 4320 17574 4324
rect 17590 4380 17654 4384
rect 17590 4324 17594 4380
rect 17594 4324 17650 4380
rect 17650 4324 17654 4380
rect 17590 4320 17654 4324
rect 17670 4380 17734 4384
rect 17670 4324 17674 4380
rect 17674 4324 17730 4380
rect 17730 4324 17734 4380
rect 17670 4320 17734 4324
rect 3480 3836 3544 3840
rect 3480 3780 3484 3836
rect 3484 3780 3540 3836
rect 3540 3780 3544 3836
rect 3480 3776 3544 3780
rect 3560 3836 3624 3840
rect 3560 3780 3564 3836
rect 3564 3780 3620 3836
rect 3620 3780 3624 3836
rect 3560 3776 3624 3780
rect 3640 3836 3704 3840
rect 3640 3780 3644 3836
rect 3644 3780 3700 3836
rect 3700 3780 3704 3836
rect 3640 3776 3704 3780
rect 3720 3836 3784 3840
rect 3720 3780 3724 3836
rect 3724 3780 3780 3836
rect 3780 3780 3784 3836
rect 3720 3776 3784 3780
rect 6580 3836 6644 3840
rect 6580 3780 6584 3836
rect 6584 3780 6640 3836
rect 6640 3780 6644 3836
rect 6580 3776 6644 3780
rect 6660 3836 6724 3840
rect 6660 3780 6664 3836
rect 6664 3780 6720 3836
rect 6720 3780 6724 3836
rect 6660 3776 6724 3780
rect 6740 3836 6804 3840
rect 6740 3780 6744 3836
rect 6744 3780 6800 3836
rect 6800 3780 6804 3836
rect 6740 3776 6804 3780
rect 6820 3836 6884 3840
rect 6820 3780 6824 3836
rect 6824 3780 6880 3836
rect 6880 3780 6884 3836
rect 6820 3776 6884 3780
rect 9680 3836 9744 3840
rect 9680 3780 9684 3836
rect 9684 3780 9740 3836
rect 9740 3780 9744 3836
rect 9680 3776 9744 3780
rect 9760 3836 9824 3840
rect 9760 3780 9764 3836
rect 9764 3780 9820 3836
rect 9820 3780 9824 3836
rect 9760 3776 9824 3780
rect 9840 3836 9904 3840
rect 9840 3780 9844 3836
rect 9844 3780 9900 3836
rect 9900 3780 9904 3836
rect 9840 3776 9904 3780
rect 9920 3836 9984 3840
rect 9920 3780 9924 3836
rect 9924 3780 9980 3836
rect 9980 3780 9984 3836
rect 9920 3776 9984 3780
rect 12780 3836 12844 3840
rect 12780 3780 12784 3836
rect 12784 3780 12840 3836
rect 12840 3780 12844 3836
rect 12780 3776 12844 3780
rect 12860 3836 12924 3840
rect 12860 3780 12864 3836
rect 12864 3780 12920 3836
rect 12920 3780 12924 3836
rect 12860 3776 12924 3780
rect 12940 3836 13004 3840
rect 12940 3780 12944 3836
rect 12944 3780 13000 3836
rect 13000 3780 13004 3836
rect 12940 3776 13004 3780
rect 13020 3836 13084 3840
rect 13020 3780 13024 3836
rect 13024 3780 13080 3836
rect 13080 3780 13084 3836
rect 13020 3776 13084 3780
rect 15880 3836 15944 3840
rect 15880 3780 15884 3836
rect 15884 3780 15940 3836
rect 15940 3780 15944 3836
rect 15880 3776 15944 3780
rect 15960 3836 16024 3840
rect 15960 3780 15964 3836
rect 15964 3780 16020 3836
rect 16020 3780 16024 3836
rect 15960 3776 16024 3780
rect 16040 3836 16104 3840
rect 16040 3780 16044 3836
rect 16044 3780 16100 3836
rect 16100 3780 16104 3836
rect 16040 3776 16104 3780
rect 16120 3836 16184 3840
rect 16120 3780 16124 3836
rect 16124 3780 16180 3836
rect 16180 3780 16184 3836
rect 16120 3776 16184 3780
rect 5030 3292 5094 3296
rect 5030 3236 5034 3292
rect 5034 3236 5090 3292
rect 5090 3236 5094 3292
rect 5030 3232 5094 3236
rect 5110 3292 5174 3296
rect 5110 3236 5114 3292
rect 5114 3236 5170 3292
rect 5170 3236 5174 3292
rect 5110 3232 5174 3236
rect 5190 3292 5254 3296
rect 5190 3236 5194 3292
rect 5194 3236 5250 3292
rect 5250 3236 5254 3292
rect 5190 3232 5254 3236
rect 5270 3292 5334 3296
rect 5270 3236 5274 3292
rect 5274 3236 5330 3292
rect 5330 3236 5334 3292
rect 5270 3232 5334 3236
rect 8130 3292 8194 3296
rect 8130 3236 8134 3292
rect 8134 3236 8190 3292
rect 8190 3236 8194 3292
rect 8130 3232 8194 3236
rect 8210 3292 8274 3296
rect 8210 3236 8214 3292
rect 8214 3236 8270 3292
rect 8270 3236 8274 3292
rect 8210 3232 8274 3236
rect 8290 3292 8354 3296
rect 8290 3236 8294 3292
rect 8294 3236 8350 3292
rect 8350 3236 8354 3292
rect 8290 3232 8354 3236
rect 8370 3292 8434 3296
rect 8370 3236 8374 3292
rect 8374 3236 8430 3292
rect 8430 3236 8434 3292
rect 8370 3232 8434 3236
rect 11230 3292 11294 3296
rect 11230 3236 11234 3292
rect 11234 3236 11290 3292
rect 11290 3236 11294 3292
rect 11230 3232 11294 3236
rect 11310 3292 11374 3296
rect 11310 3236 11314 3292
rect 11314 3236 11370 3292
rect 11370 3236 11374 3292
rect 11310 3232 11374 3236
rect 11390 3292 11454 3296
rect 11390 3236 11394 3292
rect 11394 3236 11450 3292
rect 11450 3236 11454 3292
rect 11390 3232 11454 3236
rect 11470 3292 11534 3296
rect 11470 3236 11474 3292
rect 11474 3236 11530 3292
rect 11530 3236 11534 3292
rect 11470 3232 11534 3236
rect 14330 3292 14394 3296
rect 14330 3236 14334 3292
rect 14334 3236 14390 3292
rect 14390 3236 14394 3292
rect 14330 3232 14394 3236
rect 14410 3292 14474 3296
rect 14410 3236 14414 3292
rect 14414 3236 14470 3292
rect 14470 3236 14474 3292
rect 14410 3232 14474 3236
rect 14490 3292 14554 3296
rect 14490 3236 14494 3292
rect 14494 3236 14550 3292
rect 14550 3236 14554 3292
rect 14490 3232 14554 3236
rect 14570 3292 14634 3296
rect 14570 3236 14574 3292
rect 14574 3236 14630 3292
rect 14630 3236 14634 3292
rect 14570 3232 14634 3236
rect 17430 3292 17494 3296
rect 17430 3236 17434 3292
rect 17434 3236 17490 3292
rect 17490 3236 17494 3292
rect 17430 3232 17494 3236
rect 17510 3292 17574 3296
rect 17510 3236 17514 3292
rect 17514 3236 17570 3292
rect 17570 3236 17574 3292
rect 17510 3232 17574 3236
rect 17590 3292 17654 3296
rect 17590 3236 17594 3292
rect 17594 3236 17650 3292
rect 17650 3236 17654 3292
rect 17590 3232 17654 3236
rect 17670 3292 17734 3296
rect 17670 3236 17674 3292
rect 17674 3236 17730 3292
rect 17730 3236 17734 3292
rect 17670 3232 17734 3236
rect 3480 2748 3544 2752
rect 3480 2692 3484 2748
rect 3484 2692 3540 2748
rect 3540 2692 3544 2748
rect 3480 2688 3544 2692
rect 3560 2748 3624 2752
rect 3560 2692 3564 2748
rect 3564 2692 3620 2748
rect 3620 2692 3624 2748
rect 3560 2688 3624 2692
rect 3640 2748 3704 2752
rect 3640 2692 3644 2748
rect 3644 2692 3700 2748
rect 3700 2692 3704 2748
rect 3640 2688 3704 2692
rect 3720 2748 3784 2752
rect 3720 2692 3724 2748
rect 3724 2692 3780 2748
rect 3780 2692 3784 2748
rect 3720 2688 3784 2692
rect 6580 2748 6644 2752
rect 6580 2692 6584 2748
rect 6584 2692 6640 2748
rect 6640 2692 6644 2748
rect 6580 2688 6644 2692
rect 6660 2748 6724 2752
rect 6660 2692 6664 2748
rect 6664 2692 6720 2748
rect 6720 2692 6724 2748
rect 6660 2688 6724 2692
rect 6740 2748 6804 2752
rect 6740 2692 6744 2748
rect 6744 2692 6800 2748
rect 6800 2692 6804 2748
rect 6740 2688 6804 2692
rect 6820 2748 6884 2752
rect 6820 2692 6824 2748
rect 6824 2692 6880 2748
rect 6880 2692 6884 2748
rect 6820 2688 6884 2692
rect 9680 2748 9744 2752
rect 9680 2692 9684 2748
rect 9684 2692 9740 2748
rect 9740 2692 9744 2748
rect 9680 2688 9744 2692
rect 9760 2748 9824 2752
rect 9760 2692 9764 2748
rect 9764 2692 9820 2748
rect 9820 2692 9824 2748
rect 9760 2688 9824 2692
rect 9840 2748 9904 2752
rect 9840 2692 9844 2748
rect 9844 2692 9900 2748
rect 9900 2692 9904 2748
rect 9840 2688 9904 2692
rect 9920 2748 9984 2752
rect 9920 2692 9924 2748
rect 9924 2692 9980 2748
rect 9980 2692 9984 2748
rect 9920 2688 9984 2692
rect 12780 2748 12844 2752
rect 12780 2692 12784 2748
rect 12784 2692 12840 2748
rect 12840 2692 12844 2748
rect 12780 2688 12844 2692
rect 12860 2748 12924 2752
rect 12860 2692 12864 2748
rect 12864 2692 12920 2748
rect 12920 2692 12924 2748
rect 12860 2688 12924 2692
rect 12940 2748 13004 2752
rect 12940 2692 12944 2748
rect 12944 2692 13000 2748
rect 13000 2692 13004 2748
rect 12940 2688 13004 2692
rect 13020 2748 13084 2752
rect 13020 2692 13024 2748
rect 13024 2692 13080 2748
rect 13080 2692 13084 2748
rect 13020 2688 13084 2692
rect 15880 2748 15944 2752
rect 15880 2692 15884 2748
rect 15884 2692 15940 2748
rect 15940 2692 15944 2748
rect 15880 2688 15944 2692
rect 15960 2748 16024 2752
rect 15960 2692 15964 2748
rect 15964 2692 16020 2748
rect 16020 2692 16024 2748
rect 15960 2688 16024 2692
rect 16040 2748 16104 2752
rect 16040 2692 16044 2748
rect 16044 2692 16100 2748
rect 16100 2692 16104 2748
rect 16040 2688 16104 2692
rect 16120 2748 16184 2752
rect 16120 2692 16124 2748
rect 16124 2692 16180 2748
rect 16180 2692 16184 2748
rect 16120 2688 16184 2692
rect 5030 2204 5094 2208
rect 5030 2148 5034 2204
rect 5034 2148 5090 2204
rect 5090 2148 5094 2204
rect 5030 2144 5094 2148
rect 5110 2204 5174 2208
rect 5110 2148 5114 2204
rect 5114 2148 5170 2204
rect 5170 2148 5174 2204
rect 5110 2144 5174 2148
rect 5190 2204 5254 2208
rect 5190 2148 5194 2204
rect 5194 2148 5250 2204
rect 5250 2148 5254 2204
rect 5190 2144 5254 2148
rect 5270 2204 5334 2208
rect 5270 2148 5274 2204
rect 5274 2148 5330 2204
rect 5330 2148 5334 2204
rect 5270 2144 5334 2148
rect 8130 2204 8194 2208
rect 8130 2148 8134 2204
rect 8134 2148 8190 2204
rect 8190 2148 8194 2204
rect 8130 2144 8194 2148
rect 8210 2204 8274 2208
rect 8210 2148 8214 2204
rect 8214 2148 8270 2204
rect 8270 2148 8274 2204
rect 8210 2144 8274 2148
rect 8290 2204 8354 2208
rect 8290 2148 8294 2204
rect 8294 2148 8350 2204
rect 8350 2148 8354 2204
rect 8290 2144 8354 2148
rect 8370 2204 8434 2208
rect 8370 2148 8374 2204
rect 8374 2148 8430 2204
rect 8430 2148 8434 2204
rect 8370 2144 8434 2148
rect 11230 2204 11294 2208
rect 11230 2148 11234 2204
rect 11234 2148 11290 2204
rect 11290 2148 11294 2204
rect 11230 2144 11294 2148
rect 11310 2204 11374 2208
rect 11310 2148 11314 2204
rect 11314 2148 11370 2204
rect 11370 2148 11374 2204
rect 11310 2144 11374 2148
rect 11390 2204 11454 2208
rect 11390 2148 11394 2204
rect 11394 2148 11450 2204
rect 11450 2148 11454 2204
rect 11390 2144 11454 2148
rect 11470 2204 11534 2208
rect 11470 2148 11474 2204
rect 11474 2148 11530 2204
rect 11530 2148 11534 2204
rect 11470 2144 11534 2148
rect 14330 2204 14394 2208
rect 14330 2148 14334 2204
rect 14334 2148 14390 2204
rect 14390 2148 14394 2204
rect 14330 2144 14394 2148
rect 14410 2204 14474 2208
rect 14410 2148 14414 2204
rect 14414 2148 14470 2204
rect 14470 2148 14474 2204
rect 14410 2144 14474 2148
rect 14490 2204 14554 2208
rect 14490 2148 14494 2204
rect 14494 2148 14550 2204
rect 14550 2148 14554 2204
rect 14490 2144 14554 2148
rect 14570 2204 14634 2208
rect 14570 2148 14574 2204
rect 14574 2148 14630 2204
rect 14630 2148 14634 2204
rect 14570 2144 14634 2148
rect 17430 2204 17494 2208
rect 17430 2148 17434 2204
rect 17434 2148 17490 2204
rect 17490 2148 17494 2204
rect 17430 2144 17494 2148
rect 17510 2204 17574 2208
rect 17510 2148 17514 2204
rect 17514 2148 17570 2204
rect 17570 2148 17574 2204
rect 17510 2144 17574 2148
rect 17590 2204 17654 2208
rect 17590 2148 17594 2204
rect 17594 2148 17650 2204
rect 17650 2148 17654 2204
rect 17590 2144 17654 2148
rect 17670 2204 17734 2208
rect 17670 2148 17674 2204
rect 17674 2148 17730 2204
rect 17730 2148 17734 2204
rect 17670 2144 17734 2148
rect 3480 1660 3544 1664
rect 3480 1604 3484 1660
rect 3484 1604 3540 1660
rect 3540 1604 3544 1660
rect 3480 1600 3544 1604
rect 3560 1660 3624 1664
rect 3560 1604 3564 1660
rect 3564 1604 3620 1660
rect 3620 1604 3624 1660
rect 3560 1600 3624 1604
rect 3640 1660 3704 1664
rect 3640 1604 3644 1660
rect 3644 1604 3700 1660
rect 3700 1604 3704 1660
rect 3640 1600 3704 1604
rect 3720 1660 3784 1664
rect 3720 1604 3724 1660
rect 3724 1604 3780 1660
rect 3780 1604 3784 1660
rect 3720 1600 3784 1604
rect 6580 1660 6644 1664
rect 6580 1604 6584 1660
rect 6584 1604 6640 1660
rect 6640 1604 6644 1660
rect 6580 1600 6644 1604
rect 6660 1660 6724 1664
rect 6660 1604 6664 1660
rect 6664 1604 6720 1660
rect 6720 1604 6724 1660
rect 6660 1600 6724 1604
rect 6740 1660 6804 1664
rect 6740 1604 6744 1660
rect 6744 1604 6800 1660
rect 6800 1604 6804 1660
rect 6740 1600 6804 1604
rect 6820 1660 6884 1664
rect 6820 1604 6824 1660
rect 6824 1604 6880 1660
rect 6880 1604 6884 1660
rect 6820 1600 6884 1604
rect 9680 1660 9744 1664
rect 9680 1604 9684 1660
rect 9684 1604 9740 1660
rect 9740 1604 9744 1660
rect 9680 1600 9744 1604
rect 9760 1660 9824 1664
rect 9760 1604 9764 1660
rect 9764 1604 9820 1660
rect 9820 1604 9824 1660
rect 9760 1600 9824 1604
rect 9840 1660 9904 1664
rect 9840 1604 9844 1660
rect 9844 1604 9900 1660
rect 9900 1604 9904 1660
rect 9840 1600 9904 1604
rect 9920 1660 9984 1664
rect 9920 1604 9924 1660
rect 9924 1604 9980 1660
rect 9980 1604 9984 1660
rect 9920 1600 9984 1604
rect 12780 1660 12844 1664
rect 12780 1604 12784 1660
rect 12784 1604 12840 1660
rect 12840 1604 12844 1660
rect 12780 1600 12844 1604
rect 12860 1660 12924 1664
rect 12860 1604 12864 1660
rect 12864 1604 12920 1660
rect 12920 1604 12924 1660
rect 12860 1600 12924 1604
rect 12940 1660 13004 1664
rect 12940 1604 12944 1660
rect 12944 1604 13000 1660
rect 13000 1604 13004 1660
rect 12940 1600 13004 1604
rect 13020 1660 13084 1664
rect 13020 1604 13024 1660
rect 13024 1604 13080 1660
rect 13080 1604 13084 1660
rect 13020 1600 13084 1604
rect 15880 1660 15944 1664
rect 15880 1604 15884 1660
rect 15884 1604 15940 1660
rect 15940 1604 15944 1660
rect 15880 1600 15944 1604
rect 15960 1660 16024 1664
rect 15960 1604 15964 1660
rect 15964 1604 16020 1660
rect 16020 1604 16024 1660
rect 15960 1600 16024 1604
rect 16040 1660 16104 1664
rect 16040 1604 16044 1660
rect 16044 1604 16100 1660
rect 16100 1604 16104 1660
rect 16040 1600 16104 1604
rect 16120 1660 16184 1664
rect 16120 1604 16124 1660
rect 16124 1604 16180 1660
rect 16180 1604 16184 1660
rect 16120 1600 16184 1604
rect 5030 1116 5094 1120
rect 5030 1060 5034 1116
rect 5034 1060 5090 1116
rect 5090 1060 5094 1116
rect 5030 1056 5094 1060
rect 5110 1116 5174 1120
rect 5110 1060 5114 1116
rect 5114 1060 5170 1116
rect 5170 1060 5174 1116
rect 5110 1056 5174 1060
rect 5190 1116 5254 1120
rect 5190 1060 5194 1116
rect 5194 1060 5250 1116
rect 5250 1060 5254 1116
rect 5190 1056 5254 1060
rect 5270 1116 5334 1120
rect 5270 1060 5274 1116
rect 5274 1060 5330 1116
rect 5330 1060 5334 1116
rect 5270 1056 5334 1060
rect 8130 1116 8194 1120
rect 8130 1060 8134 1116
rect 8134 1060 8190 1116
rect 8190 1060 8194 1116
rect 8130 1056 8194 1060
rect 8210 1116 8274 1120
rect 8210 1060 8214 1116
rect 8214 1060 8270 1116
rect 8270 1060 8274 1116
rect 8210 1056 8274 1060
rect 8290 1116 8354 1120
rect 8290 1060 8294 1116
rect 8294 1060 8350 1116
rect 8350 1060 8354 1116
rect 8290 1056 8354 1060
rect 8370 1116 8434 1120
rect 8370 1060 8374 1116
rect 8374 1060 8430 1116
rect 8430 1060 8434 1116
rect 8370 1056 8434 1060
rect 11230 1116 11294 1120
rect 11230 1060 11234 1116
rect 11234 1060 11290 1116
rect 11290 1060 11294 1116
rect 11230 1056 11294 1060
rect 11310 1116 11374 1120
rect 11310 1060 11314 1116
rect 11314 1060 11370 1116
rect 11370 1060 11374 1116
rect 11310 1056 11374 1060
rect 11390 1116 11454 1120
rect 11390 1060 11394 1116
rect 11394 1060 11450 1116
rect 11450 1060 11454 1116
rect 11390 1056 11454 1060
rect 11470 1116 11534 1120
rect 11470 1060 11474 1116
rect 11474 1060 11530 1116
rect 11530 1060 11534 1116
rect 11470 1056 11534 1060
rect 14330 1116 14394 1120
rect 14330 1060 14334 1116
rect 14334 1060 14390 1116
rect 14390 1060 14394 1116
rect 14330 1056 14394 1060
rect 14410 1116 14474 1120
rect 14410 1060 14414 1116
rect 14414 1060 14470 1116
rect 14470 1060 14474 1116
rect 14410 1056 14474 1060
rect 14490 1116 14554 1120
rect 14490 1060 14494 1116
rect 14494 1060 14550 1116
rect 14550 1060 14554 1116
rect 14490 1056 14554 1060
rect 14570 1116 14634 1120
rect 14570 1060 14574 1116
rect 14574 1060 14630 1116
rect 14630 1060 14634 1116
rect 14570 1056 14634 1060
rect 17430 1116 17494 1120
rect 17430 1060 17434 1116
rect 17434 1060 17490 1116
rect 17490 1060 17494 1116
rect 17430 1056 17494 1060
rect 17510 1116 17574 1120
rect 17510 1060 17514 1116
rect 17514 1060 17570 1116
rect 17570 1060 17574 1116
rect 17510 1056 17574 1060
rect 17590 1116 17654 1120
rect 17590 1060 17594 1116
rect 17594 1060 17650 1116
rect 17650 1060 17654 1116
rect 17590 1056 17654 1060
rect 17670 1116 17734 1120
rect 17670 1060 17674 1116
rect 17674 1060 17730 1116
rect 17730 1060 17734 1116
rect 17670 1056 17734 1060
rect 3480 572 3544 576
rect 3480 516 3484 572
rect 3484 516 3540 572
rect 3540 516 3544 572
rect 3480 512 3544 516
rect 3560 572 3624 576
rect 3560 516 3564 572
rect 3564 516 3620 572
rect 3620 516 3624 572
rect 3560 512 3624 516
rect 3640 572 3704 576
rect 3640 516 3644 572
rect 3644 516 3700 572
rect 3700 516 3704 572
rect 3640 512 3704 516
rect 3720 572 3784 576
rect 3720 516 3724 572
rect 3724 516 3780 572
rect 3780 516 3784 572
rect 3720 512 3784 516
rect 6580 572 6644 576
rect 6580 516 6584 572
rect 6584 516 6640 572
rect 6640 516 6644 572
rect 6580 512 6644 516
rect 6660 572 6724 576
rect 6660 516 6664 572
rect 6664 516 6720 572
rect 6720 516 6724 572
rect 6660 512 6724 516
rect 6740 572 6804 576
rect 6740 516 6744 572
rect 6744 516 6800 572
rect 6800 516 6804 572
rect 6740 512 6804 516
rect 6820 572 6884 576
rect 6820 516 6824 572
rect 6824 516 6880 572
rect 6880 516 6884 572
rect 6820 512 6884 516
rect 9680 572 9744 576
rect 9680 516 9684 572
rect 9684 516 9740 572
rect 9740 516 9744 572
rect 9680 512 9744 516
rect 9760 572 9824 576
rect 9760 516 9764 572
rect 9764 516 9820 572
rect 9820 516 9824 572
rect 9760 512 9824 516
rect 9840 572 9904 576
rect 9840 516 9844 572
rect 9844 516 9900 572
rect 9900 516 9904 572
rect 9840 512 9904 516
rect 9920 572 9984 576
rect 9920 516 9924 572
rect 9924 516 9980 572
rect 9980 516 9984 572
rect 9920 512 9984 516
rect 12780 572 12844 576
rect 12780 516 12784 572
rect 12784 516 12840 572
rect 12840 516 12844 572
rect 12780 512 12844 516
rect 12860 572 12924 576
rect 12860 516 12864 572
rect 12864 516 12920 572
rect 12920 516 12924 572
rect 12860 512 12924 516
rect 12940 572 13004 576
rect 12940 516 12944 572
rect 12944 516 13000 572
rect 13000 516 13004 572
rect 12940 512 13004 516
rect 13020 572 13084 576
rect 13020 516 13024 572
rect 13024 516 13080 572
rect 13080 516 13084 572
rect 13020 512 13084 516
rect 15880 572 15944 576
rect 15880 516 15884 572
rect 15884 516 15940 572
rect 15940 516 15944 572
rect 15880 512 15944 516
rect 15960 572 16024 576
rect 15960 516 15964 572
rect 15964 516 16020 572
rect 16020 516 16024 572
rect 15960 512 16024 516
rect 16040 572 16104 576
rect 16040 516 16044 572
rect 16044 516 16100 572
rect 16100 516 16104 572
rect 16040 512 16104 516
rect 16120 572 16184 576
rect 16120 516 16124 572
rect 16124 516 16180 572
rect 16180 516 16184 572
rect 16120 512 16184 516
rect 5030 28 5094 32
rect 5030 -28 5034 28
rect 5034 -28 5090 28
rect 5090 -28 5094 28
rect 5030 -32 5094 -28
rect 5110 28 5174 32
rect 5110 -28 5114 28
rect 5114 -28 5170 28
rect 5170 -28 5174 28
rect 5110 -32 5174 -28
rect 5190 28 5254 32
rect 5190 -28 5194 28
rect 5194 -28 5250 28
rect 5250 -28 5254 28
rect 5190 -32 5254 -28
rect 5270 28 5334 32
rect 5270 -28 5274 28
rect 5274 -28 5330 28
rect 5330 -28 5334 28
rect 5270 -32 5334 -28
rect 8130 28 8194 32
rect 8130 -28 8134 28
rect 8134 -28 8190 28
rect 8190 -28 8194 28
rect 8130 -32 8194 -28
rect 8210 28 8274 32
rect 8210 -28 8214 28
rect 8214 -28 8270 28
rect 8270 -28 8274 28
rect 8210 -32 8274 -28
rect 8290 28 8354 32
rect 8290 -28 8294 28
rect 8294 -28 8350 28
rect 8350 -28 8354 28
rect 8290 -32 8354 -28
rect 8370 28 8434 32
rect 8370 -28 8374 28
rect 8374 -28 8430 28
rect 8430 -28 8434 28
rect 8370 -32 8434 -28
rect 11230 28 11294 32
rect 11230 -28 11234 28
rect 11234 -28 11290 28
rect 11290 -28 11294 28
rect 11230 -32 11294 -28
rect 11310 28 11374 32
rect 11310 -28 11314 28
rect 11314 -28 11370 28
rect 11370 -28 11374 28
rect 11310 -32 11374 -28
rect 11390 28 11454 32
rect 11390 -28 11394 28
rect 11394 -28 11450 28
rect 11450 -28 11454 28
rect 11390 -32 11454 -28
rect 11470 28 11534 32
rect 11470 -28 11474 28
rect 11474 -28 11530 28
rect 11530 -28 11534 28
rect 11470 -32 11534 -28
rect 14330 28 14394 32
rect 14330 -28 14334 28
rect 14334 -28 14390 28
rect 14390 -28 14394 28
rect 14330 -32 14394 -28
rect 14410 28 14474 32
rect 14410 -28 14414 28
rect 14414 -28 14470 28
rect 14470 -28 14474 28
rect 14410 -32 14474 -28
rect 14490 28 14554 32
rect 14490 -28 14494 28
rect 14494 -28 14550 28
rect 14550 -28 14554 28
rect 14490 -32 14554 -28
rect 14570 28 14634 32
rect 14570 -28 14574 28
rect 14574 -28 14630 28
rect 14630 -28 14634 28
rect 14570 -32 14634 -28
rect 17430 28 17494 32
rect 17430 -28 17434 28
rect 17434 -28 17490 28
rect 17490 -28 17494 28
rect 17430 -32 17494 -28
rect 17510 28 17574 32
rect 17510 -28 17514 28
rect 17514 -28 17570 28
rect 17570 -28 17574 28
rect 17510 -32 17574 -28
rect 17590 28 17654 32
rect 17590 -28 17594 28
rect 17594 -28 17650 28
rect 17650 -28 17654 28
rect 17590 -32 17654 -28
rect 17670 28 17734 32
rect 17670 -28 17674 28
rect 17674 -28 17730 28
rect 17730 -28 17734 28
rect 17670 -32 17734 -28
<< metal4 >>
rect 3472 10368 3792 10928
rect 3472 10304 3480 10368
rect 3544 10304 3560 10368
rect 3624 10304 3640 10368
rect 3704 10304 3720 10368
rect 3784 10304 3792 10368
rect 3472 10160 3792 10304
rect 3472 9924 3514 10160
rect 3750 9924 3792 10160
rect 3472 9280 3792 9924
rect 3472 9216 3480 9280
rect 3544 9216 3560 9280
rect 3624 9216 3640 9280
rect 3704 9216 3720 9280
rect 3784 9216 3792 9280
rect 3472 8192 3792 9216
rect 3472 8128 3480 8192
rect 3544 8128 3560 8192
rect 3624 8128 3640 8192
rect 3704 8128 3720 8192
rect 3784 8128 3792 8192
rect 3472 7104 3792 8128
rect 3472 7040 3480 7104
rect 3544 7040 3560 7104
rect 3624 7040 3640 7104
rect 3704 7040 3720 7104
rect 3784 7040 3792 7104
rect 3472 6780 3792 7040
rect 3472 6544 3514 6780
rect 3750 6544 3792 6780
rect 3472 6016 3792 6544
rect 3472 5952 3480 6016
rect 3544 5952 3560 6016
rect 3624 5952 3640 6016
rect 3704 5952 3720 6016
rect 3784 5952 3792 6016
rect 3472 4928 3792 5952
rect 3472 4864 3480 4928
rect 3544 4864 3560 4928
rect 3624 4864 3640 4928
rect 3704 4864 3720 4928
rect 3784 4864 3792 4928
rect 3472 3840 3792 4864
rect 3472 3776 3480 3840
rect 3544 3776 3560 3840
rect 3624 3776 3640 3840
rect 3704 3776 3720 3840
rect 3784 3776 3792 3840
rect 3472 3400 3792 3776
rect 3472 3164 3514 3400
rect 3750 3164 3792 3400
rect 3472 2752 3792 3164
rect 3472 2688 3480 2752
rect 3544 2688 3560 2752
rect 3624 2688 3640 2752
rect 3704 2688 3720 2752
rect 3784 2688 3792 2752
rect 3472 1664 3792 2688
rect 3472 1600 3480 1664
rect 3544 1600 3560 1664
rect 3624 1600 3640 1664
rect 3704 1600 3720 1664
rect 3784 1600 3792 1664
rect 3472 576 3792 1600
rect 3472 512 3480 576
rect 3544 512 3560 576
rect 3624 512 3640 576
rect 3704 512 3720 576
rect 3784 512 3792 576
rect 3472 -48 3792 512
rect 5022 10912 5342 10928
rect 5022 10848 5030 10912
rect 5094 10848 5110 10912
rect 5174 10848 5190 10912
rect 5254 10848 5270 10912
rect 5334 10848 5342 10912
rect 5022 9824 5342 10848
rect 5022 9760 5030 9824
rect 5094 9760 5110 9824
rect 5174 9760 5190 9824
rect 5254 9760 5270 9824
rect 5334 9760 5342 9824
rect 5022 8736 5342 9760
rect 5022 8672 5030 8736
rect 5094 8672 5110 8736
rect 5174 8672 5190 8736
rect 5254 8672 5270 8736
rect 5334 8672 5342 8736
rect 5022 8470 5342 8672
rect 5022 8234 5064 8470
rect 5300 8234 5342 8470
rect 5022 7648 5342 8234
rect 5022 7584 5030 7648
rect 5094 7584 5110 7648
rect 5174 7584 5190 7648
rect 5254 7584 5270 7648
rect 5334 7584 5342 7648
rect 5022 6560 5342 7584
rect 5022 6496 5030 6560
rect 5094 6496 5110 6560
rect 5174 6496 5190 6560
rect 5254 6496 5270 6560
rect 5334 6496 5342 6560
rect 5022 5472 5342 6496
rect 5022 5408 5030 5472
rect 5094 5408 5110 5472
rect 5174 5408 5190 5472
rect 5254 5408 5270 5472
rect 5334 5408 5342 5472
rect 5022 5090 5342 5408
rect 5022 4854 5064 5090
rect 5300 4854 5342 5090
rect 5022 4384 5342 4854
rect 5022 4320 5030 4384
rect 5094 4320 5110 4384
rect 5174 4320 5190 4384
rect 5254 4320 5270 4384
rect 5334 4320 5342 4384
rect 5022 3296 5342 4320
rect 5022 3232 5030 3296
rect 5094 3232 5110 3296
rect 5174 3232 5190 3296
rect 5254 3232 5270 3296
rect 5334 3232 5342 3296
rect 5022 2208 5342 3232
rect 5022 2144 5030 2208
rect 5094 2144 5110 2208
rect 5174 2144 5190 2208
rect 5254 2144 5270 2208
rect 5334 2144 5342 2208
rect 5022 1120 5342 2144
rect 5022 1056 5030 1120
rect 5094 1056 5110 1120
rect 5174 1056 5190 1120
rect 5254 1056 5270 1120
rect 5334 1056 5342 1120
rect 5022 32 5342 1056
rect 5022 -32 5030 32
rect 5094 -32 5110 32
rect 5174 -32 5190 32
rect 5254 -32 5270 32
rect 5334 -32 5342 32
rect 5022 -48 5342 -32
rect 6572 10368 6892 10928
rect 6572 10304 6580 10368
rect 6644 10304 6660 10368
rect 6724 10304 6740 10368
rect 6804 10304 6820 10368
rect 6884 10304 6892 10368
rect 6572 10160 6892 10304
rect 6572 9924 6614 10160
rect 6850 9924 6892 10160
rect 6572 9280 6892 9924
rect 6572 9216 6580 9280
rect 6644 9216 6660 9280
rect 6724 9216 6740 9280
rect 6804 9216 6820 9280
rect 6884 9216 6892 9280
rect 6572 8192 6892 9216
rect 6572 8128 6580 8192
rect 6644 8128 6660 8192
rect 6724 8128 6740 8192
rect 6804 8128 6820 8192
rect 6884 8128 6892 8192
rect 6572 7104 6892 8128
rect 6572 7040 6580 7104
rect 6644 7040 6660 7104
rect 6724 7040 6740 7104
rect 6804 7040 6820 7104
rect 6884 7040 6892 7104
rect 6572 6780 6892 7040
rect 6572 6544 6614 6780
rect 6850 6544 6892 6780
rect 6572 6016 6892 6544
rect 6572 5952 6580 6016
rect 6644 5952 6660 6016
rect 6724 5952 6740 6016
rect 6804 5952 6820 6016
rect 6884 5952 6892 6016
rect 6572 4928 6892 5952
rect 6572 4864 6580 4928
rect 6644 4864 6660 4928
rect 6724 4864 6740 4928
rect 6804 4864 6820 4928
rect 6884 4864 6892 4928
rect 6572 3840 6892 4864
rect 6572 3776 6580 3840
rect 6644 3776 6660 3840
rect 6724 3776 6740 3840
rect 6804 3776 6820 3840
rect 6884 3776 6892 3840
rect 6572 3400 6892 3776
rect 6572 3164 6614 3400
rect 6850 3164 6892 3400
rect 6572 2752 6892 3164
rect 6572 2688 6580 2752
rect 6644 2688 6660 2752
rect 6724 2688 6740 2752
rect 6804 2688 6820 2752
rect 6884 2688 6892 2752
rect 6572 1664 6892 2688
rect 6572 1600 6580 1664
rect 6644 1600 6660 1664
rect 6724 1600 6740 1664
rect 6804 1600 6820 1664
rect 6884 1600 6892 1664
rect 6572 576 6892 1600
rect 6572 512 6580 576
rect 6644 512 6660 576
rect 6724 512 6740 576
rect 6804 512 6820 576
rect 6884 512 6892 576
rect 6572 -48 6892 512
rect 8122 10912 8442 10928
rect 8122 10848 8130 10912
rect 8194 10848 8210 10912
rect 8274 10848 8290 10912
rect 8354 10848 8370 10912
rect 8434 10848 8442 10912
rect 8122 9824 8442 10848
rect 8122 9760 8130 9824
rect 8194 9760 8210 9824
rect 8274 9760 8290 9824
rect 8354 9760 8370 9824
rect 8434 9760 8442 9824
rect 8122 8736 8442 9760
rect 8122 8672 8130 8736
rect 8194 8672 8210 8736
rect 8274 8672 8290 8736
rect 8354 8672 8370 8736
rect 8434 8672 8442 8736
rect 8122 8470 8442 8672
rect 8122 8234 8164 8470
rect 8400 8234 8442 8470
rect 8122 7648 8442 8234
rect 8122 7584 8130 7648
rect 8194 7584 8210 7648
rect 8274 7584 8290 7648
rect 8354 7584 8370 7648
rect 8434 7584 8442 7648
rect 8122 6560 8442 7584
rect 8122 6496 8130 6560
rect 8194 6496 8210 6560
rect 8274 6496 8290 6560
rect 8354 6496 8370 6560
rect 8434 6496 8442 6560
rect 8122 5472 8442 6496
rect 8122 5408 8130 5472
rect 8194 5408 8210 5472
rect 8274 5408 8290 5472
rect 8354 5408 8370 5472
rect 8434 5408 8442 5472
rect 8122 5090 8442 5408
rect 8122 4854 8164 5090
rect 8400 4854 8442 5090
rect 8122 4384 8442 4854
rect 8122 4320 8130 4384
rect 8194 4320 8210 4384
rect 8274 4320 8290 4384
rect 8354 4320 8370 4384
rect 8434 4320 8442 4384
rect 8122 3296 8442 4320
rect 8122 3232 8130 3296
rect 8194 3232 8210 3296
rect 8274 3232 8290 3296
rect 8354 3232 8370 3296
rect 8434 3232 8442 3296
rect 8122 2208 8442 3232
rect 8122 2144 8130 2208
rect 8194 2144 8210 2208
rect 8274 2144 8290 2208
rect 8354 2144 8370 2208
rect 8434 2144 8442 2208
rect 8122 1120 8442 2144
rect 8122 1056 8130 1120
rect 8194 1056 8210 1120
rect 8274 1056 8290 1120
rect 8354 1056 8370 1120
rect 8434 1056 8442 1120
rect 8122 32 8442 1056
rect 8122 -32 8130 32
rect 8194 -32 8210 32
rect 8274 -32 8290 32
rect 8354 -32 8370 32
rect 8434 -32 8442 32
rect 8122 -48 8442 -32
rect 9672 10368 9992 10928
rect 9672 10304 9680 10368
rect 9744 10304 9760 10368
rect 9824 10304 9840 10368
rect 9904 10304 9920 10368
rect 9984 10304 9992 10368
rect 9672 10160 9992 10304
rect 9672 9924 9714 10160
rect 9950 9924 9992 10160
rect 9672 9280 9992 9924
rect 9672 9216 9680 9280
rect 9744 9216 9760 9280
rect 9824 9216 9840 9280
rect 9904 9216 9920 9280
rect 9984 9216 9992 9280
rect 9672 8192 9992 9216
rect 9672 8128 9680 8192
rect 9744 8128 9760 8192
rect 9824 8128 9840 8192
rect 9904 8128 9920 8192
rect 9984 8128 9992 8192
rect 9672 7104 9992 8128
rect 9672 7040 9680 7104
rect 9744 7040 9760 7104
rect 9824 7040 9840 7104
rect 9904 7040 9920 7104
rect 9984 7040 9992 7104
rect 9672 6780 9992 7040
rect 9672 6544 9714 6780
rect 9950 6544 9992 6780
rect 9672 6016 9992 6544
rect 9672 5952 9680 6016
rect 9744 5952 9760 6016
rect 9824 5952 9840 6016
rect 9904 5952 9920 6016
rect 9984 5952 9992 6016
rect 9672 4928 9992 5952
rect 9672 4864 9680 4928
rect 9744 4864 9760 4928
rect 9824 4864 9840 4928
rect 9904 4864 9920 4928
rect 9984 4864 9992 4928
rect 9672 3840 9992 4864
rect 9672 3776 9680 3840
rect 9744 3776 9760 3840
rect 9824 3776 9840 3840
rect 9904 3776 9920 3840
rect 9984 3776 9992 3840
rect 9672 3400 9992 3776
rect 9672 3164 9714 3400
rect 9950 3164 9992 3400
rect 9672 2752 9992 3164
rect 9672 2688 9680 2752
rect 9744 2688 9760 2752
rect 9824 2688 9840 2752
rect 9904 2688 9920 2752
rect 9984 2688 9992 2752
rect 9672 1664 9992 2688
rect 9672 1600 9680 1664
rect 9744 1600 9760 1664
rect 9824 1600 9840 1664
rect 9904 1600 9920 1664
rect 9984 1600 9992 1664
rect 9672 576 9992 1600
rect 9672 512 9680 576
rect 9744 512 9760 576
rect 9824 512 9840 576
rect 9904 512 9920 576
rect 9984 512 9992 576
rect 9672 -48 9992 512
rect 11222 10912 11542 10928
rect 11222 10848 11230 10912
rect 11294 10848 11310 10912
rect 11374 10848 11390 10912
rect 11454 10848 11470 10912
rect 11534 10848 11542 10912
rect 11222 9824 11542 10848
rect 11222 9760 11230 9824
rect 11294 9760 11310 9824
rect 11374 9760 11390 9824
rect 11454 9760 11470 9824
rect 11534 9760 11542 9824
rect 11222 8736 11542 9760
rect 11222 8672 11230 8736
rect 11294 8672 11310 8736
rect 11374 8672 11390 8736
rect 11454 8672 11470 8736
rect 11534 8672 11542 8736
rect 11222 8470 11542 8672
rect 11222 8234 11264 8470
rect 11500 8234 11542 8470
rect 11222 7648 11542 8234
rect 11222 7584 11230 7648
rect 11294 7584 11310 7648
rect 11374 7584 11390 7648
rect 11454 7584 11470 7648
rect 11534 7584 11542 7648
rect 11222 6560 11542 7584
rect 11222 6496 11230 6560
rect 11294 6496 11310 6560
rect 11374 6496 11390 6560
rect 11454 6496 11470 6560
rect 11534 6496 11542 6560
rect 11222 5472 11542 6496
rect 11222 5408 11230 5472
rect 11294 5408 11310 5472
rect 11374 5408 11390 5472
rect 11454 5408 11470 5472
rect 11534 5408 11542 5472
rect 11222 5090 11542 5408
rect 11222 4854 11264 5090
rect 11500 4854 11542 5090
rect 11222 4384 11542 4854
rect 11222 4320 11230 4384
rect 11294 4320 11310 4384
rect 11374 4320 11390 4384
rect 11454 4320 11470 4384
rect 11534 4320 11542 4384
rect 11222 3296 11542 4320
rect 11222 3232 11230 3296
rect 11294 3232 11310 3296
rect 11374 3232 11390 3296
rect 11454 3232 11470 3296
rect 11534 3232 11542 3296
rect 11222 2208 11542 3232
rect 11222 2144 11230 2208
rect 11294 2144 11310 2208
rect 11374 2144 11390 2208
rect 11454 2144 11470 2208
rect 11534 2144 11542 2208
rect 11222 1120 11542 2144
rect 11222 1056 11230 1120
rect 11294 1056 11310 1120
rect 11374 1056 11390 1120
rect 11454 1056 11470 1120
rect 11534 1056 11542 1120
rect 11222 32 11542 1056
rect 11222 -32 11230 32
rect 11294 -32 11310 32
rect 11374 -32 11390 32
rect 11454 -32 11470 32
rect 11534 -32 11542 32
rect 11222 -48 11542 -32
rect 12772 10368 13092 10928
rect 12772 10304 12780 10368
rect 12844 10304 12860 10368
rect 12924 10304 12940 10368
rect 13004 10304 13020 10368
rect 13084 10304 13092 10368
rect 12772 10160 13092 10304
rect 12772 9924 12814 10160
rect 13050 9924 13092 10160
rect 12772 9280 13092 9924
rect 12772 9216 12780 9280
rect 12844 9216 12860 9280
rect 12924 9216 12940 9280
rect 13004 9216 13020 9280
rect 13084 9216 13092 9280
rect 12772 8192 13092 9216
rect 12772 8128 12780 8192
rect 12844 8128 12860 8192
rect 12924 8128 12940 8192
rect 13004 8128 13020 8192
rect 13084 8128 13092 8192
rect 12772 7104 13092 8128
rect 12772 7040 12780 7104
rect 12844 7040 12860 7104
rect 12924 7040 12940 7104
rect 13004 7040 13020 7104
rect 13084 7040 13092 7104
rect 12772 6780 13092 7040
rect 12772 6544 12814 6780
rect 13050 6544 13092 6780
rect 12772 6016 13092 6544
rect 12772 5952 12780 6016
rect 12844 5952 12860 6016
rect 12924 5952 12940 6016
rect 13004 5952 13020 6016
rect 13084 5952 13092 6016
rect 12772 4928 13092 5952
rect 12772 4864 12780 4928
rect 12844 4864 12860 4928
rect 12924 4864 12940 4928
rect 13004 4864 13020 4928
rect 13084 4864 13092 4928
rect 12772 3840 13092 4864
rect 12772 3776 12780 3840
rect 12844 3776 12860 3840
rect 12924 3776 12940 3840
rect 13004 3776 13020 3840
rect 13084 3776 13092 3840
rect 12772 3400 13092 3776
rect 12772 3164 12814 3400
rect 13050 3164 13092 3400
rect 12772 2752 13092 3164
rect 12772 2688 12780 2752
rect 12844 2688 12860 2752
rect 12924 2688 12940 2752
rect 13004 2688 13020 2752
rect 13084 2688 13092 2752
rect 12772 1664 13092 2688
rect 12772 1600 12780 1664
rect 12844 1600 12860 1664
rect 12924 1600 12940 1664
rect 13004 1600 13020 1664
rect 13084 1600 13092 1664
rect 12772 576 13092 1600
rect 12772 512 12780 576
rect 12844 512 12860 576
rect 12924 512 12940 576
rect 13004 512 13020 576
rect 13084 512 13092 576
rect 12772 -48 13092 512
rect 14322 10912 14642 10928
rect 14322 10848 14330 10912
rect 14394 10848 14410 10912
rect 14474 10848 14490 10912
rect 14554 10848 14570 10912
rect 14634 10848 14642 10912
rect 14322 9824 14642 10848
rect 14322 9760 14330 9824
rect 14394 9760 14410 9824
rect 14474 9760 14490 9824
rect 14554 9760 14570 9824
rect 14634 9760 14642 9824
rect 14322 8736 14642 9760
rect 14322 8672 14330 8736
rect 14394 8672 14410 8736
rect 14474 8672 14490 8736
rect 14554 8672 14570 8736
rect 14634 8672 14642 8736
rect 14322 8470 14642 8672
rect 14322 8234 14364 8470
rect 14600 8234 14642 8470
rect 14322 7648 14642 8234
rect 14322 7584 14330 7648
rect 14394 7584 14410 7648
rect 14474 7584 14490 7648
rect 14554 7584 14570 7648
rect 14634 7584 14642 7648
rect 14322 6560 14642 7584
rect 14322 6496 14330 6560
rect 14394 6496 14410 6560
rect 14474 6496 14490 6560
rect 14554 6496 14570 6560
rect 14634 6496 14642 6560
rect 14322 5472 14642 6496
rect 14322 5408 14330 5472
rect 14394 5408 14410 5472
rect 14474 5408 14490 5472
rect 14554 5408 14570 5472
rect 14634 5408 14642 5472
rect 14322 5090 14642 5408
rect 14322 4854 14364 5090
rect 14600 4854 14642 5090
rect 14322 4384 14642 4854
rect 14322 4320 14330 4384
rect 14394 4320 14410 4384
rect 14474 4320 14490 4384
rect 14554 4320 14570 4384
rect 14634 4320 14642 4384
rect 14322 3296 14642 4320
rect 14322 3232 14330 3296
rect 14394 3232 14410 3296
rect 14474 3232 14490 3296
rect 14554 3232 14570 3296
rect 14634 3232 14642 3296
rect 14322 2208 14642 3232
rect 14322 2144 14330 2208
rect 14394 2144 14410 2208
rect 14474 2144 14490 2208
rect 14554 2144 14570 2208
rect 14634 2144 14642 2208
rect 14322 1120 14642 2144
rect 14322 1056 14330 1120
rect 14394 1056 14410 1120
rect 14474 1056 14490 1120
rect 14554 1056 14570 1120
rect 14634 1056 14642 1120
rect 14322 32 14642 1056
rect 14322 -32 14330 32
rect 14394 -32 14410 32
rect 14474 -32 14490 32
rect 14554 -32 14570 32
rect 14634 -32 14642 32
rect 14322 -48 14642 -32
rect 15872 10368 16192 10928
rect 15872 10304 15880 10368
rect 15944 10304 15960 10368
rect 16024 10304 16040 10368
rect 16104 10304 16120 10368
rect 16184 10304 16192 10368
rect 15872 10160 16192 10304
rect 15872 9924 15914 10160
rect 16150 9924 16192 10160
rect 15872 9280 16192 9924
rect 15872 9216 15880 9280
rect 15944 9216 15960 9280
rect 16024 9216 16040 9280
rect 16104 9216 16120 9280
rect 16184 9216 16192 9280
rect 15872 8192 16192 9216
rect 15872 8128 15880 8192
rect 15944 8128 15960 8192
rect 16024 8128 16040 8192
rect 16104 8128 16120 8192
rect 16184 8128 16192 8192
rect 15872 7104 16192 8128
rect 15872 7040 15880 7104
rect 15944 7040 15960 7104
rect 16024 7040 16040 7104
rect 16104 7040 16120 7104
rect 16184 7040 16192 7104
rect 15872 6780 16192 7040
rect 15872 6544 15914 6780
rect 16150 6544 16192 6780
rect 15872 6016 16192 6544
rect 15872 5952 15880 6016
rect 15944 5952 15960 6016
rect 16024 5952 16040 6016
rect 16104 5952 16120 6016
rect 16184 5952 16192 6016
rect 15872 4928 16192 5952
rect 15872 4864 15880 4928
rect 15944 4864 15960 4928
rect 16024 4864 16040 4928
rect 16104 4864 16120 4928
rect 16184 4864 16192 4928
rect 15872 3840 16192 4864
rect 15872 3776 15880 3840
rect 15944 3776 15960 3840
rect 16024 3776 16040 3840
rect 16104 3776 16120 3840
rect 16184 3776 16192 3840
rect 15872 3400 16192 3776
rect 15872 3164 15914 3400
rect 16150 3164 16192 3400
rect 15872 2752 16192 3164
rect 15872 2688 15880 2752
rect 15944 2688 15960 2752
rect 16024 2688 16040 2752
rect 16104 2688 16120 2752
rect 16184 2688 16192 2752
rect 15872 1664 16192 2688
rect 15872 1600 15880 1664
rect 15944 1600 15960 1664
rect 16024 1600 16040 1664
rect 16104 1600 16120 1664
rect 16184 1600 16192 1664
rect 15872 576 16192 1600
rect 15872 512 15880 576
rect 15944 512 15960 576
rect 16024 512 16040 576
rect 16104 512 16120 576
rect 16184 512 16192 576
rect 15872 -48 16192 512
rect 17422 10912 17742 10928
rect 17422 10848 17430 10912
rect 17494 10848 17510 10912
rect 17574 10848 17590 10912
rect 17654 10848 17670 10912
rect 17734 10848 17742 10912
rect 17422 9824 17742 10848
rect 17422 9760 17430 9824
rect 17494 9760 17510 9824
rect 17574 9760 17590 9824
rect 17654 9760 17670 9824
rect 17734 9760 17742 9824
rect 17422 8736 17742 9760
rect 17422 8672 17430 8736
rect 17494 8672 17510 8736
rect 17574 8672 17590 8736
rect 17654 8672 17670 8736
rect 17734 8672 17742 8736
rect 17422 8470 17742 8672
rect 17422 8234 17464 8470
rect 17700 8234 17742 8470
rect 17422 7648 17742 8234
rect 17422 7584 17430 7648
rect 17494 7584 17510 7648
rect 17574 7584 17590 7648
rect 17654 7584 17670 7648
rect 17734 7584 17742 7648
rect 17422 6560 17742 7584
rect 17422 6496 17430 6560
rect 17494 6496 17510 6560
rect 17574 6496 17590 6560
rect 17654 6496 17670 6560
rect 17734 6496 17742 6560
rect 17422 5472 17742 6496
rect 17422 5408 17430 5472
rect 17494 5408 17510 5472
rect 17574 5408 17590 5472
rect 17654 5408 17670 5472
rect 17734 5408 17742 5472
rect 17422 5090 17742 5408
rect 17422 4854 17464 5090
rect 17700 4854 17742 5090
rect 17422 4384 17742 4854
rect 17422 4320 17430 4384
rect 17494 4320 17510 4384
rect 17574 4320 17590 4384
rect 17654 4320 17670 4384
rect 17734 4320 17742 4384
rect 17422 3296 17742 4320
rect 17422 3232 17430 3296
rect 17494 3232 17510 3296
rect 17574 3232 17590 3296
rect 17654 3232 17670 3296
rect 17734 3232 17742 3296
rect 17422 2208 17742 3232
rect 17422 2144 17430 2208
rect 17494 2144 17510 2208
rect 17574 2144 17590 2208
rect 17654 2144 17670 2208
rect 17734 2144 17742 2208
rect 17422 1120 17742 2144
rect 17422 1056 17430 1120
rect 17494 1056 17510 1120
rect 17574 1056 17590 1120
rect 17654 1056 17670 1120
rect 17734 1056 17742 1120
rect 17422 32 17742 1056
rect 17422 -32 17430 32
rect 17494 -32 17510 32
rect 17574 -32 17590 32
rect 17654 -32 17670 32
rect 17734 -32 17742 32
rect 17422 -48 17742 -32
<< via4 >>
rect 3514 9924 3750 10160
rect 3514 6544 3750 6780
rect 3514 3164 3750 3400
rect 5064 8234 5300 8470
rect 5064 4854 5300 5090
rect 6614 9924 6850 10160
rect 6614 6544 6850 6780
rect 6614 3164 6850 3400
rect 8164 8234 8400 8470
rect 8164 4854 8400 5090
rect 9714 9924 9950 10160
rect 9714 6544 9950 6780
rect 9714 3164 9950 3400
rect 11264 8234 11500 8470
rect 11264 4854 11500 5090
rect 12814 9924 13050 10160
rect 12814 6544 13050 6780
rect 12814 3164 13050 3400
rect 14364 8234 14600 8470
rect 14364 4854 14600 5090
rect 15914 9924 16150 10160
rect 15914 6544 16150 6780
rect 15914 3164 16150 3400
rect 17464 8234 17700 8470
rect 17464 4854 17700 5090
<< metal5 >>
rect 368 10160 18860 10202
rect 368 9924 3514 10160
rect 3750 9924 6614 10160
rect 6850 9924 9714 10160
rect 9950 9924 12814 10160
rect 13050 9924 15914 10160
rect 16150 9924 18860 10160
rect 368 9882 18860 9924
rect 368 8470 18860 8512
rect 368 8234 5064 8470
rect 5300 8234 8164 8470
rect 8400 8234 11264 8470
rect 11500 8234 14364 8470
rect 14600 8234 17464 8470
rect 17700 8234 18860 8470
rect 368 8192 18860 8234
rect 368 6780 18860 6822
rect 368 6544 3514 6780
rect 3750 6544 6614 6780
rect 6850 6544 9714 6780
rect 9950 6544 12814 6780
rect 13050 6544 15914 6780
rect 16150 6544 18860 6780
rect 368 6502 18860 6544
rect 368 5090 18860 5132
rect 368 4854 5064 5090
rect 5300 4854 8164 5090
rect 8400 4854 11264 5090
rect 11500 4854 14364 5090
rect 14600 4854 17464 5090
rect 17700 4854 18860 5090
rect 368 4812 18860 4854
rect 368 3400 18860 3442
rect 368 3164 3514 3400
rect 3750 3164 6614 3400
rect 6850 3164 9714 3400
rect 9950 3164 12814 3400
rect 13050 3164 15914 3400
rect 16150 3164 18860 3400
rect 368 3122 18860 3164
use sky130_fd_sc_hd__decap_3  PHY_2 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 368 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1636915332
transform 1 0 368 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 644 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1380 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1564 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_23 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2484 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15
timestamp 1636915332
transform 1 0 1748 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__SET_B OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2576 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 644 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_14
timestamp 1636915332
transform 1 0 1656 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_27
timestamp 1636915332
transform 1 0 2852 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40
timestamp 1636915332
transform 1 0 4048 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48
timestamp 1636915332
transform 1 0 4784 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1636915332
transform 1 0 2760 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1636915332
transform 1 0 3956 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1636915332
transform 1 0 2760 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _335_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 5152 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _336_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 5152 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _441_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 4784 0 -1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__o21ai_1  _333_
timestamp 1636915332
transform -1 0 6072 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _311_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5244 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1636915332
transform 1 0 5152 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1636915332
transform 1 0 5152 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62
timestamp 1636915332
transform 1 0 6072 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56
timestamp 1636915332
transform 1 0 5520 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53
timestamp 1636915332
transform 1 0 5244 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__RESET_B
timestamp 1636915332
transform -1 0 5520 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__nand3_1  _312_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 6440 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1636915332
transform 1 0 6348 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70
timestamp 1636915332
transform 1 0 6808 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtn_1  _442_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5520 0 -1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__xor2_1  _357_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7820 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _356_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8096 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _308_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8096 0 -1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1636915332
transform 1 0 7544 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1636915332
transform 1 0 7544 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_79
timestamp 1636915332
transform 1 0 7636 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_76
timestamp 1636915332
transform 1 0 7360 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79
timestamp 1636915332
transform 1 0 7636 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _382_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9016 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _355_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8832 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1636915332
transform 1 0 8740 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_88
timestamp 1636915332
transform 1 0 8464 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9476 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1636915332
transform 1 0 9936 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1636915332
transform 1 0 9936 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_105
timestamp 1636915332
transform 1 0 10028 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_103
timestamp 1636915332
transform 1 0 9844 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103
timestamp 1636915332
transform 1 0 9844 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__RESET_B
timestamp 1636915332
transform 1 0 10212 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1636915332
transform 1 0 11132 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _453_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10396 0 -1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_0_118
timestamp 1636915332
transform 1 0 11224 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_105
timestamp 1636915332
transform 1 0 10028 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__xor2_1  _361_
timestamp 1636915332
transform 1 0 12420 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1636915332
transform 1 0 12512 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1636915332
transform 1 0 12328 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1636915332
transform 1 0 12328 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_135
timestamp 1636915332
transform 1 0 12788 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_131
timestamp 1636915332
transform 1 0 12420 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_129
timestamp 1636915332
transform 1 0 12236 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _360_
timestamp 1636915332
transform -1 0 13432 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1636915332
transform -1 0 13800 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _290_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 14720 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1636915332
transform 1 0 13248 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1636915332
transform 1 0 13524 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_139
timestamp 1636915332
transform 1 0 13156 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_142
timestamp 1636915332
transform 1 0 13432 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_138
timestamp 1636915332
transform 1 0 13064 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__SET_B
timestamp 1636915332
transform 1 0 13800 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_144
timestamp 1636915332
transform 1 0 13616 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_1  _292_
timestamp 1636915332
transform 1 0 15088 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _291_
timestamp 1636915332
transform 1 0 14812 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1636915332
transform 1 0 14720 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1636915332
transform 1 0 14720 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_157
timestamp 1636915332
transform 1 0 14812 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__RESET_B
timestamp 1636915332
transform -1 0 15088 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1636915332
transform 1 0 15916 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_168
timestamp 1636915332
transform 1 0 15824 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _451_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 15180 0 -1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_0_170
timestamp 1636915332
transform 1 0 16008 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _401_
timestamp 1636915332
transform 1 0 17204 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _359_
timestamp 1636915332
transform 1 0 17204 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1636915332
transform 1 0 17112 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1636915332
transform 1 0 17112 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 18032 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _358_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 18032 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_190
timestamp 1636915332
transform 1 0 17848 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1636915332
transform 1 0 18308 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1636915332
transform -1 0 18860 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1636915332
transform -1 0 18860 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_196
timestamp 1636915332
transform 1 0 18400 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1636915332
transform 1 0 18400 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1636915332
transform 1 0 1380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1636915332
transform 1 0 1656 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_18
timestamp 1636915332
transform 1 0 2024 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1636915332
transform 1 0 644 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1636915332
transform 1 0 368 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1636915332
transform 1 0 1564 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtn_1  _440_
timestamp 1636915332
transform 1 0 2116 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__RESET_B
timestamp 1636915332
transform 1 0 4048 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_42
timestamp 1636915332
transform 1 0 4232 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1636915332
transform 1 0 3956 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1636915332
transform -1 0 5060 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _339_
timestamp 1636915332
transform -1 0 4784 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_51
timestamp 1636915332
transform 1 0 5060 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_63
timestamp 1636915332
transform 1 0 6164 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_72
timestamp 1636915332
transform 1 0 6992 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1636915332
transform 1 0 6348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1636915332
transform -1 0 6992 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _332_
timestamp 1636915332
transform -1 0 6716 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _385_
timestamp 1636915332
transform 1 0 5336 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _407_
timestamp 1636915332
transform 1 0 7084 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_92
timestamp 1636915332
transform 1 0 8832 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_96
timestamp 1636915332
transform 1 0 9200 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1636915332
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _381_
timestamp 1636915332
transform 1 0 9292 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1636915332
transform 1 0 7912 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_2_106
timestamp 1636915332
transform 1 0 10120 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1636915332
transform 1 0 11132 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _287_
timestamp 1636915332
transform -1 0 11592 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _288_
timestamp 1636915332
transform -1 0 11132 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _399_
timestamp 1636915332
transform 1 0 11592 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_131
timestamp 1636915332
transform 1 0 12420 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_142
timestamp 1636915332
transform 1 0 13432 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1636915332
transform 1 0 13524 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _276_
timestamp 1636915332
transform -1 0 13984 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1636915332
transform 1 0 12604 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _452_
timestamp 1636915332
transform 1 0 13984 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__RESET_B
timestamp 1636915332
transform 1 0 16100 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_170
timestamp 1636915332
transform 1 0 16008 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1636915332
transform 1 0 15916 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _427_
timestamp 1636915332
transform 1 0 16284 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1636915332
transform -1 0 18584 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_193
timestamp 1636915332
transform 1 0 18124 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1636915332
transform -1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1636915332
transform 1 0 18308 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1636915332
transform 1 0 368 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _293_
timestamp 1636915332
transform -1 0 2760 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _448_
timestamp 1636915332
transform -1 0 2484 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__RESET_B
timestamp 1636915332
transform 1 0 3772 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_30
timestamp 1636915332
transform 1 0 3128 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_45 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4508 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1636915332
transform 1 0 2760 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1636915332
transform -1 0 4232 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1636915332
transform -1 0 3128 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _296_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 3772 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _334__6
timestamp 1636915332
transform 1 0 4232 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_51
timestamp 1636915332
transform 1 0 5060 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_66
timestamp 1636915332
transform 1 0 6440 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1636915332
transform 1 0 5152 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _331_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5520 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _338_
timestamp 1636915332
transform 1 0 5244 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_83
timestamp 1636915332
transform 1 0 8004 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_94
timestamp 1636915332
transform 1 0 9016 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1636915332
transform 1 0 7544 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _281_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8648 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _286_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8188 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _309_
timestamp 1636915332
transform -1 0 8004 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 9936 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__SET_B
timestamp 1636915332
transform 1 0 11224 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_120
timestamp 1636915332
transform 1 0 11408 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1636915332
transform 1 0 9936 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _282_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 11224 0 -1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_3_128
timestamp 1636915332
transform 1 0 12144 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_131
timestamp 1636915332
transform 1 0 12420 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_147
timestamp 1636915332
transform 1 0 13892 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1636915332
transform 1 0 12328 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _279_
timestamp 1636915332
transform -1 0 13340 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _284_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 13340 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_155
timestamp 1636915332
transform 1 0 14628 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_157
timestamp 1636915332
transform 1 0 14812 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_161
timestamp 1636915332
transform 1 0 15180 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1636915332
transform 1 0 14720 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _289_
timestamp 1636915332
transform -1 0 14628 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1636915332
transform 1 0 16100 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _405_
timestamp 1636915332
transform 1 0 15272 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_180
timestamp 1636915332
transform 1 0 16928 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1636915332
transform -1 0 18860 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1636915332
transform 1 0 17112 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1636915332
transform 1 0 18032 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp 1636915332
transform 1 0 17204 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1636915332
transform 1 0 18308 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_22
timestamp 1636915332
transform 1 0 2392 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1636915332
transform 1 0 644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1636915332
transform 1 0 368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1636915332
transform 1 0 1564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o21bai_4  _295_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2576 0 1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__and2b_1  _302_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1012 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _304_
timestamp 1636915332
transform -1 0 2392 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_49
timestamp 1636915332
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1636915332
transform 1 0 3956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  rebuffer3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 4876 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_62
timestamp 1636915332
transform 1 0 6072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1636915332
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o21bai_1  _315_
timestamp 1636915332
transform -1 0 6992 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _316_
timestamp 1636915332
transform 1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _330_
timestamp 1636915332
transform -1 0 6072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _386_
timestamp 1636915332
transform 1 0 4968 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_88
timestamp 1636915332
transform 1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1636915332
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _306_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 9660 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _397_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8464 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_108
timestamp 1636915332
transform 1 0 10304 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1636915332
transform 1 0 11132 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _349_
timestamp 1636915332
transform 1 0 9660 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__dfstp_1  _454_
timestamp 1636915332
transform -1 0 13156 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer1
timestamp 1636915332
transform -1 0 11132 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__RESET_B
timestamp 1636915332
transform 1 0 13616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1636915332
transform 1 0 13524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _285_
timestamp 1636915332
transform -1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _443_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 13800 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__RESET_B
timestamp 1636915332
transform 1 0 16008 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1636915332
transform 1 0 15916 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _430_
timestamp 1636915332
transform -1 0 18308 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_4_196
timestamp 1636915332
transform 1 0 18400 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1636915332
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1636915332
transform 1 0 18308 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__SET_B
timestamp 1636915332
transform 1 0 2576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1636915332
transform 1 0 368 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _449_
timestamp 1636915332
transform 1 0 644 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp 1636915332
transform 1 0 2852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1636915332
transform 1 0 2760 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1636915332
transform 1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1636915332
transform 1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _300_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 3772 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _303_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3772 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__SET_B
timestamp 1636915332
transform 1 0 6716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_50
timestamp 1636915332
transform 1 0 4968 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_56
timestamp 1636915332
transform 1 0 5520 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_64
timestamp 1636915332
transform 1 0 6256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_68
timestamp 1636915332
transform 1 0 6624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1636915332
transform 1 0 5152 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _299_
timestamp 1636915332
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _314_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 6256 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer4
timestamp 1636915332
transform -1 0 7544 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1636915332
transform 1 0 7544 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _447_
timestamp 1636915332
transform 1 0 7636 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_5_103
timestamp 1636915332
transform 1 0 9844 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_118
timestamp 1636915332
transform 1 0 11224 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1636915332
transform 1 0 9936 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _283_
timestamp 1636915332
transform 1 0 10028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1636915332
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_2  _351_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10396 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_5_131
timestamp 1636915332
transform 1 0 12420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_137
timestamp 1636915332
transform 1 0 12972 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_144
timestamp 1636915332
transform 1 0 13616 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1636915332
transform 1 0 12328 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1636915332
transform 1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _278_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 13064 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_167
timestamp 1636915332
transform 1 0 15732 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1636915332
transform 1 0 14720 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _325_
timestamp 1636915332
transform -1 0 15732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _329_
timestamp 1636915332
transform 1 0 14812 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  split2
timestamp 1636915332
transform 1 0 16284 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_177
timestamp 1636915332
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_181
timestamp 1636915332
transform 1 0 17020 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_183
timestamp 1636915332
transform 1 0 17204 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_195
timestamp 1636915332
transform 1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1636915332
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1636915332
transform 1 0 17112 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _301__4
timestamp 1636915332
transform -1 0 1012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1636915332
transform 1 0 368 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1636915332
transform 1 0 368 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_7
timestamp 1636915332
transform 1 0 1012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1636915332
transform 1 0 644 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1636915332
transform 1 0 1564 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_18
timestamp 1636915332
transform 1 0 2024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 1636915332
transform 1 0 1656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__RESET_B
timestamp 1636915332
transform 1 0 2484 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtn_1  _450_
timestamp 1636915332
transform 1 0 2116 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _446_
timestamp 1636915332
transform 1 0 644 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 1636915332
transform 1 0 2944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1636915332
transform 1 0 2760 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_31
timestamp 1636915332
transform 1 0 3220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_27
timestamp 1636915332
transform 1 0 2852 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_25
timestamp 1636915332
transform 1 0 2668 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  rebuffer10 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _340_
timestamp 1636915332
transform -1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1636915332
transform 1 0 3956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_37
timestamp 1636915332
transform 1 0 3772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _363_
timestamp 1636915332
transform 1 0 4508 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_7_41
timestamp 1636915332
transform 1 0 4140 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_46
timestamp 1636915332
transform 1 0 4600 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__RESET_B
timestamp 1636915332
transform 1 0 4416 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _403_
timestamp 1636915332
transform 1 0 5520 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _313_
timestamp 1636915332
transform -1 0 5520 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1636915332
transform 1 0 5152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1636915332
transform 1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_56
timestamp 1636915332
transform 1 0 5520 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_52
timestamp 1636915332
transform 1 0 5152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1636915332
transform -1 0 7176 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _364_
timestamp 1636915332
transform -1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1636915332
transform 1 0 6348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_69
timestamp 1636915332
transform 1 0 6716 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_64
timestamp 1636915332
transform 1 0 6256 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _362_
timestamp 1636915332
transform -1 0 7544 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _342_
timestamp 1636915332
transform -1 0 8740 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _341_
timestamp 1636915332
transform 1 0 7452 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _305__5
timestamp 1636915332
transform 1 0 7728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1636915332
transform 1 0 7544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_79
timestamp 1636915332
transform 1 0 7636 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1636915332
transform 1 0 8004 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer9
timestamp 1636915332
transform 1 0 8832 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1636915332
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1636915332
transform 1 0 9476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _439_
timestamp 1636915332
transform 1 0 8004 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _411_
timestamp 1636915332
transform 1 0 10212 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _350_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9936 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1636915332
transform 1 0 9936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_105
timestamp 1636915332
transform 1 0 10028 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_111
timestamp 1636915332
transform 1 0 10580 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_103
timestamp 1636915332
transform 1 0 9844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _348_
timestamp 1636915332
transform 1 0 11040 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1636915332
transform 1 0 11132 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_119
timestamp 1636915332
transform 1 0 11316 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_118
timestamp 1636915332
transform 1 0 11224 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _416_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 11316 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__RESET_B
timestamp 1636915332
transform 1 0 12144 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_148
timestamp 1636915332
transform 1 0 13984 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_127
timestamp 1636915332
transform 1 0 12052 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1636915332
transform 1 0 12328 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1636915332
transform 1 0 13524 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _326_
timestamp 1636915332
transform 1 0 13248 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _327_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 12788 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _328_
timestamp 1636915332
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _432_
timestamp 1636915332
transform 1 0 12420 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__or2b_1  _323_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 15548 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1636915332
transform 1 0 14720 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_157
timestamp 1636915332
transform 1 0 14812 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_154
timestamp 1636915332
transform 1 0 14536 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_1  _324_
timestamp 1636915332
transform -1 0 16100 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1636915332
transform 1 0 15916 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_171
timestamp 1636915332
transform 1 0 16100 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_170
timestamp 1636915332
transform 1 0 16008 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_166
timestamp 1636915332
transform 1 0 15640 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__SET_B
timestamp 1636915332
transform 1 0 15732 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_4  _431_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 18308 0 1 3264
box -38 -48 2246 592
use sky130_fd_sc_hd__dfxtp_1  _414_
timestamp 1636915332
transform 1 0 14168 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1636915332
transform 1 0 17112 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_179
timestamp 1636915332
transform 1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_191
timestamp 1636915332
transform 1 0 17940 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_183
timestamp 1636915332
transform 1 0 17204 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1636915332
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1636915332
transform 1 0 18308 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1636915332
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1636915332
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_196
timestamp 1636915332
transform 1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1636915332
transform -1 0 18308 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_14
timestamp 1636915332
transform 1 0 1656 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_18
timestamp 1636915332
transform 1 0 2024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1636915332
transform 1 0 644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1636915332
transform 1 0 368 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1636915332
transform 1 0 1564 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _318_
timestamp 1636915332
transform -1 0 1564 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _445_
timestamp 1636915332
transform 1 0 2116 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1636915332
transform 1 0 3956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_1  _317_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _319_
timestamp 1636915332
transform 1 0 4048 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_53
timestamp 1636915332
transform 1 0 5244 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_59
timestamp 1636915332
transform 1 0 5796 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_63
timestamp 1636915332
transform 1 0 6164 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1636915332
transform 1 0 6348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _321_
timestamp 1636915332
transform 1 0 6440 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1636915332
transform 1 0 5888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__SET_B
timestamp 1636915332
transform 1 0 7820 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_75
timestamp 1636915332
transform 1 0 7268 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_83
timestamp 1636915332
transform 1 0 8004 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_92
timestamp 1636915332
transform 1 0 8832 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1636915332
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__RESET_B
timestamp 1636915332
transform 1 0 9844 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__RESET_B
timestamp 1636915332
transform 1 0 10948 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_100
timestamp 1636915332
transform 1 0 9568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_105
timestamp 1636915332
transform 1 0 10028 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_113
timestamp 1636915332
transform 1 0 10764 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1636915332
transform 1 0 11132 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _429_
timestamp 1636915332
transform -1 0 13064 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_8_138
timestamp 1636915332
transform 1 0 13064 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_142
timestamp 1636915332
transform 1 0 13432 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_144
timestamp 1636915332
transform 1 0 13616 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1636915332
transform 1 0 13524 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _415_
timestamp 1636915332
transform 1 0 14076 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  split5
timestamp 1636915332
transform -1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__SET_B
timestamp 1636915332
transform 1 0 16192 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_165
timestamp 1636915332
transform 1 0 15548 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_170
timestamp 1636915332
transform 1 0 16008 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1636915332
transform 1 0 15916 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_196
timestamp 1636915332
transform 1 0 18400 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1636915332
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1636915332
transform 1 0 18308 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _428_
timestamp 1636915332
transform -1 0 18308 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_9_15
timestamp 1636915332
transform 1 0 1748 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_23
timestamp 1636915332
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1636915332
transform 1 0 644 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1636915332
transform 1 0 368 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__RESET_B
timestamp 1636915332
transform 1 0 3956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1636915332
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_41
timestamp 1636915332
transform 1 0 4140 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_49
timestamp 1636915332
transform 1 0 4876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1636915332
transform 1 0 2760 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__SET_B
timestamp 1636915332
transform 1 0 5428 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1636915332
transform 1 0 5244 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1636915332
transform 1 0 5152 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_2  _444_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5612 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_9_79
timestamp 1636915332
transform 1 0 7636 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_87
timestamp 1636915332
transform 1 0 8372 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_99
timestamp 1636915332
transform 1 0 9476 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1636915332
transform 1 0 7544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _369_
timestamp 1636915332
transform 1 0 8832 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _370_
timestamp 1636915332
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1636915332
transform 1 0 9936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _424_
timestamp 1636915332
transform -1 0 11868 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_pll_clk
timestamp 1636915332
transform 1 0 9568 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__RESET_B
timestamp 1636915332
transform 1 0 12696 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_125
timestamp 1636915332
transform 1 0 11868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_129
timestamp 1636915332
transform 1 0 12236 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_131
timestamp 1636915332
transform 1 0 12420 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1636915332
transform 1 0 12328 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _469_
timestamp 1636915332
transform 1 0 12880 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_9_157
timestamp 1636915332
transform 1 0 14812 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1636915332
transform 1 0 14720 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_2  _268_
timestamp 1636915332
transform 1 0 16192 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _377_
timestamp 1636915332
transform 1 0 15548 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1636915332
transform -1 0 18308 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_183
timestamp 1636915332
transform 1 0 17204 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_191
timestamp 1636915332
transform 1 0 17940 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1636915332
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1636915332
transform 1 0 17112 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1636915332
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1636915332
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_14
timestamp 1636915332
transform 1 0 1656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1636915332
transform 1 0 644 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1636915332
transform 1 0 368 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1636915332
transform 1 0 1564 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtn_1  _460_
timestamp 1636915332
transform 1 0 2024 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__RESET_B
timestamp 1636915332
transform 1 0 4048 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1636915332
transform 1 0 3864 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1636915332
transform 1 0 3956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 1636915332
transform 1 0 4232 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__SET_B
timestamp 1636915332
transform 1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_62
timestamp 1636915332
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1636915332
transform 1 0 6348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _464_
timestamp 1636915332
transform -1 0 8740 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_pll_clk
timestamp 1636915332
transform -1 0 6808 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1636915332
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 10672 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__463__RESET_B
timestamp 1636915332
transform 1 0 10948 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk_A
timestamp 1636915332
transform 1 0 10672 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_114
timestamp 1636915332
transform 1 0 10856 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1636915332
transform 1 0 11132 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _463_
timestamp 1636915332
transform 1 0 11224 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_10_139
timestamp 1636915332
transform 1 0 13156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_147
timestamp 1636915332
transform 1 0 13892 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1636915332
transform 1 0 13524 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _204_
timestamp 1636915332
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1636915332
transform 1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__RESET_B
timestamp 1636915332
transform 1 0 15732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_165
timestamp 1636915332
transform 1 0 15548 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_170
timestamp 1636915332
transform 1 0 16008 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1636915332
transform 1 0 15916 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _373_
timestamp 1636915332
transform 1 0 14904 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _376_
timestamp 1636915332
transform -1 0 16468 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_196
timestamp 1636915332
transform 1 0 18400 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1636915332
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1636915332
transform 1 0 18308 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _470_
timestamp 1636915332
transform 1 0 16468 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__SET_B
timestamp 1636915332
transform 1 0 2576 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1636915332
transform 1 0 368 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _461_
timestamp 1636915332
transform 1 0 644 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__RESET_B
timestamp 1636915332
transform 1 0 4048 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_35
timestamp 1636915332
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_39
timestamp 1636915332
transform 1 0 3956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_42
timestamp 1636915332
transform 1 0 4232 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1636915332
transform 1 0 2760 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _245_
timestamp 1636915332
transform -1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_50
timestamp 1636915332
transform 1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1636915332
transform 1 0 5244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1636915332
transform 1 0 5152 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _228_
timestamp 1636915332
transform -1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _388_
timestamp 1636915332
transform 1 0 6716 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _389_
timestamp 1636915332
transform 1 0 5888 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_79
timestamp 1636915332
transform 1 0 7636 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_87
timestamp 1636915332
transform 1 0 8372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_97
timestamp 1636915332
transform 1 0 9292 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1636915332
transform 1 0 7544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1636915332
transform 1 0 9016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _221_
timestamp 1636915332
transform -1 0 9016 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_103
timestamp 1636915332
transform 1 0 9844 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1636915332
transform 1 0 10028 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1636915332
transform 1 0 10580 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1636915332
transform 1 0 9936 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _233_
timestamp 1636915332
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1636915332
transform 1 0 11408 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_129
timestamp 1636915332
transform 1 0 12236 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_140
timestamp 1636915332
transform 1 0 13248 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_146
timestamp 1636915332
transform 1 0 13800 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1636915332
transform 1 0 12328 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _273_
timestamp 1636915332
transform -1 0 14168 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1636915332
transform 1 0 12420 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__SET_B
timestamp 1636915332
transform 1 0 16100 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_160
timestamp 1636915332
transform 1 0 15088 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_170
timestamp 1636915332
transform 1 0 16008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1636915332
transform 1 0 14720 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1636915332
transform -1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _271_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 14168 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _387_
timestamp 1636915332
transform -1 0 17112 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _410_
timestamp 1636915332
transform 1 0 15180 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1636915332
transform -1 0 18308 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_192
timestamp 1636915332
transform 1 0 18032 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1636915332
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1636915332
transform 1 0 17112 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _206_
timestamp 1636915332
transform 1 0 17204 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1636915332
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_14
timestamp 1636915332
transform 1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_24
timestamp 1636915332
transform 1 0 2576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1636915332
transform 1 0 644 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1636915332
transform 1 0 1012 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1636915332
transform 1 0 368 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1636915332
transform 1 0 1564 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2ai_1  _241_
timestamp 1636915332
transform 1 0 1932 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _242__1
timestamp 1636915332
transform -1 0 1012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _244_
timestamp 1636915332
transform -1 0 1564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_38
timestamp 1636915332
transform 1 0 3864 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1636915332
transform 1 0 3956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _234_
timestamp 1636915332
transform -1 0 3864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1636915332
transform -1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _236_
timestamp 1636915332
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _237_
timestamp 1636915332
transform -1 0 4600 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  rebuffer8
timestamp 1636915332
transform -1 0 4968 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_50
timestamp 1636915332
transform 1 0 4968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_60
timestamp 1636915332
transform 1 0 5888 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_64
timestamp 1636915332
transform 1 0 6256 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1636915332
transform 1 0 6348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1636915332
transform 1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _229_
timestamp 1636915332
transform -1 0 5888 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _371_
timestamp 1636915332
transform 1 0 6440 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_12_88
timestamp 1636915332
transform 1 0 8464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_92
timestamp 1636915332
transform 1 0 8832 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1636915332
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _230_
timestamp 1636915332
transform 1 0 7360 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _231_
timestamp 1636915332
transform 1 0 7728 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _391_
timestamp 1636915332
transform 1 0 9016 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk90_A
timestamp 1636915332
transform -1 0 11408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_103
timestamp 1636915332
transform 1 0 9844 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_116
timestamp 1636915332
transform 1 0 11040 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_120
timestamp 1636915332
transform 1 0 11408 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1636915332
transform 1 0 11132 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _232_
timestamp 1636915332
transform 1 0 10396 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1636915332
transform 1 0 10764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__SET_B
timestamp 1636915332
transform 1 0 13340 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_126
timestamp 1636915332
transform 1 0 11960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_131
timestamp 1636915332
transform 1 0 12420 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_139
timestamp 1636915332
transform 1 0 13156 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1636915332
transform 1 0 13524 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _368_
timestamp 1636915332
transform 1 0 12052 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _455_
timestamp 1636915332
transform 1 0 13616 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_12_165
timestamp 1636915332
transform 1 0 15548 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1636915332
transform 1 0 15916 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1636915332
transform -1 0 15916 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _372_
timestamp 1636915332
transform 1 0 16008 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_196
timestamp 1636915332
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1636915332
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1636915332
transform 1 0 18308 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _468_
timestamp 1636915332
transform 1 0 16376 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1636915332
transform 1 0 368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1636915332
transform 1 0 368 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1636915332
transform 1 0 644 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1636915332
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _254_
timestamp 1636915332
transform -1 0 2852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _240_
timestamp 1636915332
transform 1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1636915332
transform 1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1636915332
transform 1 0 1564 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_21
timestamp 1636915332
transform 1 0 2300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_14
timestamp 1636915332
transform 1 0 1656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtn_1  _462_
timestamp 1636915332
transform 1 0 644 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__and2b_1  _243_
timestamp 1636915332
transform -1 0 3864 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1636915332
transform -1 0 3128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1636915332
transform 1 0 2760 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_27
timestamp 1636915332
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__462__RESET_B
timestamp 1636915332
transform 1 0 3128 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _384_
timestamp 1636915332
transform 1 0 4048 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1636915332
transform 1 0 3680 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1636915332
transform 1 0 3956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_35
timestamp 1636915332
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_38
timestamp 1636915332
transform 1 0 3864 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _255_
timestamp 1636915332
transform -1 0 5428 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _247_
timestamp 1636915332
transform 1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_46
timestamp 1636915332
transform 1 0 4600 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer7
timestamp 1636915332
transform 1 0 6072 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _390_
timestamp 1636915332
transform 1 0 5244 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _225_
timestamp 1636915332
transform 1 0 5796 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _215_
timestamp 1636915332
transform -1 0 5796 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1636915332
transform 1 0 5152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_pll_clk90
timestamp 1636915332
transform -1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _224_
timestamp 1636915332
transform 1 0 7176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _217_
timestamp 1636915332
transform -1 0 7176 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1636915332
transform 1 0 6348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__459__SET_B
timestamp 1636915332
transform 1 0 6164 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_1  _459_
timestamp 1636915332
transform 1 0 6808 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _246__2
timestamp 1636915332
transform -1 0 7912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1636915332
transform 1 0 7544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_86
timestamp 1636915332
transform 1 0 8280 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_82
timestamp 1636915332
transform 1 0 7912 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _392_
timestamp 1636915332
transform 1 0 8372 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _213_
timestamp 1636915332
transform -1 0 9936 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1636915332
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_96
timestamp 1636915332
transform 1 0 9200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_92
timestamp 1636915332
transform 1 0 8832 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_96
timestamp 1636915332
transform 1 0 9200 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk90
timestamp 1636915332
transform -1 0 11132 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__SET_B
timestamp 1636915332
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1636915332
transform 1 0 9936 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1636915332
transform 1 0 11132 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _210_
timestamp 1636915332
transform -1 0 12052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _223_
timestamp 1636915332
transform 1 0 10028 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _226_
timestamp 1636915332
transform -1 0 11132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _227_
timestamp 1636915332
transform 1 0 11132 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _466_
timestamp 1636915332
transform 1 0 11224 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _353_
timestamp 1636915332
transform 1 0 12604 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1636915332
transform 1 0 12328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_131
timestamp 1636915332
transform 1 0 12420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_127
timestamp 1636915332
transform 1 0 12052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_pll_clk90
timestamp 1636915332
transform 1 0 13156 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _272_
timestamp 1636915332
transform -1 0 14444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1636915332
transform 1 0 13616 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1636915332
transform 1 0 13524 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_147
timestamp 1636915332
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_148
timestamp 1636915332
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_140
timestamp 1636915332
transform 1 0 13248 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2ai_2  _354_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 15088 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__RESET_B
timestamp 1636915332
transform 1 0 15088 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__RESET_B
timestamp 1636915332
transform 1 0 16008 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1636915332
transform 1 0 14720 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1636915332
transform 1 0 15916 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1636915332
transform 1 0 14444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _352_
timestamp 1636915332
transform -1 0 15088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _413_
timestamp 1636915332
transform 1 0 15088 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _433_
timestamp 1636915332
transform -1 0 17112 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _436_
timestamp 1636915332
transform 1 0 16192 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_12  FILLER_13_186
timestamp 1636915332
transform 1 0 17480 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_196
timestamp 1636915332
transform 1 0 18400 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1636915332
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1636915332
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1636915332
transform 1 0 17112 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1636915332
transform 1 0 18308 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _207_
timestamp 1636915332
transform 1 0 17204 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__456__RESET_B
timestamp 1636915332
transform 1 0 2484 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1636915332
transform 1 0 368 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _456_
timestamp 1636915332
transform 1 0 644 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_15_25
timestamp 1636915332
transform 1 0 2668 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_49
timestamp 1636915332
transform 1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1636915332
transform 1 0 2760 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _259_
timestamp 1636915332
transform 1 0 3128 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _266_
timestamp 1636915332
transform -1 0 3128 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _383_
timestamp 1636915332
transform -1 0 4876 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_53
timestamp 1636915332
transform 1 0 5244 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_68
timestamp 1636915332
transform 1 0 6624 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1636915332
transform 1 0 5152 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _250_
timestamp 1636915332
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _256_
timestamp 1636915332
transform -1 0 5888 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _257_
timestamp 1636915332
transform -1 0 6624 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__RESET_B
timestamp 1636915332
transform 1 0 8648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_76
timestamp 1636915332
transform 1 0 7360 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_79
timestamp 1636915332
transform 1 0 7636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_83
timestamp 1636915332
transform 1 0 8004 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_87
timestamp 1636915332
transform 1 0 8372 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1636915332
transform 1 0 7544 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _212_
timestamp 1636915332
transform 1 0 8832 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _214_
timestamp 1636915332
transform 1 0 9292 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1636915332
transform -1 0 8372 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_105
timestamp 1636915332
transform 1 0 10028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1636915332
transform 1 0 9936 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _208_
timestamp 1636915332
transform 1 0 10396 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _209_
timestamp 1636915332
transform 1 0 10948 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _211_
timestamp 1636915332
transform -1 0 9936 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _218_
timestamp 1636915332
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_127
timestamp 1636915332
transform 1 0 12052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_131
timestamp 1636915332
transform 1 0 12420 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1636915332
transform 1 0 12328 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _417_
timestamp 1636915332
transform -1 0 14168 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__SET_B
timestamp 1636915332
transform 1 0 14536 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_150
timestamp 1636915332
transform 1 0 14168 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1636915332
transform 1 0 14720 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _434_
timestamp 1636915332
transform 1 0 14812 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__SET_B
timestamp 1636915332
transform 1 0 16744 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1636915332
transform 1 0 18400 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_180
timestamp 1636915332
transform 1 0 16928 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_183
timestamp 1636915332
transform 1 0 17204 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1636915332
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1636915332
transform 1 0 17112 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1636915332
transform 1 0 17756 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  split6
timestamp 1636915332
transform -1 0 18400 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1636915332
transform -1 0 1196 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1636915332
transform 1 0 644 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1636915332
transform 1 0 368 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1636915332
transform 1 0 1564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _267_
timestamp 1636915332
transform -1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  input3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1656 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_16_33
timestamp 1636915332
transform 1 0 3404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_43
timestamp 1636915332
transform 1 0 4324 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1636915332
transform 1 0 3956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _258_
timestamp 1636915332
transform 1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1636915332
transform -1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_55
timestamp 1636915332
transform 1 0 5428 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_63
timestamp 1636915332
transform 1 0 6164 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1636915332
transform 1 0 6348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _409_
timestamp 1636915332
transform 1 0 6440 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1636915332
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _419_
timestamp 1636915332
transform 1 0 7268 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _426_
timestamp 1636915332
transform 1 0 8832 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__RESET_B
timestamp 1636915332
transform 1 0 10948 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_112
timestamp 1636915332
transform 1 0 10672 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1636915332
transform 1 0 11132 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _467_
timestamp 1636915332
transform 1 0 11224 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__RESET_B
timestamp 1636915332
transform 1 0 13892 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1636915332
transform 1 0 13340 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_144
timestamp 1636915332
transform 1 0 13616 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1636915332
transform 1 0 13524 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _435_
timestamp 1636915332
transform 1 0 14076 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1636915332
transform 1 0 15916 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _437_
timestamp 1636915332
transform 1 0 16008 0 1 8704
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_1  FILLER_16_194
timestamp 1636915332
transform 1 0 18216 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_196
timestamp 1636915332
transform 1 0 18400 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1636915332
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1636915332
transform 1 0 18308 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1636915332
transform 1 0 368 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _260_
timestamp 1636915332
transform -1 0 2760 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _458_
timestamp 1636915332
transform 1 0 644 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__SET_B
timestamp 1636915332
transform 1 0 3956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__RESET_B
timestamp 1636915332
transform 1 0 4140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_34
timestamp 1636915332
transform 1 0 3496 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_38
timestamp 1636915332
transform 1 0 3864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1636915332
transform 1 0 2760 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1636915332
transform -1 0 3864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _253_
timestamp 1636915332
transform -1 0 3220 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _263_
timestamp 1636915332
transform -1 0 3496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _396_
timestamp 1636915332
transform 1 0 4324 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_62
timestamp 1636915332
transform 1 0 6072 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_74
timestamp 1636915332
transform 1 0 7176 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1636915332
transform 1 0 5152 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _395_
timestamp 1636915332
transform 1 0 5244 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1636915332
transform -1 0 7176 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_79
timestamp 1636915332
transform 1 0 7636 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_87
timestamp 1636915332
transform 1 0 8372 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1636915332
transform 1 0 7544 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _418_
timestamp 1636915332
transform 1 0 8464 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_105
timestamp 1636915332
transform 1 0 10028 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_109
timestamp 1636915332
transform 1 0 10396 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_119
timestamp 1636915332
transform 1 0 11316 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1636915332
transform 1 0 9936 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _394_
timestamp 1636915332
transform 1 0 11500 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1636915332
transform -1 0 11316 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1636915332
transform 1 0 12328 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _423_
timestamp 1636915332
transform 1 0 12788 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_ext_clk
timestamp 1636915332
transform -1 0 12788 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1636915332
transform 1 0 14720 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _438_
timestamp 1636915332
transform -1 0 16928 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1636915332
transform -1 0 18308 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_180
timestamp 1636915332
transform 1 0 16928 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_183
timestamp 1636915332
transform 1 0 17204 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_191
timestamp 1636915332
transform 1 0 17940 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1636915332
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1636915332
transform 1 0 17112 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1636915332
transform 1 0 18308 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_11
timestamp 1636915332
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1636915332
transform 1 0 644 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1636915332
transform 1 0 368 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1636915332
transform 1 0 1564 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _261_
timestamp 1636915332
transform -1 0 2024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _457_
timestamp 1636915332
transform 1 0 2024 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_18_40
timestamp 1636915332
transform 1 0 4048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1636915332
transform 1 0 3956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_2  _249_
timestamp 1636915332
transform 1 0 4784 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _367_
timestamp 1636915332
transform 1 0 4140 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_18_66
timestamp 1636915332
transform 1 0 6440 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1636915332
transform 1 0 6348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _365_
timestamp 1636915332
transform 1 0 5704 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _420_
timestamp 1636915332
transform 1 0 7176 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_ext_clk_A
timestamp 1636915332
transform 1 0 9108 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_90
timestamp 1636915332
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_92
timestamp 1636915332
transform 1 0 8832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1636915332
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ext_clk
timestamp 1636915332
transform 1 0 9292 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1636915332
transform 1 0 11132 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _425_
timestamp 1636915332
transform 1 0 11224 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__SET_B
timestamp 1636915332
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__SET_B
timestamp 1636915332
transform 1 0 13064 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_140
timestamp 1636915332
transform 1 0 13248 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_144
timestamp 1636915332
transform 1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1636915332
transform 1 0 13524 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _422_
timestamp 1636915332
transform 1 0 13984 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__SET_B
timestamp 1636915332
transform 1 0 16008 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1636915332
transform 1 0 15916 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _421_
timestamp 1636915332
transform 1 0 16192 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_18_193
timestamp 1636915332
transform 1 0 18124 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_196
timestamp 1636915332
transform 1 0 18400 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1636915332
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1636915332
transform 1 0 18308 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1636915332
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_14
timestamp 1636915332
transform 1 0 1656 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_18
timestamp 1636915332
transform 1 0 2024 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1636915332
transform 1 0 644 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1636915332
transform 1 0 368 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1636915332
transform 1 0 1564 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1636915332
transform -1 0 2668 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262__3
timestamp 1636915332
transform -1 0 2392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_25
timestamp 1636915332
transform 1 0 2668 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_31
timestamp 1636915332
transform 1 0 3220 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_40
timestamp 1636915332
transform 1 0 4048 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1636915332
transform 1 0 2760 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1636915332
transform 1 0 3956 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _264_
timestamp 1636915332
transform -1 0 3220 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_56
timestamp 1636915332
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_64
timestamp 1636915332
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_66
timestamp 1636915332
transform 1 0 6440 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1636915332
transform 1 0 5152 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1636915332
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _344_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 6900 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _366_
timestamp 1636915332
transform 1 0 5244 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_ext_clk
timestamp 1636915332
transform 1 0 7176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output10
timestamp 1636915332
transform -1 0 6900 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__S
timestamp 1636915332
transform 1 0 8556 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_79
timestamp 1636915332
transform 1 0 7636 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1636915332
transform 1 0 7544 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1636915332
transform 1 0 8740 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _343_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7728 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8832 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__RESET_B
timestamp 1636915332
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_100
timestamp 1636915332
transform 1 0 9568 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_108
timestamp 1636915332
transform 1 0 10304 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_116
timestamp 1636915332
transform 1 0 11040 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_120
timestamp 1636915332
transform 1 0 11408 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1636915332
transform 1 0 9936 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1636915332
transform 1 0 11132 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  output12
timestamp 1636915332
transform 1 0 10028 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1636915332
transform 1 0 12144 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_140
timestamp 1636915332
transform 1 0 13248 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1636915332
transform 1 0 12328 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1636915332
transform 1 0 13524 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _378__13 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 14260 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _393_
timestamp 1636915332
transform -1 0 13248 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1636915332
transform -1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__RESET_B
timestamp 1636915332
transform 1 0 14812 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_151
timestamp 1636915332
transform 1 0 14260 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_155
timestamp 1636915332
transform 1 0 14628 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1636915332
transform 1 0 14996 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_167
timestamp 1636915332
transform 1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_170
timestamp 1636915332
transform 1 0 16008 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1636915332
transform 1 0 14720 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1636915332
transform 1 0 15916 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1636915332
transform -1 0 18308 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_183
timestamp 1636915332
transform 1 0 17204 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_196
timestamp 1636915332
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1636915332
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1636915332
transform 1 0 17112 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1636915332
transform 1 0 18308 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _375_
timestamp 1636915332
transform -1 0 18124 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1636915332
transform -1 0 17848 0 -1 10880
box -38 -48 314 592
<< labels >>
rlabel metal5 s 368 4812 18860 5132 6 VGND
port 0 nsew ground input
rlabel metal5 s 368 8192 18860 8512 6 VGND
port 0 nsew ground input
rlabel metal4 s 5022 -48 5342 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 8122 -48 8442 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 11222 -48 11542 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 14322 -48 14642 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 17422 -48 17742 10928 6 VGND
port 0 nsew ground input
rlabel metal5 s 368 3122 18860 3442 6 VPWR
port 1 nsew power input
rlabel metal5 s 368 6502 18860 6822 6 VPWR
port 1 nsew power input
rlabel metal5 s 368 9882 18860 10202 6 VPWR
port 1 nsew power input
rlabel metal4 s 3472 -48 3792 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 6572 -48 6892 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 9672 -48 9992 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 12772 -48 13092 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 15872 -48 16192 10928 6 VPWR
port 1 nsew power input
rlabel metal2 s 7102 11200 7158 12000 6 core_clk
port 2 nsew signal tristate
rlabel metal2 s 4250 11200 4306 12000 6 ext_clk
port 3 nsew signal input
rlabel metal3 s 19200 688 20000 808 6 ext_clk_sel
port 4 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 ext_reset
port 5 nsew signal input
rlabel metal2 s 15658 11200 15714 12000 6 pll_clk
port 6 nsew signal input
rlabel metal2 s 18510 11200 18566 12000 6 pll_clk90
port 7 nsew signal input
rlabel metal2 s 1398 11200 1454 12000 6 resetb
port 8 nsew signal input
rlabel metal2 s 12806 11200 12862 12000 6 resetb_sync
port 9 nsew signal tristate
rlabel metal3 s 19200 6672 20000 6792 6 sel2[0]
port 10 nsew signal input
rlabel metal3 s 19200 8168 20000 8288 6 sel2[1]
port 11 nsew signal input
rlabel metal3 s 19200 9664 20000 9784 6 sel2[2]
port 12 nsew signal input
rlabel metal3 s 19200 2184 20000 2304 6 sel[0]
port 13 nsew signal input
rlabel metal3 s 19200 3680 20000 3800 6 sel[1]
port 14 nsew signal input
rlabel metal3 s 19200 5176 20000 5296 6 sel[2]
port 15 nsew signal input
rlabel metal2 s 9954 11200 10010 12000 6 user_clk
port 16 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 12000
<< end >>
