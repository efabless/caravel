magic
tech sky130A
magscale 1 2
timestamp 1684835651
<< metal5 >>
rect 78610 1018624 90778 1030788
rect 130010 1018624 142178 1030788
rect 181410 1018624 193578 1030788
rect 231810 1018624 243978 1030788
rect 284410 1018624 296578 1030788
rect 334810 1018624 346978 1030788
rect 386210 1018624 398378 1030788
rect 475210 1018624 487378 1030788
rect 526610 1018624 538778 1030788
rect 577010 1018624 589178 1030788
rect 628410 1018624 640578 1030788
rect 19178 968893 19501 969216
rect 710938 965293 711261 965616
rect 19821 925053 20141 925373
rect 711581 920653 711901 920973
rect 19178 883493 19501 883816
rect 698230 876147 698523 876440
rect 19178 841293 19501 841616
rect 710938 832093 711261 832416
rect 6316 799147 6609 799440
rect 698230 786947 698523 787240
rect 6316 755947 6609 756240
rect 698230 741947 698523 742240
rect 6316 712747 6609 713040
rect 698230 696947 698523 697240
rect 6316 669547 6609 669840
rect 698230 651747 698523 652040
rect 6316 626347 6609 626640
rect 698230 606747 698523 607040
rect 6316 583147 6609 583440
rect 698230 561547 698523 561840
rect 6316 539947 6609 540240
rect 710938 517493 711261 517816
rect 19178 496693 19501 497016
rect 711581 472853 711901 473173
rect 19821 453853 20141 454173
rect 710938 429293 711261 429616
rect 6316 412347 6609 412640
rect 698230 384347 698523 384640
rect 6316 369147 6609 369440
rect 698230 339147 698523 339440
rect 6316 325947 6609 326240
rect 698230 294147 698523 294440
rect 6316 282747 6609 283040
rect 698230 249147 698523 249440
rect 6316 239547 6609 239840
rect 698230 203947 698523 204240
rect 6316 196347 6609 196640
rect 698230 158947 698523 159240
rect 19178 123893 19501 124216
rect 698230 113747 698523 114040
rect 19821 81053 20141 81373
rect 254320 19754 254640 20074
rect 187371 19088 187694 19411
rect 295971 19088 296294 19411
rect 350771 19088 351094 19411
rect 405571 19088 405894 19411
rect 460371 19088 460694 19411
rect 515171 19088 515494 19411
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use caravel_logo  caravel_logo
timestamp 0
transform 1 0 216000 0 1 5100
box 0 0 1 1
use caravel_motto  caravel_motto
timestamp 0
transform 1 0 270000 0 1 -7000
box 0 0 1 1
use caravan_core  chip_core
timestamp 0
transform 1 0 42300 0 1 42100
box 0 0 1 1
use copyright_block  copyright_block
timestamp 0
transform 1 0 96400 0 1 17000
box 0 0 1 1
use open_source  open_source
timestamp 0
transform 1 0 153600 0 1 3000
box 0 0 1 1
use chip_io_alt  padframe
timestamp 0
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use user_id_textblock  user_id_textblock
timestamp 0
transform 1 0 35000 0 1 7000
box 0 0 1 1
<< labels >>
flabel metal5 s 187371 19088 187694 19411 0 FreeSans 2560 0 0 0 clock
port 0 nsew signal input
flabel metal5 s 350771 19088 351094 19411 0 FreeSans 2560 0 0 0 flash_clk
port 1 nsew signal tristate
flabel metal5 s 295971 19088 296294 19411 0 FreeSans 2560 0 0 0 flash_csb
port 2 nsew signal tristate
flabel metal5 s 405571 19088 405894 19411 0 FreeSans 2560 0 0 0 flash_io0
port 3 nsew signal tristate
flabel metal5 s 460371 19088 460694 19411 0 FreeSans 2560 0 0 0 flash_io1
port 4 nsew signal tristate
flabel metal5 s 515171 19088 515494 19411 0 FreeSans 2560 0 0 0 gpio
port 5 nsew signal bidirectional
flabel metal5 s 698230 113747 698523 114040 0 FreeSans 2560 0 0 0 mprj_io[0]
port 6 nsew signal bidirectional
flabel metal5 s 698230 696947 698523 697240 0 FreeSans 2560 0 0 0 mprj_io[10]
port 7 nsew signal bidirectional
flabel metal5 s 698230 741947 698523 742240 0 FreeSans 2560 0 0 0 mprj_io[11]
port 8 nsew signal bidirectional
flabel metal5 s 698230 786947 698523 787240 0 FreeSans 2560 0 0 0 mprj_io[12]
port 9 nsew signal bidirectional
flabel metal5 s 698230 876147 698523 876440 0 FreeSans 2560 0 0 0 mprj_io[13]
port 10 nsew signal bidirectional
flabel metal5 s 710938 965293 711261 965616 0 FreeSans 2560 0 0 0 mprj_io[14]
port 11 nsew signal bidirectional
flabel metal5 s 628410 1018624 640578 1030788 0 FreeSans 81920 0 0 0 mprj_io[15]
port 12 nsew signal bidirectional
flabel metal5 s 526610 1018624 538778 1030788 0 FreeSans 81920 0 0 0 mprj_io[16]
port 13 nsew signal bidirectional
flabel metal5 s 475210 1018624 487378 1030788 0 FreeSans 81920 0 0 0 mprj_io[17]
port 14 nsew signal bidirectional
flabel metal5 s 386210 1018624 398378 1030788 0 FreeSans 81920 0 0 0 mprj_io[18]
port 15 nsew signal bidirectional
flabel metal5 s 284410 1018624 296578 1030788 0 FreeSans 81920 0 0 0 mprj_io[19]
port 16 nsew signal bidirectional
flabel metal5 s 698230 158947 698523 159240 0 FreeSans 2560 0 0 0 mprj_io[1]
port 17 nsew signal bidirectional
flabel metal5 s 231810 1018624 243978 1030788 0 FreeSans 81920 0 0 0 mprj_io[20]
port 18 nsew signal bidirectional
flabel metal5 s 181410 1018624 193578 1030788 0 FreeSans 81920 0 0 0 mprj_io[21]
port 19 nsew signal bidirectional
flabel metal5 s 130010 1018624 142178 1030788 0 FreeSans 81920 0 0 0 mprj_io[22]
port 20 nsew signal bidirectional
flabel metal5 s 78610 1018624 90778 1030788 0 FreeSans 81920 0 0 0 mprj_io[23]
port 21 nsew signal bidirectional
flabel metal5 s 19178 968893 19501 969216 0 FreeSans 2560 0 0 0 mprj_io[24]
port 22 nsew signal bidirectional
flabel metal5 s 6316 799147 6609 799440 0 FreeSans 2560 0 0 0 mprj_io[25]
port 23 nsew signal bidirectional
flabel metal5 s 6316 755947 6609 756240 0 FreeSans 2560 0 0 0 mprj_io[26]
port 24 nsew signal bidirectional
flabel metal5 s 6316 712747 6609 713040 0 FreeSans 2560 0 0 0 mprj_io[27]
port 25 nsew signal bidirectional
flabel metal5 s 6316 669547 6609 669840 0 FreeSans 2560 0 0 0 mprj_io[28]
port 26 nsew signal bidirectional
flabel metal5 s 6316 626347 6609 626640 0 FreeSans 2560 0 0 0 mprj_io[29]
port 27 nsew signal bidirectional
flabel metal5 s 698230 203947 698523 204240 0 FreeSans 2560 0 0 0 mprj_io[2]
port 28 nsew signal bidirectional
flabel metal5 s 6316 583147 6609 583440 0 FreeSans 2560 0 0 0 mprj_io[30]
port 29 nsew signal bidirectional
flabel metal5 s 6316 539947 6609 540240 0 FreeSans 2560 0 0 0 mprj_io[31]
port 30 nsew signal bidirectional
flabel metal5 s 6316 412347 6609 412640 0 FreeSans 2560 0 0 0 mprj_io[32]
port 31 nsew signal bidirectional
flabel metal5 s 6316 369147 6609 369440 0 FreeSans 2560 0 0 0 mprj_io[33]
port 32 nsew signal bidirectional
flabel metal5 s 6316 325947 6609 326240 0 FreeSans 2560 0 0 0 mprj_io[34]
port 33 nsew signal bidirectional
flabel metal5 s 6316 282747 6609 283040 0 FreeSans 2560 0 0 0 mprj_io[35]
port 34 nsew signal bidirectional
flabel metal5 s 6316 239547 6609 239840 0 FreeSans 2560 0 0 0 mprj_io[36]
port 35 nsew signal bidirectional
flabel metal5 s 6316 196347 6609 196640 0 FreeSans 2560 0 0 0 mprj_io[37]
port 36 nsew signal bidirectional
flabel metal5 s 698230 249147 698523 249440 0 FreeSans 2560 0 0 0 mprj_io[3]
port 37 nsew signal bidirectional
flabel metal5 s 698230 294147 698523 294440 0 FreeSans 2560 0 0 0 mprj_io[4]
port 38 nsew signal bidirectional
flabel metal5 s 698230 339147 698523 339440 0 FreeSans 2560 0 0 0 mprj_io[5]
port 39 nsew signal bidirectional
flabel metal5 s 698230 384347 698523 384640 0 FreeSans 2560 0 0 0 mprj_io[6]
port 40 nsew signal bidirectional
flabel metal5 s 698230 561547 698523 561840 0 FreeSans 2560 0 0 0 mprj_io[7]
port 41 nsew signal bidirectional
flabel metal5 s 698230 606747 698523 607040 0 FreeSans 2560 0 0 0 mprj_io[8]
port 42 nsew signal bidirectional
flabel metal5 s 698230 651747 698523 652040 0 FreeSans 2560 0 0 0 mprj_io[9]
port 43 nsew signal bidirectional
flabel metal5 s 136713 7143 144149 18309 0 FreeSans 81920 0 0 0 resetb
port 44 nsew signal input
flabel metal5 s 19821 81053 20141 81373 0 FreeSans 2560 0 0 0 vccd
port 45 nsew signal bidirectional
flabel metal5 s 711581 920653 711901 920973 0 FreeSans 2560 0 0 0 vccd1
port 46 nsew signal bidirectional
flabel metal5 s 19821 925053 20141 925373 0 FreeSans 2560 0 0 0 vccd2
port 47 nsew signal bidirectional
flabel metal5 s 624222 6811 636390 18975 0 FreeSans 81920 0 0 0 vdda
port 48 nsew signal bidirectional
flabel metal5 s 710938 832093 711261 832416 0 FreeSans 2560 0 0 0 vdda1
port 49 nsew signal bidirectional
flabel metal5 s 710938 517493 711261 517816 0 FreeSans 2560 0 0 0 vdda1_2
port 50 nsew signal bidirectional
flabel metal5 s 19178 496693 19501 497016 0 FreeSans 2560 0 0 0 vdda2
port 51 nsew signal bidirectional
flabel metal5 s 19178 123893 19501 124216 0 FreeSans 2560 0 0 0 vddio
port 52 nsew signal bidirectional
flabel metal5 s 19178 883493 19501 883816 0 FreeSans 2560 0 0 0 vddio_2
port 53 nsew signal bidirectional
flabel metal5 s 80222 6811 92390 18975 0 FreeSans 81920 0 0 0 vssa
port 54 nsew signal bidirectional
flabel metal5 s 577010 1018624 589178 1030788 0 FreeSans 81920 0 0 0 vssa1
port 55 nsew signal bidirectional
flabel metal5 s 710938 429293 711261 429616 0 FreeSans 2560 0 0 0 vssa1_2
port 56 nsew signal bidirectional
flabel metal5 s 19178 841293 19501 841616 0 FreeSans 2560 0 0 0 vssa2
port 57 nsew signal bidirectional
flabel metal5 s 254320 19754 254640 20074 0 FreeSans 2560 0 0 0 vssd
port 58 nsew signal bidirectional
flabel metal5 s 711581 472853 711901 473173 0 FreeSans 2560 0 0 0 vssd1
port 59 nsew signal bidirectional
flabel metal5 s 19821 453853 20141 454173 0 FreeSans 2560 0 0 0 vssd2
port 60 nsew signal bidirectional
flabel metal5 s 570422 6811 582590 18975 0 FreeSans 81920 0 0 0 vssio
port 61 nsew signal bidirectional
flabel metal5 s 334810 1018624 346978 1030788 0 FreeSans 81920 0 0 0 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
