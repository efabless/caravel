magic
tech sky130A
timestamp 1638586442
<< metal5 >>
tri 2970 7740 3060 7830 se
rect 3060 7740 3960 8010
tri 3960 7740 4050 7830 sw
tri 2880 7470 2970 7560 se
rect 2970 7470 4050 7740
tri 4050 7470 4140 7560 sw
tri 1440 7291 1619 7470 se
tri 1619 7380 1709 7470 sw
rect 1619 7291 1799 7380
rect 1440 7290 1799 7291
tri 1799 7290 1889 7380 sw
rect 2880 7290 4140 7470
tri 5311 7380 5401 7470 se
tri 5131 7290 5221 7380 se
rect 5221 7291 5401 7380
tri 5401 7291 5580 7470 sw
rect 5221 7290 5580 7291
tri 1080 6930 1440 7290 se
rect 1440 7200 1979 7290
tri 1979 7200 2069 7290 sw
rect 1440 7020 2159 7200
tri 2159 7020 2339 7200 sw
tri 2609 7110 2789 7290 se
rect 2789 7110 4231 7290
tri 4231 7110 4411 7290 sw
tri 4951 7200 5041 7290 se
rect 5041 7200 5580 7290
tri 2339 7020 2429 7110 se
rect 2429 7020 4591 7110
tri 4591 7020 4681 7110 sw
tri 4681 7020 4861 7200 se
rect 4861 7020 5580 7200
rect 1440 6930 5580 7020
tri 5580 6930 5940 7290 sw
tri 1080 6750 1260 6930 ne
rect 1260 6660 5760 6930
tri 5760 6750 5940 6930 nw
tri 1260 6390 1530 6660 ne
tri 1440 6030 1530 6120 se
rect 1530 6030 5490 6660
tri 5490 6390 5760 6660 nw
tri 5490 6030 5580 6120 sw
rect 7056 6101 7356 6161
rect 7776 6101 8076 6161
rect 8436 6101 8856 6161
rect 9096 6101 9516 6161
rect 10296 6101 10716 6161
rect 11016 6101 11316 6161
rect 6996 6041 7416 6101
rect 7716 6041 8136 6101
rect 1440 5940 3240 6030
tri 3240 5940 3330 6030 nw
tri 3690 5940 3780 6030 ne
rect 3780 5940 5580 6030
tri 1260 5670 1440 5850 se
rect 1440 5670 2700 5940
tri 810 5580 900 5670 se
rect 900 5580 2700 5670
rect 540 4770 2700 5580
tri 2700 5490 3150 5940 nw
tri 3870 5490 4320 5940 ne
rect 4320 5670 5580 5940
rect 6936 5921 7476 6041
tri 5580 5670 5760 5850 sw
rect 4320 5580 6120 5670
tri 6120 5580 6210 5670 sw
rect 4320 4770 6480 5580
rect 6936 5501 7116 5921
rect 7296 5501 7476 5921
rect 6936 5381 7476 5501
rect 7656 5921 8196 6041
rect 7656 5501 7836 5921
rect 8016 5501 8196 5921
rect 7656 5381 8196 5501
rect 8376 5981 8916 6101
rect 8376 5801 8556 5981
rect 8736 5801 8916 5981
rect 8376 5681 8916 5801
rect 9096 6041 9576 6101
rect 10236 6041 10716 6101
rect 10956 6041 11376 6101
rect 9096 5921 9636 6041
rect 8376 5621 8856 5681
rect 8376 5441 8556 5621
rect 6996 5321 7416 5381
rect 7656 5321 8136 5381
rect 8376 5321 8916 5441
rect 7056 5261 7356 5321
rect 7656 5261 8076 5321
rect 8436 5261 8916 5321
rect 9096 5261 9276 5921
rect 9456 5261 9636 5921
rect 10176 5981 10716 6041
rect 10176 5801 10416 5981
rect 10896 5921 11436 6041
rect 10176 5741 10596 5801
rect 10236 5681 10656 5741
rect 10296 5621 10716 5681
rect 10476 5441 10716 5621
rect 10176 5381 10716 5441
rect 10896 5501 11076 5921
rect 11256 5501 11436 5921
rect 10896 5381 11436 5501
rect 11616 5501 11796 6161
rect 11976 5501 12156 6161
rect 11616 5381 12156 5501
rect 12336 6101 12756 6161
rect 13176 6101 13476 6161
rect 13836 6101 14256 6161
rect 12336 6041 12816 6101
rect 13116 6041 13536 6101
rect 12336 5921 12876 6041
rect 10176 5321 10656 5381
rect 10956 5321 11376 5381
rect 11676 5321 12096 5381
rect 10176 5261 10596 5321
rect 11016 5261 11316 5321
rect 11736 5261 12036 5321
rect 12336 5261 12516 5921
rect 12696 5801 12876 5921
rect 13056 5921 13596 6041
rect 13056 5501 13236 5921
rect 13416 5801 13596 5921
rect 13776 5981 14316 6101
rect 13776 5801 13956 5981
rect 14136 5801 14316 5981
rect 13776 5681 14316 5801
rect 13776 5621 14256 5681
rect 13416 5501 13596 5621
rect 13056 5381 13596 5501
rect 13776 5441 13956 5621
rect 13116 5321 13536 5381
rect 13776 5321 14316 5441
rect 13176 5261 13476 5321
rect 13836 5261 14316 5321
rect 7656 4901 7836 5261
rect 10176 4901 10356 5261
rect 7656 4841 8076 4901
rect 8376 4841 8856 4901
rect 9096 4841 9516 4901
rect 9936 4841 10356 4901
rect 7656 4781 8136 4841
tri 810 4680 900 4770 ne
rect 900 4680 2700 4770
tri 1170 4500 1350 4680 ne
rect 1350 4410 2700 4680
tri 2700 4410 3060 4770 sw
rect 1350 4320 3060 4410
tri 1350 4230 1440 4320 ne
rect 1440 4230 3060 4320
rect 1440 4140 2970 4230
tri 2970 4140 3060 4230 nw
tri 3960 4410 4320 4770 se
rect 4320 4680 6120 4770
tri 6120 4680 6210 4770 nw
rect 4320 4410 5670 4680
tri 5670 4500 5850 4680 nw
rect 7656 4661 8196 4781
rect 8376 4721 8916 4841
rect 3960 4320 5670 4410
rect 3960 4230 5580 4320
tri 5580 4230 5670 4320 nw
tri 3960 4140 4050 4230 ne
rect 4050 4140 5580 4230
tri 1440 4050 1530 4140 ne
tri 1440 3960 1530 4050 se
rect 1530 3960 2970 4140
tri 1260 3690 1440 3870 se
rect 1440 3780 2880 3960
tri 2880 3870 2970 3960 nw
rect 4050 3960 5490 4140
tri 5490 4050 5580 4140 nw
tri 5490 3960 5580 4050 sw
rect 7656 4001 7836 4661
rect 8016 4001 8196 4661
rect 8736 4541 8916 4721
rect 8376 4361 8916 4541
rect 8376 4181 8556 4361
rect 8736 4181 8916 4361
rect 8376 4061 8916 4181
rect 8436 4001 8916 4061
rect 9096 4781 9576 4841
rect 9876 4781 10356 4841
rect 9096 4661 9636 4781
rect 9096 4001 9276 4661
rect 9456 4541 9636 4661
rect 9816 4661 10356 4781
rect 9816 4241 9996 4661
rect 10176 4241 10356 4661
rect 9816 4121 10356 4241
rect 10536 4241 10716 4901
rect 10896 4241 11076 4901
rect 11256 4241 11436 4901
rect 11616 4841 12096 4901
rect 12336 4841 12756 4901
rect 13116 4841 13536 4901
rect 11616 4721 12156 4841
rect 11976 4541 12156 4721
rect 11676 4481 12156 4541
rect 10536 4121 11436 4241
rect 11616 4361 12156 4481
rect 11616 4181 11796 4361
rect 11976 4181 12156 4361
rect 9876 4061 10356 4121
rect 10596 4061 11376 4121
rect 11616 4061 12156 4181
rect 9936 4001 10356 4061
rect 10656 4001 10896 4061
rect 11076 4001 11316 4061
rect 11676 4001 12156 4061
rect 12336 4781 12816 4841
rect 12336 4661 12876 4781
rect 12336 4001 12516 4661
rect 12696 4541 12876 4661
rect 13056 4721 13596 4841
rect 13056 4541 13236 4721
rect 13416 4541 13596 4721
rect 13056 4361 13596 4541
rect 13056 4181 13236 4361
rect 13056 4061 13596 4181
rect 13116 4001 13596 4061
tri 4050 3870 4140 3960 ne
rect 1440 3690 2790 3780
tri 2790 3690 2880 3780 nw
rect 4140 3780 5580 3960
tri 4140 3690 4230 3780 ne
rect 4230 3690 5580 3780
tri 5580 3690 5760 3870 sw
tri 1080 3420 1260 3600 se
rect 1260 3510 2790 3690
rect 1260 3420 2700 3510
tri 2700 3420 2790 3510 nw
rect 4230 3510 5760 3690
tri 4230 3420 4320 3510 ne
rect 4320 3420 5760 3510
tri 5760 3420 5940 3600 sw
tri 1080 2880 1620 3420 ne
rect 1620 3330 2700 3420
rect 1620 3240 2634 3330
tri 2634 3264 2700 3330 nw
rect 4320 3330 5400 3420
tri 4320 3264 4386 3330 ne
rect 1620 3150 2160 3240
tri 2160 3150 2250 3240 nw
rect 1620 3060 1980 3150
tri 1980 3060 2070 3150 nw
tri 2315 3060 2495 3240 ne
rect 2495 3174 2634 3240
rect 2495 3060 2520 3174
tri 2520 3060 2634 3174 nw
rect 4386 3240 5400 3330
rect 4386 3174 4525 3240
tri 4386 3060 4500 3174 ne
rect 4500 3060 4525 3174
tri 4525 3060 4705 3240 nw
tri 4770 3150 4860 3240 ne
rect 4860 3150 5400 3240
tri 4950 3060 5040 3150 ne
rect 5040 3060 5400 3150
rect 1620 2880 1710 3060
tri 1710 2880 1890 3060 nw
tri 5130 2880 5310 3060 ne
rect 5310 2880 5400 3060
tri 5400 2880 5940 3420 nw
<< fillblock >>
rect 376 2582 6603 8121
rect 6796 3824 14515 6352
<< end >>
