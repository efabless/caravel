* NGSPICE file created from mgmt_protect.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_8 abstract view
.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_2 abstract view
.subckt sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_4 abstract view
.subckt sky130_fd_sc_hd__einvp_4 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for mprj2_logic_high abstract view
.subckt mprj2_logic_high HI vccd2 vssd2
.ends

* Black-box entry subcircuit for mprj_logic_high abstract view
.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[287] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295]
+ HI[296] HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304]
+ HI[305] HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314]
+ HI[315] HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334]
+ HI[335] HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344]
+ HI[345] HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354]
+ HI[355] HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374]
+ HI[375] HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384]
+ HI[385] HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394]
+ HI[395] HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403]
+ HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413]
+ HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423]
+ HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[42] HI[430] HI[431] HI[432] HI[433]
+ HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443]
+ HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453]
+ HI[454] HI[455] HI[456] HI[457] HI[458] HI[459] HI[45] HI[460] HI[461] HI[462] HI[46]
+ HI[47] HI[48] HI[49] HI[4] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57]
+ HI[58] HI[59] HI[5] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68]
+ HI[69] HI[6] HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79]
+ HI[7] HI[80] HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8]
+ HI[90] HI[91] HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1
+ vssd1
.ends

* Black-box entry subcircuit for mgmt_protect_hv abstract view
.subckt mgmt_protect_hv mprj2_vdd_logic1 mprj_vdd_logic1 vccd vssd vdda1 vssa1 vdda2
+ vssa2
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102]
+ la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107]
+ la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[10] la_iena_mprj[110] la_iena_mprj[111]
+ la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116]
+ la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[11] la_iena_mprj[120]
+ la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125]
+ la_iena_mprj[126] la_iena_mprj[127] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14]
+ la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19]
+ la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23]
+ la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28]
+ la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32]
+ la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37]
+ la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3] la_iena_mprj[40] la_iena_mprj[41]
+ la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46]
+ la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[4] la_iena_mprj[50]
+ la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55]
+ la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[5]
+ la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64]
+ la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69]
+ la_iena_mprj[6] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73]
+ la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78]
+ la_iena_mprj[79] la_iena_mprj[7] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82]
+ la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87]
+ la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[8] la_iena_mprj[90] la_iena_mprj[91]
+ la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96]
+ la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[9] la_oenb_core[0]
+ la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104]
+ la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109]
+ la_oenb_core[10] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113]
+ la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118]
+ la_oenb_core[119] la_oenb_core[11] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122]
+ la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127]
+ la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16]
+ la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[1] la_oenb_core[20]
+ la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25]
+ la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[2]
+ la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34]
+ la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39]
+ la_oenb_core[3] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43]
+ la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48]
+ la_oenb_core[49] la_oenb_core[4] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52]
+ la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57]
+ la_oenb_core[58] la_oenb_core[59] la_oenb_core[5] la_oenb_core[60] la_oenb_core[61]
+ la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66]
+ la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[6] la_oenb_core[70]
+ la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75]
+ la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[7]
+ la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84]
+ la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89]
+ la_oenb_core[8] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93]
+ la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98]
+ la_oenb_core[99] la_oenb_core[9] la_oenb_mprj[0] la_oenb_mprj[100] la_oenb_mprj[101]
+ la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106]
+ la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[10] la_oenb_mprj[110]
+ la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115]
+ la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[11]
+ la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124]
+ la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] la_oenb_mprj[12] la_oenb_mprj[13]
+ la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18]
+ la_oenb_mprj[19] la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22]
+ la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27]
+ la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31]
+ la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36]
+ la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40]
+ la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45]
+ la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4]
+ la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54]
+ la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59]
+ la_oenb_mprj[5] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63]
+ la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68]
+ la_oenb_mprj[69] la_oenb_mprj[6] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72]
+ la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77]
+ la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[7] la_oenb_mprj[80] la_oenb_mprj[81]
+ la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86]
+ la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[8] la_oenb_mprj[90]
+ la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95]
+ la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[9]
+ mprj_ack_i_core mprj_ack_i_user mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11]
+ mprj_adr_o_core[12] mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15]
+ mprj_adr_o_core[16] mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19]
+ mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23]
+ mprj_adr_o_core[24] mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27]
+ mprj_adr_o_core[28] mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31]
+ mprj_adr_o_core[3] mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7]
+ mprj_adr_o_core[8] mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11]
+ mprj_adr_o_user[12] mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15]
+ mprj_adr_o_user[16] mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19]
+ mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23]
+ mprj_adr_o_user[24] mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27]
+ mprj_adr_o_user[28] mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31]
+ mprj_adr_o_user[3] mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7]
+ mprj_adr_o_user[8] mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0]
+ mprj_dat_i_core[10] mprj_dat_i_core[11] mprj_dat_i_core[12] mprj_dat_i_core[13]
+ mprj_dat_i_core[14] mprj_dat_i_core[15] mprj_dat_i_core[16] mprj_dat_i_core[17]
+ mprj_dat_i_core[18] mprj_dat_i_core[19] mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21]
+ mprj_dat_i_core[22] mprj_dat_i_core[23] mprj_dat_i_core[24] mprj_dat_i_core[25]
+ mprj_dat_i_core[26] mprj_dat_i_core[27] mprj_dat_i_core[28] mprj_dat_i_core[29]
+ mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31] mprj_dat_i_core[3] mprj_dat_i_core[4]
+ mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7] mprj_dat_i_core[8] mprj_dat_i_core[9]
+ mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11] mprj_dat_i_user[12] mprj_dat_i_user[13]
+ mprj_dat_i_user[14] mprj_dat_i_user[15] mprj_dat_i_user[16] mprj_dat_i_user[17]
+ mprj_dat_i_user[18] mprj_dat_i_user[19] mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21]
+ mprj_dat_i_user[22] mprj_dat_i_user[23] mprj_dat_i_user[24] mprj_dat_i_user[25]
+ mprj_dat_i_user[26] mprj_dat_i_user[27] mprj_dat_i_user[28] mprj_dat_i_user[29]
+ mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31] mprj_dat_i_user[3] mprj_dat_i_user[4]
+ mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7] mprj_dat_i_user[8] mprj_dat_i_user[9]
+ mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13]
+ mprj_dat_o_core[14] mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17]
+ mprj_dat_o_core[18] mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21]
+ mprj_dat_o_core[22] mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25]
+ mprj_dat_o_core[26] mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29]
+ mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4]
+ mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9]
+ mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13]
+ mprj_dat_o_user[14] mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17]
+ mprj_dat_o_user[18] mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21]
+ mprj_dat_o_user[22] mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25]
+ mprj_dat_o_user[26] mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29]
+ mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4]
+ mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9]
+ mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2] mprj_sel_o_core[3]
+ mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3] mprj_stb_o_core
+ mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood user1_vdd_powergood
+ user2_vcc_powergood user2_vdd_powergood user_clock user_clock2 user_irq[0] user_irq[1]
+ user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2] user_irq_ena[0] user_irq_ena[1]
+ user_irq_ena[2] user_reset vccd vccd1 vccd2 vssd vssd1 vssd2 vccd2_uq0 vccd2_uq1
+ vccd2_uq2 vccd2_uq3 vccd2_uq4 vccd2_uq5 vccd2_uq6 vccd1_uq0 vccd1_uq1 vccd1_uq2
+ vccd1_uq3 vccd1_uq4 vccd1_uq5 vssd2_uq0 vssd2_uq1 vssd2_uq2 vssd2_uq3 vssd2_uq4
+ vssd2_uq5 vssd1_uq0 vssd1_uq1 vssd1_uq2 vssd1_uq4 vdda2_uq0 vdda1_uq0
XTAP_177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_29 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[34\]_A input59/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[72\] input357/X mprj_logic_high_inst/HI[402] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[72\]/B sky130_fd_sc_hd__and2_1
XFILLER_4_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input127_A la_data_out_core[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[50\] _642_/A la_buf_enable\[50\]/B vssd vssd vccd vccd la_buf\[50\]/TE
+ sky130_fd_sc_hd__and2b_1
X_501_ _501_/A vssd vssd vccd vccd _501_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_432_ _432_/A vssd vssd vccd vccd _432_/Y sky130_fd_sc_hd__inv_6
XTAP_1844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_363_ _363_/A vssd vssd vccd vccd _363_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input496_A la_oenb_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input92_A la_data_out_core[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[36\] _500_/Y la_buf\[36\]/TE vssd vssd vccd vccd output684/A sky130_fd_sc_hd__einvp_8
XFILLER_6_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[108\] input269/X mprj_logic_high_inst/HI[438] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[108\]/B sky130_fd_sc_hd__and2_1
Xuser_wb_dat_gates\[8\] input580/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[8\]/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_10_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[25\]_A input49/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_45 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output882_A output882/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[25\] input49/X user_to_mprj_in_gates\[25\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[25\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[16\]_A input39/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[100\]_A input5/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output1077_A output1077/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[76\] _339_/Y mprj_logic_high_inst/HI[278] vssd vssd vccd
+ vccd output984/A sky130_fd_sc_hd__einvp_2
XFILLER_2_346 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput990 output990/A vssd vssd vccd vccd la_oenb_core[81] sky130_fd_sc_hd__buf_2
Xla_buf_enable\[98\] _361_/A la_buf_enable\[98\]/B vssd vssd vccd vccd la_buf\[98\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[24\] _456_/Y mprj_dat_buf\[24\]/TE vssd vssd vccd vccd output1093/A
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input244_A la_data_out_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[104\]_TE mprj_logic_high_inst/HI[306] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input411_A la_oenb_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input509_A la_oenb_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_415_ _415_/A vssd vssd vccd vccd _415_/Y sky130_fd_sc_hd__inv_12
XTAP_1696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_346_ _346_/A vssd vssd vccd vccd _346_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput1106 output1106/A vssd vssd vccd vccd mprj_dat_o_user[7] sky130_fd_sc_hd__buf_2
XFILLER_5_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput1117 output1117/A vssd vssd vccd vccd user2_vcc_powergood sky130_fd_sc_hd__buf_2
XANTENNA_output630_A output630/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output728_A output728/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[122\]_A input285/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[4\] _596_/A la_buf_enable\[4\]/B vssd vssd vccd vccd la_buf\[4\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_31_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[127\]_TE mprj_logic_high_inst/HI[329] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[113\]_A input275/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[35\] input316/X mprj_logic_high_inst/HI[365] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[35\]/B sky130_fd_sc_hd__and2_1
XFILLER_3_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[13\] _605_/A la_buf_enable\[13\]/B vssd vssd vccd vccd la_buf\[13\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_7_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input194_A la_data_out_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input361_A la_iena_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[41\]_TE la_buf\[41\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input459_A la_oenb_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input55_A la_data_out_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input626_A user_irq_ena[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[26\]_TE mprj_logic_high_inst/HI[228] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_50 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[92\]_A_N _355_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[104\]_A input265/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[30\]_A_N _622_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output678_A output678/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_329_ _329_/A vssd vssd vccd vccd _329_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[45\]_A_N _637_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output845_A output845/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[92\] input123/X user_to_mprj_in_gates\[92\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[92\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[64\]_TE la_buf\[64\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[49\]_TE mprj_logic_high_inst/HI[251] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput515 la_oenb_mprj[9] vssd vssd vccd vccd _601_/A sky130_fd_sc_hd__clkbuf_2
Xinput504 la_oenb_mprj[8] vssd vssd vccd vccd _600_/A sky130_fd_sc_hd__buf_2
Xinput526 mprj_adr_o_core[18] vssd vssd vccd vccd _418_/A sky130_fd_sc_hd__buf_2
Xinput537 mprj_adr_o_core[28] vssd vssd vccd vccd _428_/A sky130_fd_sc_hd__buf_2
Xinput559 mprj_dat_i_user[18] vssd vssd vccd vccd input559/X sky130_fd_sc_hd__buf_12
Xuser_to_mprj_oen_buffers\[109\] _372_/Y mprj_logic_high_inst/HI[311] vssd vssd vccd
+ vccd output893/A sky130_fd_sc_hd__einvp_2
XFILLER_25_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput548 mprj_adr_o_core[9] vssd vssd vccd vccd _409_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[93\]_A input380/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[39\] _631_/Y mprj_logic_high_inst/HI[241] vssd vssd vccd
+ vccd output943/A sky130_fd_sc_hd__einvp_8
XFILLER_16_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input207_A la_data_out_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_41 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input576_A mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[13\]_TE mprj_dat_buf\[13\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__402__A _402_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[84\]_A input370/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[62\] user_to_mprj_in_gates\[62\]/Y vssd vssd vccd vccd output841/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_1_1842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output795_A output795/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output962_A output962/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[87\]_TE la_buf\[87\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_wb_dat_gates\[20\] input562/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[20\]/Y
+ sky130_fd_sc_hd__nand2_4
XFILLER_50_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[75\]_A input360/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_54 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[80\] _343_/A la_buf_enable\[80\]/B vssd vssd vccd vccd la_buf\[80\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_27_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput301 la_iena_mprj[21] vssd vssd vccd vccd input301/X sky130_fd_sc_hd__clkbuf_1
Xinput312 la_iena_mprj[31] vssd vssd vccd vccd input312/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input157_A la_data_out_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput334 la_iena_mprj[51] vssd vssd vccd vccd input334/X sky130_fd_sc_hd__clkbuf_1
Xinput323 la_iena_mprj[41] vssd vssd vccd vccd input323/X sky130_fd_sc_hd__clkbuf_1
Xinput345 la_iena_mprj[61] vssd vssd vccd vccd input345/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_74 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input324_A la_iena_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput356 la_iena_mprj[71] vssd vssd vccd vccd input356/X sky130_fd_sc_hd__clkbuf_1
Xinput367 la_iena_mprj[81] vssd vssd vccd vccd input367/X sky130_fd_sc_hd__clkbuf_1
Xinput378 la_iena_mprj[91] vssd vssd vccd vccd input378/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_in_ena_buf\[66\]_A input350/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input18_A la_data_out_core[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput389 la_oenb_mprj[100] vssd vssd vccd vccd _363_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[66\] _530_/Y la_buf\[66\]/TE vssd vssd vccd vccd output717/A sky130_fd_sc_hd__einvp_8
XFILLER_44_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_594_ _594_/A vssd vssd vccd vccd _594_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_38_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[122\] _586_/Y la_buf\[122\]/TE vssd vssd vccd vccd output652/A sky130_fd_sc_hd__einvp_2
XFILLER_32_1195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput808 output808/A vssd vssd vccd vccd la_data_in_mprj[32] sky130_fd_sc_hd__buf_2
Xoutput819 output819/A vssd vssd vccd vccd la_data_in_mprj[42] sky130_fd_sc_hd__buf_2
XFILLER_4_750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[70\]_B user_to_mprj_in_gates\[70\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output710_A output710/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output808_A output808/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[57\]_A input340/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[55\] input82/X user_to_mprj_in_gates\[55\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[55\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[61\]_B user_to_mprj_in_gates\[61\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[48\]_A input330/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input274_A la_iena_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[52\]_B user_to_mprj_in_gates\[52\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input441_A la_oenb_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input539_A mprj_adr_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput120 la_data_out_core[8] vssd vssd vccd vccd input120/X sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput131 la_data_out_core[9] vssd vssd vccd vccd input131/X sky130_fd_sc_hd__buf_2
XFILLER_7_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput142 la_data_out_mprj[109] vssd vssd vccd vccd _573_/A sky130_fd_sc_hd__clkbuf_4
Xinput153 la_data_out_mprj[119] vssd vssd vccd vccd _583_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_ena_buf\[39\]_A input320/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput164 la_data_out_mprj[13] vssd vssd vccd vccd _477_/A sky130_fd_sc_hd__clkbuf_2
Xinput175 la_data_out_mprj[23] vssd vssd vccd vccd _487_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput186 la_data_out_mprj[33] vssd vssd vccd vccd _497_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput197 la_data_out_mprj[43] vssd vssd vccd vccd _507_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_646_ _646_/A vssd vssd vccd vccd _646_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_654 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_577_ _577_/A vssd vssd vccd vccd _577_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[6\]_A _438_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output660_A output660/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[25\] user_to_mprj_in_gates\[25\]/Y vssd vssd vccd vccd output800/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_16_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output758_A output758/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput627 output627/A vssd vssd vccd vccd la_data_in_core[0] sky130_fd_sc_hd__buf_2
XFILLER_12_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[43\]_B user_to_mprj_in_gates\[43\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output925_A output925/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput638 output638/A vssd vssd vccd vccd la_data_in_core[10] sky130_fd_sc_hd__buf_2
Xoutput649 output649/A vssd vssd vccd vccd la_data_in_core[11] sky130_fd_sc_hd__buf_2
XANTENNA_la_buf\[112\]_TE la_buf\[112\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[27\]_TE mprj_adr_buf\[27\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_19 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[34\]_B user_to_mprj_in_gates\[34\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[95\]_A user_to_mprj_in_gates\[95\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output1022_A output1022/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__500__A _500_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[65\] input349/X mprj_logic_high_inst/HI[395] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[65\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_500_ _500_/A vssd vssd vccd vccd _500_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[3\] _595_/Y mprj_logic_high_inst/HI[205] vssd vssd vccd
+ vccd output944/A sky130_fd_sc_hd__einvp_2
X_431_ _431_/A vssd vssd vccd vccd _431_/Y sky130_fd_sc_hd__clkinv_8
Xuser_to_mprj_oen_buffers\[21\] _613_/Y mprj_logic_high_inst/HI[223] vssd vssd vccd
+ vccd output924/A sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[43\] _635_/A la_buf_enable\[43\]/B vssd vssd vccd vccd la_buf\[43\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_1277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_362_ _362_/A vssd vssd vccd vccd _362_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input489_A la_oenb_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input391_A la_oenb_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input85_A la_data_out_core[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[122\]_A _586_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[29\] _493_/Y la_buf\[29\]/TE vssd vssd vccd vccd output676/A sky130_fd_sc_hd__einvp_8
XFILLER_13_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[25\]_B user_to_mprj_in_gates\[25\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[86\]_A user_to_mprj_in_gates\[86\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__410__A _410_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[10\]_A user_to_mprj_in_gates\[10\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_629_ _629_/A vssd vssd vccd vccd _629_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output875_A output875/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[18\] input41/X user_to_mprj_in_gates\[18\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[18\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_buffers\[124\]_A user_to_mprj_in_gates\[124\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[113\]_A _577_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[16\]_B user_to_mprj_in_gates\[16\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[77\]_A user_to_mprj_in_gates\[77\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[28\] user_wb_dat_gates\[28\]/Y vssd vssd vccd vccd output1065/A
+ sky130_fd_sc_hd__inv_6
XFILLER_47_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[50\]_A _514_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[100\]_B user_to_mprj_in_gates\[100\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[82\]_TE mprj_logic_high_inst/HI[284] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[115\]_A user_to_mprj_in_gates\[115\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[104\]_A _568_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[68\]_A user_to_mprj_in_gates\[68\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[41\]_A _505_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput980 output980/A vssd vssd vccd vccd la_oenb_core[72] sky130_fd_sc_hd__buf_2
Xoutput991 output991/A vssd vssd vccd vccd la_oenb_core[82] sky130_fd_sc_hd__buf_2
XFILLER_2_369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[69\] _332_/Y mprj_logic_high_inst/HI[271] vssd vssd vccd
+ vccd output976/A sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[17\] _449_/Y mprj_dat_buf\[17\]/TE vssd vssd vccd vccd output1085/A
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input237_A la_data_out_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input404_A la_oenb_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1074 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_414_ _414_/A vssd vssd vccd vccd _414_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_53_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_345_ _345_/A vssd vssd vccd vccd _345_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[120\] input283/X mprj_logic_high_inst/HI[450] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[120\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_buffers\[106\]_A user_to_mprj_in_gates\[106\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__405__A _405_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[59\]_A user_to_mprj_in_gates\[59\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xoutput1107 output1107/A vssd vssd vccd vccd mprj_dat_o_user[8] sky130_fd_sc_hd__buf_2
XANTENNA_la_buf\[32\]_A _496_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput1118 output1118/A vssd vssd vccd vccd user2_vdd_powergood sky130_fd_sc_hd__buf_2
Xmprj_adr_buf\[12\] _412_/Y mprj_adr_buf\[12\]/TE vssd vssd vccd vccd output1015/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_42_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[50\]_B la_buf_enable\[50\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[126\] user_to_mprj_in_gates\[126\]/Y vssd vssd vccd vccd
+ output784/A sky130_fd_sc_hd__clkinv_4
XFILLER_46_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[92\] user_to_mprj_in_gates\[92\]/Y vssd vssd vccd vccd output874/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_42_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output992_A output992/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[122\]_B mprj_logic_high_inst/HI[452] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[99\]_A _563_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[2\] user_wb_dat_gates\[2\]/Y vssd vssd vccd vccd output1067/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_36_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[23\]_A _487_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[41\]_B la_buf_enable\[41\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[113\]_B mprj_logic_high_inst/HI[443] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_16_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[28\] input308/X mprj_logic_high_inst/HI[358] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[28\]/B sky130_fd_sc_hd__and2_1
XFILLER_3_1394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input187_A la_data_out_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[14\]_A _478_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[32\]_B la_buf_enable\[32\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input354_A la_iena_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input48_A la_data_out_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[1\]_A input299/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input521_A mprj_adr_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input619_A mprj_stb_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[111\] _374_/A la_buf_enable\[111\]/B vssd vssd vccd vccd la_buf\[111\]/TE
+ sky130_fd_sc_hd__and2b_1
Xla_buf\[96\] _560_/Y la_buf\[96\]/TE vssd vssd vccd vccd output750/A sky130_fd_sc_hd__einvp_4
Xuser_to_mprj_in_ena_buf\[1\] input299/X mprj_logic_high_inst/HI[331] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[1\]/B sky130_fd_sc_hd__and2_1
XFILLER_4_1103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[104\]_B mprj_logic_high_inst/HI[434] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_2140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[99\]_B la_buf_enable\[99\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output740_A output740/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output838_A output838/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[23\]_B la_buf_enable\[23\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[85\] input115/X user_to_mprj_in_gates\[85\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[85\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_516 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[92\]_A _355_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[14\]_B la_buf_enable\[14\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput516 mprj_ack_i_user vssd vssd vccd vccd input516/X sky130_fd_sc_hd__buf_12
Xinput505 la_oenb_mprj[90] vssd vssd vccd vccd _353_/A sky130_fd_sc_hd__buf_2
Xinput527 mprj_adr_o_core[19] vssd vssd vccd vccd _419_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_output1102_A output1102/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput549 mprj_cyc_o_core vssd vssd vccd vccd _393_/A sky130_fd_sc_hd__clkbuf_2
Xinput538 mprj_adr_o_core[29] vssd vssd vccd vccd _429_/A sky130_fd_sc_hd__buf_2
XFILLER_29_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[93\]_B mprj_logic_high_inst/HI[423] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input102_A la_data_out_core[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[83\]_A _346_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input471_A la_oenb_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input569_A mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[7\] _471_/Y la_buf\[7\]/TE vssd vssd vccd vccd output732/A sky130_fd_sc_hd__einvp_8
Xla_buf\[11\] _475_/Y la_buf\[11\]/TE vssd vssd vccd vccd output649/A sky130_fd_sc_hd__einvp_8
XFILLER_4_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[4\] _404_/Y mprj_adr_buf\[4\]/TE vssd vssd vccd vccd output1038/A sky130_fd_sc_hd__einvp_4
XFILLER_47_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[84\]_B mprj_logic_high_inst/HI[414] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[55\] user_to_mprj_in_gates\[55\]/Y vssd vssd vccd vccd output833/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output690_A output690/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output788_A output788/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[117\]_TE mprj_logic_high_inst/HI[319] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[74\]_A _337_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[13\] input554/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[13\]/Y
+ sky130_fd_sc_hd__nand2_2
XANTENNA_output955_A output955/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_buffers\[10\] user_wb_dat_gates\[10\]/Y vssd vssd vccd vccd output1046/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_48_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[1\]_A input561/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[75\]_B mprj_logic_high_inst/HI[405] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[111\] input17/X user_to_mprj_in_gates\[111\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[111\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1618 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[31\]_TE la_buf\[31\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[1\]_A input43/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[65\]_A _657_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[16\]_TE mprj_logic_high_inst/HI[218] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[91\]_A_N _354_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1052_A output1052/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__503__A _503_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[95\] input382/X mprj_logic_high_inst/HI[425] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[95\]/B sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[121\] _384_/Y mprj_logic_high_inst/HI[323] vssd vssd vccd
+ vccd output907/A sky130_fd_sc_hd__einvp_4
XFILLER_7_2208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_sel_buf\[2\] _398_/Y mprj_sel_buf\[2\]/TE vssd vssd vccd vccd output1111/A sky130_fd_sc_hd__einvp_8
Xinput302 la_iena_mprj[22] vssd vssd vccd vccd input302/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput335 la_iena_mprj[52] vssd vssd vccd vccd input335/X sky130_fd_sc_hd__clkbuf_1
Xinput324 la_iena_mprj[42] vssd vssd vccd vccd input324/X sky130_fd_sc_hd__clkbuf_1
Xinput313 la_iena_mprj[32] vssd vssd vccd vccd input313/X sky130_fd_sc_hd__clkbuf_1
Xuser_to_mprj_oen_buffers\[51\] _643_/Y mprj_logic_high_inst/HI[253] vssd vssd vccd
+ vccd output957/A sky130_fd_sc_hd__einvp_2
Xla_buf_enable\[73\] _336_/A la_buf_enable\[73\]/B vssd vssd vccd vccd la_buf\[73\]/TE
+ sky130_fd_sc_hd__and2b_1
Xinput346 la_iena_mprj[62] vssd vssd vccd vccd input346/X sky130_fd_sc_hd__clkbuf_1
Xinput357 la_iena_mprj[72] vssd vssd vccd vccd input357/X sky130_fd_sc_hd__clkbuf_1
Xinput368 la_iena_mprj[82] vssd vssd vccd vccd input368/X sky130_fd_sc_hd__clkbuf_1
Xinput379 la_iena_mprj[92] vssd vssd vccd vccd input379/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_in_ena_buf\[66\]_B mprj_logic_high_inst/HI[396] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input317_A la_iena_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[44\]_A_N _636_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_593_ _593_/A vssd vssd vccd vccd _593_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[59\] _523_/Y la_buf\[59\]/TE vssd vssd vccd vccd output709/A sky130_fd_sc_hd__einvp_8
XFILLER_44_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[59\]_A_N _651_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[56\]_A _648_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput809 output809/A vssd vssd vccd vccd la_data_in_mprj[33] sky130_fd_sc_hd__buf_2
XFILLER_49_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[115\] _579_/Y la_buf\[115\]/TE vssd vssd vccd vccd output644/A sky130_fd_sc_hd__einvp_4
XANTENNA__413__A _413_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output703_A output703/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[57\]_B mprj_logic_high_inst/HI[387] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[54\]_TE la_buf\[54\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[39\]_TE mprj_logic_high_inst/HI[241] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[48\] input74/X user_to_mprj_in_gates\[48\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[48\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_50_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[47\]_A _639_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[48\]_B mprj_logic_high_inst/HI[378] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[10\] input271/X mprj_logic_high_inst/HI[340] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[10\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[38\]_A _630_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_76 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[99\] _362_/Y mprj_logic_high_inst/HI[301] vssd vssd vccd
+ vccd output1009/A sky130_fd_sc_hd__einvp_8
XANTENNA_input267_A la_iena_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj2_vdd_pwrgood mprj2_vdd_pwrgood/A vssd vssd vccd vccd output1118/A sky130_fd_sc_hd__buf_6
XFILLER_1_732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput110 la_data_out_core[80] vssd vssd vccd vccd input110/X sky130_fd_sc_hd__buf_4
XFILLER_46_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[77\]_TE la_buf\[77\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input434_A la_oenb_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input30_A la_data_out_core[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput121 la_data_out_core[90] vssd vssd vccd vccd input121/X sky130_fd_sc_hd__buf_4
Xinput143 la_data_out_mprj[10] vssd vssd vccd vccd _474_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput132 la_data_out_mprj[0] vssd vssd vccd vccd _464_/A sky130_fd_sc_hd__clkbuf_2
Xinput154 la_data_out_mprj[11] vssd vssd vccd vccd _475_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput165 la_data_out_mprj[14] vssd vssd vccd vccd _478_/A sky130_fd_sc_hd__clkbuf_2
Xinput176 la_data_out_mprj[24] vssd vssd vccd vccd _488_/A sky130_fd_sc_hd__clkbuf_2
Xinput187 la_data_out_mprj[34] vssd vssd vccd vccd _498_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input601_A mprj_dat_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[39\]_B mprj_logic_high_inst/HI[369] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput198 la_data_out_mprj[44] vssd vssd vccd vccd _508_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_645_ _645_/A vssd vssd vccd vccd _645_/Y sky130_fd_sc_hd__clkinv_2
X_576_ _576_/A vssd vssd vccd vccd _576_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__408__A _408_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[29\]_A _621_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[18\] user_to_mprj_in_gates\[18\]/Y vssd vssd vccd vccd output792/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output653_A output653/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput639 output639/A vssd vssd vccd vccd la_data_in_core[110] sky130_fd_sc_hd__buf_2
Xoutput628 output628/A vssd vssd vccd vccd la_data_in_core[100] sky130_fd_sc_hd__buf_2
XANTENNA_output918_A output918/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output820_A output820/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[25\]_A _425_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1674 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[26\]_TE mprj_dat_buf\[26\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[5\]_TE mprj_logic_high_inst/HI[207] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_23_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_488 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[2\]_A _594_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[16\]_A _416_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1015_A output1015/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[58\] input341/X mprj_logic_high_inst/HI[388] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[58\]/B sky130_fd_sc_hd__and2_1
XTAP_680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_430_ _430_/A vssd vssd vccd vccd _430_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_26_452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_54 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[14\] _606_/Y mprj_logic_high_inst/HI[216] vssd vssd vccd
+ vccd output916/A sky130_fd_sc_hd__einvp_4
X_361_ _361_/A vssd vssd vccd vccd _361_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[36\] _628_/A la_buf_enable\[36\]/B vssd vssd vccd vccd la_buf\[36\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_1879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input384_A la_iena_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input78_A la_data_out_core[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input551_A mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_sel_buf\[0\]_TE mprj_sel_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_628_ _628_/A vssd vssd vccd vccd _628_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1710 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_559_ _559_/A vssd vssd vccd vccd _559_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output770_A output770/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output868_A output868/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__601__A _601_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput981 output981/A vssd vssd vccd vccd la_oenb_core[73] sky130_fd_sc_hd__buf_2
Xoutput970 output970/A vssd vssd vccd vccd la_oenb_core[63] sky130_fd_sc_hd__buf_2
XFILLER_47_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__511__A _511_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput992 output992/A vssd vssd vccd vccd la_oenb_core[83] sky130_fd_sc_hd__buf_2
XFILLER_8_1443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input132_A la_data_out_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_413_ _413_/A vssd vssd vccd vccd _413_/Y sky130_fd_sc_hd__inv_6
XFILLER_42_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input599_A mprj_dat_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[102\]_TE la_buf\[102\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_344_ _344_/A vssd vssd vccd vccd _344_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[41\] _505_/Y la_buf\[41\]/TE vssd vssd vccd vccd output690/A sky130_fd_sc_hd__einvp_8
XFILLER_30_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[113\] input275/X mprj_logic_high_inst/HI[443] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[113\]/B sky130_fd_sc_hd__and2_1
XFILLER_31_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[17\]_TE mprj_adr_buf\[17\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput1108 output1108/A vssd vssd vccd vccd mprj_dat_o_user[9] sky130_fd_sc_hd__buf_2
Xoutput1119 output1119/A vssd vssd vccd vccd user_clock sky130_fd_sc_hd__buf_2
XANTENNA_mprj_adr_buf\[1\]_TE mprj_adr_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__421__A _421_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[119\] user_to_mprj_in_gates\[119\]/Y vssd vssd vccd vccd
+ output776/A sky130_fd_sc_hd__clkinv_4
XFILLER_42_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[29\]_A _461_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[85\] user_to_mprj_in_gates\[85\]/Y vssd vssd vccd vccd output866/A
+ sky130_fd_sc_hd__inv_2
XFILLER_49_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output985_A output985/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[30\] input55/X user_to_mprj_in_gates\[30\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[30\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[1\]_A _401_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__331__A _331_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[5\]_TE mprj_dat_buf\[5\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[27\]_A user_wb_dat_gates\[27\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_5_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[125\]_TE la_buf\[125\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_ack_gate_A input516/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output1082_A output1082/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__506__A _506_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[81\] _344_/Y mprj_logic_high_inst/HI[283] vssd vssd vccd
+ vccd output990/A sky130_fd_sc_hd__einvp_4
XFILLER_30_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input347_A la_iena_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[1\]_B mprj_logic_high_inst/HI[331] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[18\]_A user_wb_dat_gates\[18\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_48_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input514_A la_oenb_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[89\] _553_/Y la_buf\[89\]/TE vssd vssd vccd vccd output742/A sky130_fd_sc_hd__einvp_8
XFILLER_4_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[104\] _367_/A la_buf_enable\[104\]/B vssd vssd vccd vccd la_buf\[104\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_2141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[72\]_TE mprj_logic_high_inst/HI[274] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__416__A _416_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output733_A output733/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output900_A output900/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[78\] input107/X user_to_mprj_in_gates\[78\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[78\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[122\]_B la_buf_enable\[122\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[91\]_A input122/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj2_pwrgood_A mprj2_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput506 la_oenb_mprj[91] vssd vssd vccd vccd _354_/A sky130_fd_sc_hd__clkbuf_4
Xinput517 mprj_adr_o_core[0] vssd vssd vccd vccd _400_/A sky130_fd_sc_hd__buf_12
Xinput528 mprj_adr_o_core[1] vssd vssd vccd vccd _401_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput539 mprj_adr_o_core[2] vssd vssd vccd vccd _402_/A sky130_fd_sc_hd__buf_12
XFILLER_28_300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[113\]_B la_buf_enable\[113\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[40\] input322/X mprj_logic_high_inst/HI[370] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[40\]/B sky130_fd_sc_hd__and2_1
XFILLER_44_826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[95\]_TE mprj_logic_high_inst/HI[297] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input297_A la_iena_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[4\]_A user_wb_dat_gates\[4\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[82\]_A input112/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input60_A la_data_out_core[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input464_A la_oenb_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[7\]_A _471_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[104\]_B la_buf_enable\[104\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[48\] user_to_mprj_in_gates\[48\]/Y vssd vssd vccd vccd output825/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_15_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output683_A output683/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output850_A output850/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output948_A output948/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[73\]_A input102/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[1\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[104\] input9/X user_to_mprj_in_gates\[104\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[104\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[1\]_B user_to_mprj_in_gates\[1\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[64\]_A input92/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output1045_A output1045/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[88\] input374/X mprj_logic_high_inst/HI[418] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[88\]/B sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[114\] _377_/Y mprj_logic_high_inst/HI[316] vssd vssd vccd
+ vccd output899/A sky130_fd_sc_hd__einvp_4
Xinput303 la_iena_mprj[23] vssd vssd vccd vccd input303/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput336 la_iena_mprj[53] vssd vssd vccd vccd input336/X sky130_fd_sc_hd__clkbuf_1
Xinput325 la_iena_mprj[43] vssd vssd vccd vccd input325/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput314 la_iena_mprj[33] vssd vssd vccd vccd input314/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput347 la_iena_mprj[63] vssd vssd vccd vccd input347/X sky130_fd_sc_hd__clkbuf_1
Xinput358 la_iena_mprj[73] vssd vssd vccd vccd input358/X sky130_fd_sc_hd__clkbuf_1
Xinput369 la_iena_mprj[83] vssd vssd vccd vccd input369/X sky130_fd_sc_hd__clkbuf_1
Xuser_to_mprj_oen_buffers\[44\] _636_/Y mprj_logic_high_inst/HI[246] vssd vssd vccd
+ vccd output949/A sky130_fd_sc_hd__einvp_2
Xla_buf_enable\[66\] _329_/A la_buf_enable\[66\]/B vssd vssd vccd vccd la_buf\[66\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_29_642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_irq_buffers\[2\] user_irq_gates\[2\]/Y vssd vssd vccd vccd output1123/A sky130_fd_sc_hd__clkinv_4
XFILLER_44_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_592_ _592_/A vssd vssd vccd vccd _592_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input212_A la_data_out_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input581_A mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[55\]_A input82/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_69 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[108\] _572_/Y la_buf\[108\]/TE vssd vssd vccd vccd output636/A sky130_fd_sc_hd__einvp_4
XTAP_317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[101\] user_to_mprj_in_gates\[101\]/Y vssd vssd vccd vccd
+ output757/A sky130_fd_sc_hd__clkinv_4
XFILLER_48_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1878 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output898_A output898/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[5\]_A user_to_mprj_in_gates\[5\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1674 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__604__A _604_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[46\]_A input72/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[0\] _432_/Y mprj_dat_buf\[0\]/TE vssd vssd vccd vccd output1077/A sky130_fd_sc_hd__einvp_8
XTAP_862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_464 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__514__A _514_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[121\]_A input28/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[37\]_A input62/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_88 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input162_A la_data_out_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput111 la_data_out_core[81] vssd vssd vccd vccd input111/X sky130_fd_sc_hd__buf_4
Xinput100 la_data_out_core[71] vssd vssd vccd vccd input100/X sky130_fd_sc_hd__buf_4
XFILLER_42_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput122 la_data_out_core[91] vssd vssd vccd vccd input122/X sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[107\]_TE mprj_logic_high_inst/HI[309] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input427_A la_oenb_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput133 la_data_out_mprj[100] vssd vssd vccd vccd _564_/A sky130_fd_sc_hd__buf_2
Xinput144 la_data_out_mprj[110] vssd vssd vccd vccd _574_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input23_A la_data_out_core[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput166 la_data_out_mprj[15] vssd vssd vccd vccd _479_/A sky130_fd_sc_hd__clkbuf_2
Xinput177 la_data_out_mprj[25] vssd vssd vccd vccd _489_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput155 la_data_out_mprj[120] vssd vssd vccd vccd _584_/A sky130_fd_sc_hd__clkbuf_2
X_644_ _644_/A vssd vssd vccd vccd _644_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput199 la_data_out_mprj[45] vssd vssd vccd vccd _509_/A sky130_fd_sc_hd__clkbuf_2
Xinput188 la_data_out_mprj[35] vssd vssd vccd vccd _499_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xla_buf\[71\] _535_/Y la_buf\[71\]/TE vssd vssd vccd vccd output723/A sky130_fd_sc_hd__einvp_4
XFILLER_45_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_575_ _575_/A vssd vssd vccd vccd _575_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__424__A _424_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[28\]_A input52/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[112\]_A input18/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput629 output629/A vssd vssd vccd vccd la_data_in_core[101] sky130_fd_sc_hd__buf_2
XANTENNA_output646_A output646/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[21\]_TE la_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output813_A output813/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[90\]_A_N _353_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[60\] input88/X user_to_mprj_in_gates\[60\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[60\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[19\]_A input42/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__334__A _334_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[103\]_A input8/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[43\]_A_N _635_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[58\]_A_N _650_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output1008_A output1008/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__509__A _509_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_360_ _360_/A vssd vssd vccd vccd _360_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[29\] _621_/A la_buf_enable\[29\]/B vssd vssd vccd vccd la_buf\[29\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_42_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[44\]_TE la_buf\[44\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input377_A la_iena_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[29\]_TE mprj_logic_high_inst/HI[231] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input544_A mprj_adr_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_627_ _627_/A vssd vssd vccd vccd _627_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__419__A _419_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_558_ _558_/A vssd vssd vccd vccd _558_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_489_ _489_/A vssd vssd vccd vccd _489_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[30\] user_to_mprj_in_gates\[30\]/Y vssd vssd vccd vccd output806/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_51_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output763_A output763/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output930_A output930/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[1\]_B la_buf_enable\[1\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[125\]_A input288/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__329__A _329_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[67\]_TE la_buf\[67\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput982 output982/A vssd vssd vccd vccd la_oenb_core[74] sky130_fd_sc_hd__buf_2
Xoutput971 output971/A vssd vssd vccd vccd la_oenb_core[64] sky130_fd_sc_hd__buf_2
Xoutput960 output960/A vssd vssd vccd vccd la_oenb_core[54] sky130_fd_sc_hd__buf_2
XFILLER_28_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[70\] input355/X mprj_logic_high_inst/HI[400] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[70\]/B sky130_fd_sc_hd__and2_1
Xoutput993 output993/A vssd vssd vccd vccd la_oenb_core[84] sky130_fd_sc_hd__buf_2
XFILLER_47_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[116\]_A input278/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input125_A la_data_out_core[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_412_ _412_/A vssd vssd vccd vccd _412_/Y sky130_fd_sc_hd__inv_8
XFILLER_53_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_343_ _343_/A vssd vssd vccd vccd _343_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input494_A la_oenb_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input90_A la_data_out_core[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[34\] _498_/Y la_buf\[34\]/TE vssd vssd vccd vccd output682/A sky130_fd_sc_hd__einvp_8
XFILLER_31_1218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[106\] input267/X mprj_logic_high_inst/HI[436] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[106\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[6\] input578/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[6\]/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_13_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_9 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[16\]_TE mprj_dat_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput1109 output1109/A vssd vssd vccd vccd mprj_sel_o_user[0] sky130_fd_sc_hd__buf_2
XFILLER_48_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[107\]_A input268/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[78\] user_to_mprj_in_gates\[78\]/Y vssd vssd vccd vccd output858/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_40_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output978_A output978/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output880_A output880/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[23\] input47/X user_to_mprj_in_gates\[23\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[23\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__612__A _612_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_ack_gate_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output1075_A output1075/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__522__A _522_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[74\] _337_/Y mprj_logic_high_inst/HI[276] vssd vssd vccd
+ vccd output982/A sky130_fd_sc_hd__einvp_4
Xla_buf_enable\[96\] _359_/A la_buf_enable\[96\]/B vssd vssd vccd vccd la_buf\[96\]/TE
+ sky130_fd_sc_hd__and2b_1
Xoutput790 output790/A vssd vssd vccd vccd la_data_in_mprj[16] sky130_fd_sc_hd__buf_2
XFILLER_43_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[22\] _454_/Y mprj_dat_buf\[22\]/TE vssd vssd vccd vccd output1091/A
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input242_A la_data_out_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[96\]_A input383/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input507_A la_oenb_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[20\]_A input300/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__432__A _432_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output726_A output726/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[87\]_A input373/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__607__A _607_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[11\]_A input282/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[2\] _594_/A la_buf_enable\[2\]/B vssd vssd vccd vccd la_buf\[2\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_20_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[91\]_B user_to_mprj_in_gates\[91\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__342__A _342_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput507 la_oenb_mprj[92] vssd vssd vccd vccd _355_/A sky130_fd_sc_hd__buf_2
Xinput518 mprj_adr_o_core[10] vssd vssd vccd vccd _410_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_in_ena_buf\[78\]_A input363/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2076 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput529 mprj_adr_o_core[20] vssd vssd vccd vccd _420_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[33\] input314/X mprj_logic_high_inst/HI[363] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[33\]/B sky130_fd_sc_hd__and2_1
XFILLER_43_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__517__A _517_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[11\] _603_/A la_buf_enable\[11\]/B vssd vssd vccd vccd la_buf\[11\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_8_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input192_A la_data_out_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[82\]_B user_to_mprj_in_gates\[82\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input457_A la_oenb_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input53_A la_data_out_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input624_A user_irq_ena[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[69\]_A input353/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__427__A _427_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output676_A output676/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[73\]_B user_to_mprj_in_gates\[73\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output843_A output843/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[115\]_TE la_buf\[115\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[90\] input121/X user_to_mprj_in_gates\[90\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[90\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__337__A _337_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[64\]_B user_to_mprj_in_gates\[64\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1038_A output1038/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[62\]_TE mprj_logic_high_inst/HI[264] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput326 la_iena_mprj[44] vssd vssd vccd vccd input326/X sky130_fd_sc_hd__clkbuf_1
Xinput304 la_iena_mprj[24] vssd vssd vccd vccd input304/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput315 la_iena_mprj[34] vssd vssd vccd vccd input315/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[107\] _370_/Y mprj_logic_high_inst/HI[309] vssd vssd vccd
+ vccd output891/A sky130_fd_sc_hd__einvp_4
XFILLER_29_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput337 la_iena_mprj[54] vssd vssd vccd vccd input337/X sky130_fd_sc_hd__clkbuf_1
Xinput348 la_iena_mprj[64] vssd vssd vccd vccd input348/X sky130_fd_sc_hd__clkbuf_1
Xinput359 la_iena_mprj[74] vssd vssd vccd vccd input359/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[59\] _651_/A la_buf_enable\[59\]/B vssd vssd vccd vccd la_buf\[59\]/TE
+ sky130_fd_sc_hd__and2b_1
X_591_ _591_/A vssd vssd vccd vccd _591_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[37\] _629_/Y mprj_logic_high_inst/HI[239] vssd vssd vccd
+ vccd output941/A sky130_fd_sc_hd__einvp_4
XFILLER_44_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input205_A la_data_out_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input574_A mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[55\]_B user_to_mprj_in_gates\[55\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[40\]_A user_to_mprj_in_gates\[40\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[60\] user_to_mprj_in_gates\[60\]/Y vssd vssd vccd vccd output839/A
+ sky130_fd_sc_hd__inv_2
XFILLER_34_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[9\]_A _441_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output793_A output793/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output960_A output960/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[46\]_B user_to_mprj_in_gates\[46\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[80\]_A _544_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[85\]_TE mprj_logic_high_inst/HI[287] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__620__A _620_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[31\]_A user_to_mprj_in_gates\[31\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[98\]_A user_to_mprj_in_gates\[98\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[37\]_B user_to_mprj_in_gates\[37\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[71\]_A _535_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[121\]_B user_to_mprj_in_gates\[121\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__530__A _530_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput101 la_data_out_core[72] vssd vssd vccd vccd input101/X sky130_fd_sc_hd__buf_4
XFILLER_46_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input155_A la_data_out_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput123 la_data_out_core[92] vssd vssd vccd vccd input123/X sky130_fd_sc_hd__buf_4
Xinput112 la_data_out_core[82] vssd vssd vccd vccd input112/X sky130_fd_sc_hd__buf_4
XFILLER_49_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput134 la_data_out_mprj[101] vssd vssd vccd vccd _565_/A sky130_fd_sc_hd__buf_2
Xinput145 la_data_out_mprj[111] vssd vssd vccd vccd _575_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input322_A la_iena_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput167 la_data_out_mprj[16] vssd vssd vccd vccd _480_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput178 la_data_out_mprj[26] vssd vssd vccd vccd _490_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput156 la_data_out_mprj[121] vssd vssd vccd vccd _585_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_input16_A la_data_out_core[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_643_ _643_/A vssd vssd vccd vccd _643_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[22\]_A user_to_mprj_in_gates\[22\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_17_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput189 la_data_out_mprj[36] vssd vssd vccd vccd _500_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_44_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2020 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[64\] _528_/Y la_buf\[64\]/TE vssd vssd vccd vccd output715/A sky130_fd_sc_hd__einvp_8
XFILLER_45_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[30\]_A input573/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_574_ _574_/A vssd vssd vccd vccd _574_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[125\]_A _589_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[28\]_B user_to_mprj_in_gates\[28\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[89\]_A user_to_mprj_in_gates\[89\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[62\]_A _526_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[112\]_B user_to_mprj_in_gates\[112\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf\[120\] _584_/Y la_buf\[120\]/TE vssd vssd vccd vccd output650/A sky130_fd_sc_hd__einvp_2
Xmprj_adr_buf\[28\] _428_/Y mprj_adr_buf\[28\]/TE vssd vssd vccd vccd output1032/A
+ sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[80\]_B la_buf_enable\[80\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output639_A output639/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__440__A _440_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output806_A output806/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[53\] input80/X user_to_mprj_in_gates\[53\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[53\]/Y sky130_fd_sc_hd__nand2_2
XANTENNA_user_to_mprj_in_buffers\[13\]_A user_to_mprj_in_gates\[13\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[21\]_A input563/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[127\]_A user_to_mprj_in_gates\[127\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[116\]_A _580_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__615__A _615_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[19\]_B user_to_mprj_in_gates\[19\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[53\]_A _517_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_B user_to_mprj_in_gates\[103\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1046 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[71\]_B la_buf_enable\[71\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__350__A _350_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input8_A la_data_out_core[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[12\]_A input553/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[118\]_A user_to_mprj_in_gates\[118\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[107\]_A _571_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__525__A _525_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[44\]_A _508_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[62\]_B la_buf_enable\[62\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input272_A la_iena_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input537_A mprj_adr_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[127\] _390_/A la_buf_enable\[127\]/B vssd vssd vccd vccd la_buf\[127\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_24_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_626_ _626_/A vssd vssd vccd vccd _626_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_557_ _557_/A vssd vssd vccd vccd _557_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_2337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[109\]_A user_to_mprj_in_gates\[109\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_488_ _488_/A vssd vssd vccd vccd _488_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__435__A _435_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[35\]_A _499_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[23\] user_to_mprj_in_gates\[23\]/Y vssd vssd vccd vccd output798/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output756_A output756/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[53\]_B la_buf_enable\[53\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output923_A output923/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[120\]_A _383_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[125\]_B mprj_logic_high_inst/HI[455] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__345__A _345_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[26\]_A _490_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[44\]_B la_buf_enable\[44\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput972 output972/A vssd vssd vccd vccd la_oenb_core[65] sky130_fd_sc_hd__buf_2
Xoutput961 output961/A vssd vssd vccd vccd la_oenb_core[55] sky130_fd_sc_hd__buf_2
Xoutput950 output950/A vssd vssd vccd vccd la_oenb_core[45] sky130_fd_sc_hd__buf_2
XFILLER_47_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput983 output983/A vssd vssd vccd vccd la_oenb_core[75] sky130_fd_sc_hd__buf_2
Xoutput994 output994/A vssd vssd vccd vccd la_oenb_core[85] sky130_fd_sc_hd__buf_2
XANTENNA_output1020_A output1020/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1118_A output1118/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[111\]_A _374_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[63\] input347/X mprj_logic_high_inst/HI[393] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[63\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[116\]_B mprj_logic_high_inst/HI[446] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input118_A la_data_out_core[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[1\] _593_/Y mprj_logic_high_inst/HI[203] vssd vssd vccd
+ vccd output922/A sky130_fd_sc_hd__einvp_4
Xla_buf_enable\[41\] _633_/A la_buf_enable\[41\]/B vssd vssd vccd vccd la_buf\[41\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_26_273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_411_ _411_/A vssd vssd vccd vccd _411_/Y sky130_fd_sc_hd__inv_6
XFILLER_42_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[11\]_TE la_buf\[11\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_342_ _342_/A vssd vssd vccd vccd _342_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_2089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input83_A la_data_out_core[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input487_A la_oenb_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[27\] _491_/Y la_buf\[27\]/TE vssd vssd vccd vccd output674/A sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[17\]_A _481_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[35\]_B la_buf_enable\[35\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[4\]_A input332/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[102\]_A _365_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[107\]_B mprj_logic_high_inst/HI[437] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[42\]_A_N _634_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_609_ _609_/A vssd vssd vccd vccd _609_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_53_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output873_A output873/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[29\] input571/X repeater1125/X vssd vssd vccd vccd user_wb_dat_gates\[29\]/Y
+ sky130_fd_sc_hd__nand2_8
XFILLER_32_287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[16\] input39/X user_to_mprj_in_gates\[16\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[16\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA_la_buf_enable\[57\]_A_N _649_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[26\] user_wb_dat_gates\[26\]/Y vssd vssd vccd vccd output1063/A
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_la_buf_enable\[26\]_B la_buf_enable\[26\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[127\] input34/X user_to_mprj_in_gates\[127\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[127\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[34\]_TE la_buf\[34\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[19\]_TE mprj_logic_high_inst/HI[221] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[95\]_A _358_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_298 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output1068_A output1068/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[17\]_B la_buf_enable\[17\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput780 output780/A vssd vssd vccd vccd la_data_in_mprj[122] sky130_fd_sc_hd__buf_2
XFILLER_47_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[67\] _330_/Y mprj_logic_high_inst/HI[269] vssd vssd vccd
+ vccd output974/A sky130_fd_sc_hd__einvp_2
Xoutput791 output791/A vssd vssd vccd vccd la_data_in_mprj[17] sky130_fd_sc_hd__buf_2
XFILLER_8_1220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[96\]_B mprj_logic_high_inst/HI[426] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[89\] _352_/A la_buf_enable\[89\]/B vssd vssd vccd vccd la_buf\[89\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_48_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[15\] _447_/Y mprj_dat_buf\[15\]/TE vssd vssd vccd vccd output1083/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_19_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input235_A la_data_out_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_39 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input402_A la_oenb_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[86\]_A _349_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[2\]_TE la_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[20\]_B mprj_logic_high_inst/HI[350] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_7 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[10\] _410_/Y mprj_adr_buf\[10\]/TE vssd vssd vccd vccd output1013/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_26_1800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[124\] user_to_mprj_in_gates\[124\]/Y vssd vssd vccd vccd
+ output782/A sky130_fd_sc_hd__clkinv_4
XANTENNA_output719_A output719/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[10\]_A _602_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[87\]_B mprj_logic_high_inst/HI[417] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[57\]_TE la_buf\[57\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[90\] user_to_mprj_in_gates\[90\]/Y vssd vssd vccd vccd output872/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_42_1178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output990_A output990/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[0\] user_wb_dat_gates\[0\]/Y vssd vssd vccd vccd output1045/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_18_582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[77\]_A _340_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[11\]_B mprj_logic_high_inst/HI[341] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__623__A _623_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[4\]_A input576/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput508 la_oenb_mprj[93] vssd vssd vccd vccd _356_/A sky130_fd_sc_hd__buf_2
Xinput519 mprj_adr_o_core[11] vssd vssd vccd vccd _411_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[78\]_B mprj_logic_high_inst/HI[408] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2066 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[4\]_A input76/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[26\] input306/X mprj_logic_high_inst/HI[356] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[26\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[68\]_A _331_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__533__A _533_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input185_A la_data_out_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input352_A la_iena_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input46_A la_data_out_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[69\]_B mprj_logic_high_inst/HI[399] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[94\] _558_/Y la_buf\[94\]/TE vssd vssd vccd vccd output748/A sky130_fd_sc_hd__einvp_4
XFILLER_8_1061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input617_A mprj_sel_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[59\]_A _651_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output669_A output669/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__443__A _443_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output836_A output836/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[83\] input113/X user_to_mprj_in_gates\[83\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[83\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[29\]_TE mprj_dat_buf\[29\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_71 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__618__A _618_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[8\]_TE mprj_logic_high_inst/HI[210] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__353__A _353_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput327 la_iena_mprj[45] vssd vssd vccd vccd input327/X sky130_fd_sc_hd__clkbuf_1
Xinput305 la_iena_mprj[25] vssd vssd vccd vccd input305/X sky130_fd_sc_hd__clkbuf_1
Xinput316 la_iena_mprj[35] vssd vssd vccd vccd input316/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_output1100_A output1100/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput338 la_iena_mprj[55] vssd vssd vccd vccd input338/X sky130_fd_sc_hd__clkbuf_1
Xinput349 la_iena_mprj[65] vssd vssd vccd vccd input349/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_590_ _590_/A vssd vssd vccd vccd _590_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__528__A _528_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input100_A la_data_out_core[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_820 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input567_A mprj_dat_i_user[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[5\] _469_/Y la_buf\[5\]/TE vssd vssd vccd vccd output710/A sky130_fd_sc_hd__einvp_8
XFILLER_6_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_pwrgood_A mprj_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[3\]_TE mprj_sel_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[2\] _402_/Y mprj_adr_buf\[2\]/TE vssd vssd vccd vccd output1034/A sky130_fd_sc_hd__einvp_4
XFILLER_43_1273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__438__A _438_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[53\] user_to_mprj_in_gates\[53\]/Y vssd vssd vccd vccd output831/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_37_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output786_A output786/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_dat_buf\[10\]_A _442_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_gates\[11\] input552/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[11\]/Y
+ sky130_fd_sc_hd__nand2_2
XANTENNA_output953_A output953/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[28\]_A _428_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__348__A _348_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[5\]_A _597_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1050_A output1050/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[93\] input380/X mprj_logic_high_inst/HI[423] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[93\]/B sky130_fd_sc_hd__and2_1
XANTENNA_mprj_adr_buf\[19\]_A _419_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput102 la_data_out_core[73] vssd vssd vccd vccd input102/X sky130_fd_sc_hd__buf_4
XFILLER_44_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_sel_buf\[0\] _396_/Y mprj_sel_buf\[0\]/TE vssd vssd vccd vccd output1109/A sky130_fd_sc_hd__einvp_8
Xinput124 la_data_out_core[93] vssd vssd vccd vccd input124/X sky130_fd_sc_hd__buf_4
Xinput113 la_data_out_core[83] vssd vssd vccd vccd input113/X sky130_fd_sc_hd__buf_4
Xoutput1090 output1090/A vssd vssd vccd vccd mprj_dat_o_user[21] sky130_fd_sc_hd__buf_2
XFILLER_1_779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput135 la_data_out_mprj[102] vssd vssd vccd vccd _566_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input148_A la_data_out_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[71\] _334_/A la_buf_enable\[71\]/B vssd vssd vccd vccd la_buf\[71\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_40_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput168 la_data_out_mprj[17] vssd vssd vccd vccd _481_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput146 la_data_out_mprj[112] vssd vssd vccd vccd _576_/A sky130_fd_sc_hd__clkbuf_4
Xinput157 la_data_out_mprj[122] vssd vssd vccd vccd _586_/A sky130_fd_sc_hd__clkbuf_2
X_642_ _642_/A vssd vssd vccd vccd _642_/Y sky130_fd_sc_hd__clkinv_2
Xinput179 la_data_out_mprj[27] vssd vssd vccd vccd _491_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input315_A la_iena_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[30\]_B repeater1125/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_573_ _573_/A vssd vssd vccd vccd _573_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[57\] _521_/Y la_buf\[57\]/TE vssd vssd vccd vccd output707/A sky130_fd_sc_hd__einvp_8
XFILLER_44_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[105\]_TE la_buf\[105\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_buffers\[2\]_A user_irq_gates\[2\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[113\] _577_/Y la_buf\[113\]/TE vssd vssd vccd vccd output642/A sky130_fd_sc_hd__einvp_4
XANTENNA_mprj_adr_buf\[4\]_TE mprj_adr_buf\[4\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output701_A output701/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[21\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[46\] input72/X user_to_mprj_in_gates\[46\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[46\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[52\]_TE mprj_logic_high_inst/HI[254] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__631__A _631_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[8\]_TE mprj_dat_buf\[8\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[8\] input120/X user_to_mprj_in_gates\[8\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[8\]/Y sky130_fd_sc_hd__nand2_2
XTAP_650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[12\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output1098_A output1098/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[97\] _360_/Y mprj_logic_high_inst/HI[299] vssd vssd vccd
+ vccd output1007/A sky130_fd_sc_hd__einvp_2
XFILLER_13_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__541__A _541_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input265_A la_iena_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input432_A la_oenb_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[90\]_TE la_buf\[90\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_625_ _625_/A vssd vssd vccd vccd _625_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_oen_buffers\[75\]_TE mprj_logic_high_inst/HI[277] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_556_ _556_/A vssd vssd vccd vccd _556_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_487_ _487_/A vssd vssd vccd vccd _487_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_51_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2040 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[16\] user_to_mprj_in_gates\[16\]/Y vssd vssd vccd vccd output790/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output651_A output651/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output749_A output749/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__451__A _451_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output916_A output916/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__626__A _626_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[4\]_A _404_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__361__A _361_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput973 output973/A vssd vssd vccd vccd la_oenb_core[66] sky130_fd_sc_hd__buf_2
Xoutput962 output962/A vssd vssd vccd vccd la_oenb_core[56] sky130_fd_sc_hd__buf_2
Xoutput951 output951/A vssd vssd vccd vccd la_oenb_core[46] sky130_fd_sc_hd__buf_2
Xoutput940 output940/A vssd vssd vccd vccd la_oenb_core[36] sky130_fd_sc_hd__buf_2
Xoutput995 output995/A vssd vssd vccd vccd la_oenb_core[86] sky130_fd_sc_hd__buf_2
Xoutput984 output984/A vssd vssd vccd vccd la_oenb_core[76] sky130_fd_sc_hd__buf_2
XFILLER_47_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output1013_A output1013/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[56\] input339/X mprj_logic_high_inst/HI[386] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[56\]/B sky130_fd_sc_hd__and2_1
XTAP_491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[98\]_TE mprj_logic_high_inst/HI[300] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_410_ _410_/A vssd vssd vccd vccd _410_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_14_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_341_ _341_/A vssd vssd vccd vccd _341_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__536__A _536_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[12\] _604_/Y mprj_logic_high_inst/HI[214] vssd vssd vccd
+ vccd output914/A sky130_fd_sc_hd__einvp_4
Xla_buf_enable\[34\] _626_/A la_buf_enable\[34\]/B vssd vssd vccd vccd la_buf\[34\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[8\] user_to_mprj_in_gates\[8\]/Y vssd vssd vccd vccd output871/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_35_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input382_A la_iena_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input76_A la_data_out_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[4\]_B mprj_logic_high_inst/HI[334] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_830 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_stb_buf _394_/Y mprj_stb_buf/TE vssd vssd vccd vccd output1113/A sky130_fd_sc_hd__einvp_8
XFILLER_2_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_712 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_608_ _608_/A vssd vssd vccd vccd _608_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_1669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output699_A output699/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__446__A _446_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_539_ _539_/A vssd vssd vccd vccd _539_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1598 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output866_A output866/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_buffers\[19\] user_wb_dat_gates\[19\]/Y vssd vssd vccd vccd output1055/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_25_2215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[125\]_B la_buf_enable\[125\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__356__A _356_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_542 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[94\]_A input125/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput770 output770/A vssd vssd vccd vccd la_data_in_mprj[113] sky130_fd_sc_hd__buf_2
Xoutput781 output781/A vssd vssd vccd vccd la_data_in_mprj[123] sky130_fd_sc_hd__buf_2
XFILLER_43_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput792 output792/A vssd vssd vccd vccd la_data_in_mprj[18] sky130_fd_sc_hd__buf_2
XFILLER_8_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[116\]_B la_buf_enable\[116\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input130_A la_data_out_core[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input228_A la_data_out_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2319 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_buffers\[7\]_A user_wb_dat_gates\[7\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input597_A mprj_dat_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[85\]_A input115/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[111\] input273/X mprj_logic_high_inst/HI[441] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[111\]/B sky130_fd_sc_hd__and2_1
XFILLER_11_951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_clk_buf_A _391_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[30\]_TE mprj_adr_buf\[30\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[117\] user_to_mprj_in_gates\[117\]/Y vssd vssd vccd vccd
+ output774/A sky130_fd_sc_hd__inv_2
XFILLER_38_804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[107\]_B la_buf_enable\[107\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[83\] user_to_mprj_in_gates\[83\]/Y vssd vssd vccd vccd output864/A
+ sky130_fd_sc_hd__clkinv_2
XFILLER_24_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output983_A output983/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_A input105/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[4\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput509 la_oenb_mprj[94] vssd vssd vccd vccd _357_/A sky130_fd_sc_hd__buf_2
XFILLER_9_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[4\]_B user_to_mprj_in_gates\[4\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1716 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output1080_A output1080/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[19\] input298/X mprj_logic_high_inst/HI[349] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[19\]/B sky130_fd_sc_hd__and2_1
XFILLER_51_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[67\]_A input95/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input178_A la_data_out_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[41\]_A_N _633_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input345_A la_iena_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input39_A la_data_out_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[56\]_A_N _648_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input512_A la_oenb_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[87\] _551_/Y la_buf\[87\]/TE vssd vssd vccd vccd output740/A sky130_fd_sc_hd__einvp_4
XFILLER_21_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[102\] _365_/A la_buf_enable\[102\]/B vssd vssd vccd vccd la_buf\[102\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_21_1742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1786 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[58\]_A input85/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[24\]_TE la_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output731_A output731/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output829_A output829/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[76\] input105/X user_to_mprj_in_gates\[76\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[76\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_1703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[8\]_A user_to_mprj_in_gates\[8\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_38_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_61 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__634__A _634_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[49\]_A input75/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput306 la_iena_mprj[26] vssd vssd vccd vccd input306/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput317 la_iena_mprj[36] vssd vssd vccd vccd input317/X sky130_fd_sc_hd__clkbuf_1
Xinput339 la_iena_mprj[56] vssd vssd vccd vccd input339/X sky130_fd_sc_hd__clkbuf_1
Xinput328 la_iena_mprj[46] vssd vssd vccd vccd input328/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__544__A _544_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[124\]_A input31/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input295_A la_iena_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[47\]_TE la_buf\[47\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input462_A la_oenb_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_irq_ena_buf\[2\] input626/X user_irq_ena_buf\[2\]/B vssd vssd vccd vccd user_irq_gates\[2\]/B
+ sky130_fd_sc_hd__and2_1
XFILLER_3_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output681_A output681/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[46\] user_to_mprj_in_gates\[46\]/Y vssd vssd vccd vccd output823/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_34_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__454__A _454_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[115\]_A input21/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output779_A output779/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output946_A output946/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__629__A _629_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[102\] input7/X user_to_mprj_in_gates\[102\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[102\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__364__A _364_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_A input11/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_47 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output1043_A output1043/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[86\] input372/X mprj_logic_high_inst/HI[416] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[86\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput125 la_data_out_core[94] vssd vssd vccd vccd input125/X sky130_fd_sc_hd__buf_4
Xinput114 la_data_out_core[84] vssd vssd vccd vccd input114/X sky130_fd_sc_hd__buf_4
Xinput103 la_data_out_core[74] vssd vssd vccd vccd input103/X sky130_fd_sc_hd__buf_4
Xoutput1091 output1091/A vssd vssd vccd vccd mprj_dat_o_user[22] sky130_fd_sc_hd__buf_2
Xoutput1080 output1080/A vssd vssd vccd vccd mprj_dat_o_user[12] sky130_fd_sc_hd__buf_2
XFILLER_49_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[112\] _375_/Y mprj_logic_high_inst/HI[314] vssd vssd vccd
+ vccd output897/A sky130_fd_sc_hd__einvp_4
Xinput136 la_data_out_mprj[103] vssd vssd vccd vccd _567_/A sky130_fd_sc_hd__clkbuf_4
Xinput169 la_data_out_mprj[18] vssd vssd vccd vccd _482_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput147 la_data_out_mprj[113] vssd vssd vccd vccd _577_/A sky130_fd_sc_hd__clkbuf_4
Xinput158 la_data_out_mprj[123] vssd vssd vccd vccd _587_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_641_ _641_/A vssd vssd vccd vccd _641_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[42\] _634_/Y mprj_logic_high_inst/HI[244] vssd vssd vccd
+ vccd output947/A sky130_fd_sc_hd__einvp_2
Xla_buf_enable\[64\] _656_/A la_buf_enable\[64\]/B vssd vssd vccd vccd la_buf\[64\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA__539__A _539_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_buffers\[0\] user_irq_gates\[0\]/Y vssd vssd vccd vccd output1121/A sky130_fd_sc_hd__clkinv_4
XFILLER_44_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_572_ _572_/A vssd vssd vccd vccd _572_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input210_A la_data_out_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input308_A la_iena_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1532 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[19\]_TE mprj_dat_buf\[19\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[106\] _570_/Y la_buf\[106\]/TE vssd vssd vccd vccd output634/A sky130_fd_sc_hd__einvp_8
XFILLER_45_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__449__A _449_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output896_A output896/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[39\] input64/X user_to_mprj_in_gates\[39\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[39\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_82 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[4\]_B la_buf_enable\[4\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__359__A _359_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1352 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input258_A la_data_out_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input160_A la_data_out_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[119\]_A input281/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input425_A la_oenb_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input21_A la_data_out_core[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[120\]_TE mprj_logic_high_inst/HI[322] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_624_ _624_/A vssd vssd vccd vccd _624_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_17_445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_555_ _555_/A vssd vssd vccd vccd _555_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_33_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_486_ _486_/A vssd vssd vccd vccd _486_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_51_2030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_we_buf _395_/Y mprj_we_buf/TE vssd vssd vccd vccd output1114/A sky130_fd_sc_hd__einvp_8
XFILLER_18_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[50\]_A input333/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output644_A output644/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_pwrgood mprj_pwrgood/A vssd vssd vccd vccd output1115/A sky130_fd_sc_hd__buf_8
XANTENNA_output811_A output811/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output909_A output909/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[41\]_A input323/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__642__A _642_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput930 output930/A vssd vssd vccd vccd la_oenb_core[27] sky130_fd_sc_hd__buf_2
Xoutput941 output941/A vssd vssd vccd vccd la_oenb_core[37] sky130_fd_sc_hd__buf_2
Xoutput963 output963/A vssd vssd vccd vccd la_oenb_core[57] sky130_fd_sc_hd__buf_2
Xoutput952 output952/A vssd vssd vccd vccd la_oenb_core[47] sky130_fd_sc_hd__buf_2
Xoutput985 output985/A vssd vssd vccd vccd la_oenb_core[77] sky130_fd_sc_hd__buf_2
Xoutput996 output996/A vssd vssd vccd vccd la_oenb_core[87] sky130_fd_sc_hd__buf_2
Xoutput974 output974/A vssd vssd vccd vccd la_oenb_core[67] sky130_fd_sc_hd__buf_2
XFILLER_43_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output1006_A output1006/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[49\] input331/X mprj_logic_high_inst/HI[379] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[49\]/B sky130_fd_sc_hd__and2_1
XFILLER_2_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_340_ _340_/A vssd vssd vccd vccd _340_/Y sky130_fd_sc_hd__inv_2
XTAP_1658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[32\]_A input313/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[27\] _619_/A la_buf_enable\[27\]/B vssd vssd vccd vccd la_buf\[27\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_35_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__552__A _552_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input375_A la_iena_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input69_A la_data_out_core[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[99\]_A input386/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input542_A mprj_adr_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[42\]_TE mprj_logic_high_inst/HI[244] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_607_ _607_/A vssd vssd vccd vccd _607_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_17_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_538_ _538_/A vssd vssd vccd vccd _538_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_ena_buf\[23\]_A input303/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_469_ _469_/A vssd vssd vccd vccd _469_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__462__A _462_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output859_A output859/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output761_A output761/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[118\]_TE la_buf\[118\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_72 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__637__A _637_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[14\]_A input293/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[94\]_B user_to_mprj_in_gates\[94\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__372__A _372_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[80\]_TE la_buf\[80\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[65\]_TE mprj_logic_high_inst/HI[267] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_7 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output1123_A output1123/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput760 output760/A vssd vssd vccd vccd la_data_in_mprj[104] sky130_fd_sc_hd__buf_2
Xoutput771 output771/A vssd vssd vccd vccd la_data_in_mprj[114] sky130_fd_sc_hd__buf_2
XFILLER_47_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput793 output793/A vssd vssd vccd vccd la_data_in_mprj[19] sky130_fd_sc_hd__buf_2
Xoutput782 output782/A vssd vssd vccd vccd la_data_in_mprj[124] sky130_fd_sc_hd__buf_2
XFILLER_43_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input123_A la_data_out_core[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__547__A _547_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_irq_ena_buf\[1\]_A input625/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_we_buf_A _395_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input492_A la_oenb_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[85\]_B user_to_mprj_in_gates\[85\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[32\] _496_/Y la_buf\[32\]/TE vssd vssd vccd vccd output680/A sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[104\] input265/X mprj_logic_high_inst/HI[434] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[104\]/B sky130_fd_sc_hd__and2_1
Xuser_wb_dat_gates\[4\] input576/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[4\]/Y
+ sky130_fd_sc_hd__nand2_4
XFILLER_52_1490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[70\]_A user_to_mprj_in_gates\[70\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[76\] user_to_mprj_in_gates\[76\]/Y vssd vssd vccd vccd output856/A
+ sky130_fd_sc_hd__inv_2
XFILLER_4_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__457__A _457_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output976_A output976/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[21\] input45/X user_to_mprj_in_gates\[21\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[21\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[76\]_B user_to_mprj_in_gates\[76\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[88\]_TE mprj_logic_high_inst/HI[290] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[31\] user_wb_dat_gates\[31\]/Y vssd vssd vccd vccd output1069/A
+ sky130_fd_sc_hd__inv_6
XFILLER_44_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[9\] _441_/Y mprj_dat_buf\[9\]/TE vssd vssd vccd vccd output1108/A sky130_fd_sc_hd__einvp_8
XFILLER_9_1520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[61\]_A user_to_mprj_in_gates\[61\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__367__A _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[67\]_B user_to_mprj_in_gates\[67\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1073_A output1073/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[72\] _335_/Y mprj_logic_high_inst/HI[274] vssd vssd vccd
+ vccd output980/A sky130_fd_sc_hd__einvp_4
Xla_buf_enable\[94\] _357_/A la_buf_enable\[94\]/B vssd vssd vccd vccd la_buf\[94\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_47_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[20\] _452_/Y mprj_dat_buf\[20\]/TE vssd vssd vccd vccd output1089/A
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input338_A la_iena_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input240_A la_data_out_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[52\]_A user_to_mprj_in_gates\[52\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input505_A la_oenb_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[58\]_B user_to_mprj_in_gates\[58\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[92\]_A _556_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output724_A output724/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[43\]_A user_to_mprj_in_gates\[43\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_40 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[69\] input97/X user_to_mprj_in_gates\[69\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[69\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_51 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[49\]_B user_to_mprj_in_gates\[49\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[83\]_A _547_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[0\] _592_/A la_buf_enable\[0\]/B vssd vssd vccd vccd la_buf\[0\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA__650__A _650_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput307 la_iena_mprj[27] vssd vssd vccd vccd input307/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput318 la_iena_mprj[37] vssd vssd vccd vccd input318/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_47 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[34\]_A user_to_mprj_in_gates\[34\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xinput329 la_iena_mprj[47] vssd vssd vccd vccd input329/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[31\] input312/X mprj_logic_high_inst/HI[361] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[31\]/B sky130_fd_sc_hd__and2_1
XFILLER_45_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[20\]_TE mprj_adr_buf\[20\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_682 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[74\]_A _538_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[124\]_B user_to_mprj_in_gates\[124\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1878 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input190_A la_data_out_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[92\]_B la_buf_enable\[92\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input288_A la_iena_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__560__A _560_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input455_A la_oenb_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input51_A la_data_out_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input622_A user_irq_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[25\]_A user_to_mprj_in_gates\[25\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[65\]_A _529_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[115\]_B user_to_mprj_in_gates\[115\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[39\] user_to_mprj_in_gates\[39\]/Y vssd vssd vccd vccd output815/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output674_A output674/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[83\]_B la_buf_enable\[83\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output939_A output939/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__470__A _470_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output841_A output841/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[16\]_A user_to_mprj_in_gates\[16\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[24\]_A input566/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__645__A _645_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[119\]_A _583_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[40\]_A_N _632_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[56\]_A _520_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_B user_to_mprj_in_gates\[106\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[55\]_A_N _647_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[74\]_B la_buf_enable\[74\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__380__A _380_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output1036_A output1036/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[79\] input364/X mprj_logic_high_inst/HI[409] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[79\]/B sky130_fd_sc_hd__and2_1
Xinput126 la_data_out_core[95] vssd vssd vccd vccd input126/X sky130_fd_sc_hd__buf_4
Xinput115 la_data_out_core[85] vssd vssd vccd vccd input115/X sky130_fd_sc_hd__buf_4
Xinput104 la_data_out_core[75] vssd vssd vccd vccd input104/X sky130_fd_sc_hd__buf_4
Xoutput1081 output1081/A vssd vssd vccd vccd mprj_dat_o_user[13] sky130_fd_sc_hd__buf_2
Xoutput1092 output1092/A vssd vssd vccd vccd mprj_dat_o_user[23] sky130_fd_sc_hd__buf_2
XFILLER_40_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput1070 output1070/A vssd vssd vccd vccd mprj_dat_i_core[3] sky130_fd_sc_hd__buf_2
XFILLER_40_1404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[105\] _368_/Y mprj_logic_high_inst/HI[307] vssd vssd vccd
+ vccd output889/A sky130_fd_sc_hd__einvp_4
Xinput137 la_data_out_mprj[104] vssd vssd vccd vccd _568_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput148 la_data_out_mprj[114] vssd vssd vccd vccd _578_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput159 la_data_out_mprj[124] vssd vssd vccd vccd _588_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_wb_dat_gates\[15\]_A input556/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_640_ _640_/A vssd vssd vccd vccd _640_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[57\] _649_/A la_buf_enable\[57\]/B vssd vssd vccd vccd la_buf\[57\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_44_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_571_ _571_/A vssd vssd vccd vccd _571_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[35\] _627_/Y mprj_logic_high_inst/HI[237] vssd vssd vccd
+ vccd output939/A sky130_fd_sc_hd__einvp_2
XFILLER_5_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[14\]_TE la_buf\[14\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input203_A la_data_out_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__555__A _555_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input99_A la_data_out_core[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[47\]_A _511_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input572_A mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[65\]_B la_buf_enable\[65\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_81 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output791_A output791/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output889_A output889/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__465__A _465_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[38\]_A _502_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[56\]_B la_buf_enable\[56\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[123\]_A _386_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[37\]_TE la_buf\[37\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__375__A _375_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1842 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[29\]_A _493_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_858 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[47\]_B la_buf_enable\[47\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[114\]_A _377_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_578 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input153_A la_data_out_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[119\]_B mprj_logic_high_inst/HI[449] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input320_A la_iena_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_623_ _623_/A vssd vssd vccd vccd _623_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_24_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input418_A la_oenb_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input14_A la_data_out_core[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[62\] _526_/Y la_buf\[62\]/TE vssd vssd vccd vccd output713/A sky130_fd_sc_hd__einvp_8
XFILLER_2_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_554_ _554_/A vssd vssd vccd vccd _554_/Y sky130_fd_sc_hd__inv_2
X_485_ _485_/A vssd vssd vccd vccd _485_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[5\]_TE la_buf\[5\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[50\]_B mprj_logic_high_inst/HI[380] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[38\]_B la_buf_enable\[38\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[26\] _426_/Y mprj_adr_buf\[26\]/TE vssd vssd vccd vccd output1030/A
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[7\]_A input365/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output637_A output637/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[40\]_A _632_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[105\]_A _368_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output804_A output804/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput490 la_oenb_mprj[77] vssd vssd vccd vccd _340_/A sky130_fd_sc_hd__buf_2
Xuser_to_mprj_in_gates\[51\] input78/X user_to_mprj_in_gates\[51\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[51\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[41\]_B mprj_logic_high_inst/HI[371] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_23_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[29\]_B la_buf_enable\[29\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput920 output920/A vssd vssd vccd vccd la_oenb_core[18] sky130_fd_sc_hd__buf_2
XFILLER_2_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput953 output953/A vssd vssd vccd vccd la_oenb_core[48] sky130_fd_sc_hd__buf_2
Xoutput964 output964/A vssd vssd vccd vccd la_oenb_core[58] sky130_fd_sc_hd__buf_2
Xoutput942 output942/A vssd vssd vccd vccd la_oenb_core[38] sky130_fd_sc_hd__buf_2
Xoutput931 output931/A vssd vssd vccd vccd la_oenb_core[28] sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_oen_buffers\[31\]_A _623_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput997 output997/A vssd vssd vccd vccd la_oenb_core[88] sky130_fd_sc_hd__buf_2
Xoutput986 output986/A vssd vssd vccd vccd la_oenb_core[78] sky130_fd_sc_hd__buf_2
Xoutput975 output975/A vssd vssd vccd vccd la_oenb_core[68] sky130_fd_sc_hd__buf_2
XFILLER_28_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input6_A la_data_out_core[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[98\]_A _361_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_298 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[32\]_B mprj_logic_high_inst/HI[362] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_41_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input368_A la_iena_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input270_A la_iena_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[22\]_A _614_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[99\]_B mprj_logic_high_inst/HI[429] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input535_A mprj_adr_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[125\] _388_/A la_buf_enable\[125\]/B vssd vssd vccd vccd la_buf\[125\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_8_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[89\]_A _352_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_606_ _606_/A vssd vssd vccd vccd _606_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_537_ _537_/A vssd vssd vccd vccd _537_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[23\]_B mprj_logic_high_inst/HI[353] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_468_ _468_/A vssd vssd vccd vccd _468_/Y sky130_fd_sc_hd__clkinv_2
X_399_ _399_/A vssd vssd vccd vccd _399_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[21\] user_to_mprj_in_gates\[21\]/Y vssd vssd vccd vccd output796/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_9_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output754_A output754/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output921_A output921/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[13\]_A _605_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[99\] input130/X user_to_mprj_in_gates\[99\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[99\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_1674 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[14\]_B mprj_logic_high_inst/HI[344] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_23_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__653__A _653_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[7\]_A input579/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[110\]_TE mprj_logic_high_inst/HI[312] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput750 output750/A vssd vssd vccd vccd la_data_in_core[96] sky130_fd_sc_hd__buf_2
Xoutput761 output761/A vssd vssd vccd vccd la_data_in_mprj[105] sky130_fd_sc_hd__buf_2
Xoutput772 output772/A vssd vssd vccd vccd la_data_in_mprj[115] sky130_fd_sc_hd__buf_2
XFILLER_47_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput794 output794/A vssd vssd vccd vccd la_data_in_mprj[1] sky130_fd_sc_hd__buf_2
Xoutput783 output783/A vssd vssd vccd vccd la_data_in_mprj[125] sky130_fd_sc_hd__buf_2
XANTENNA_output1116_A output1116/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[61\] input345/X mprj_logic_high_inst/HI[391] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[61\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[7\]_A input109/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input116_A la_data_out_core[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_irq_ena_buf\[1\]_B user_irq_ena_buf\[1\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__563__A _563_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input81_A la_data_out_core[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input485_A la_oenb_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[25\] _489_/Y la_buf\[25\]/TE vssd vssd vccd vccd output672/A sky130_fd_sc_hd__einvp_8
XFILLER_6_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_319 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[69\] user_to_mprj_in_gates\[69\]/Y vssd vssd vccd vccd output848/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_45_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1954 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output871_A output871/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output969_A output969/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[27\] input569/X repeater1125/X vssd vssd vccd vccd user_wb_dat_gates\[27\]/Y
+ sky130_fd_sc_hd__nand2_8
XTAP_1990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__473__A _473_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[14\] input37/X user_to_mprj_in_gates\[14\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[14\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_1277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[24\] user_wb_dat_gates\[24\]/Y vssd vssd vccd vccd output1061/A
+ sky130_fd_sc_hd__inv_6
XFILLER_29_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[125\] input32/X user_to_mprj_in_gates\[125\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[125\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA__648__A _648_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[31\]_A _463_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__383__A _383_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[32\]_TE mprj_logic_high_inst/HI[234] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1066_A output1066/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[65\] _657_/Y mprj_logic_high_inst/HI[267] vssd vssd vccd
+ vccd output972/A sky130_fd_sc_hd__einvp_8
XFILLER_43_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[87\] _350_/A la_buf_enable\[87\]/B vssd vssd vccd vccd la_buf\[87\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_43_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[13\] _445_/Y mprj_dat_buf\[13\]/TE vssd vssd vccd vccd output1081/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_19_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input233_A la_data_out_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__558__A _558_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[108\]_TE la_buf\[108\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input400_A la_oenb_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[22\]_A _454_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[7\]_TE mprj_adr_buf\[7\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[122\] user_to_mprj_in_gates\[122\]/Y vssd vssd vccd vccd
+ output780/A sky130_fd_sc_hd__inv_2
XFILLER_26_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output717_A output717/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__468__A _468_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2080 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[70\]_TE la_buf\[70\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[13\]_A _445_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[20\]_A user_wb_dat_gates\[20\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[55\]_TE mprj_logic_high_inst/HI[257] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput308 la_iena_mprj[28] vssd vssd vccd vccd input308/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput319 la_iena_mprj[38] vssd vssd vccd vccd input319/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__378__A _378_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[8\]_A _600_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_buffers\[11\]_A user_wb_dat_gates\[11\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_24_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[24\] input304/X mprj_logic_high_inst/HI[354] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[24\]/B sky130_fd_sc_hd__and2_1
XFILLER_12_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input183_A la_data_out_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input448_A la_oenb_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input350_A la_iena_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input44_A la_data_out_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[92\] _556_/Y la_buf\[92\]/TE vssd vssd vccd vccd output746/A sky130_fd_sc_hd__einvp_4
XFILLER_19_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[93\]_TE la_buf\[93\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input615_A mprj_sel_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[78\]_TE mprj_logic_high_inst/HI[280] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_vdd_pwrgood mprj_vdd_pwrgood/A vssd vssd vccd vccd output1116/A sky130_fd_sc_hd__buf_6
XFILLER_31_812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output667_A output667/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output834_A output834/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[81\] input111/X user_to_mprj_in_gates\[81\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[81\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[24\]_B repeater1125/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_458 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output1029_A output1029/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput1060 output1060/A vssd vssd vccd vccd mprj_dat_i_core[23] sky130_fd_sc_hd__buf_2
Xinput127 la_data_out_core[96] vssd vssd vccd vccd input127/X sky130_fd_sc_hd__buf_4
Xinput116 la_data_out_core[86] vssd vssd vccd vccd input116/X sky130_fd_sc_hd__buf_4
Xinput105 la_data_out_core[76] vssd vssd vccd vccd input105/X sky130_fd_sc_hd__buf_4
Xoutput1093 output1093/A vssd vssd vccd vccd mprj_dat_o_user[24] sky130_fd_sc_hd__buf_2
Xoutput1082 output1082/A vssd vssd vccd vccd mprj_dat_o_user[14] sky130_fd_sc_hd__buf_2
XFILLER_49_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput1071 output1071/A vssd vssd vccd vccd mprj_dat_i_core[4] sky130_fd_sc_hd__buf_2
Xinput138 la_data_out_mprj[105] vssd vssd vccd vccd _569_/A sky130_fd_sc_hd__clkbuf_2
Xinput149 la_data_out_mprj[115] vssd vssd vccd vccd _579_/A sky130_fd_sc_hd__buf_2
XFILLER_45_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[9\]_A_N _601_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[15\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_570_ _570_/A vssd vssd vccd vccd _570_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[28\] _620_/Y mprj_logic_high_inst/HI[230] vssd vssd vccd
+ vccd output931/A sky130_fd_sc_hd__einvp_2
XPHY_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[0\]_A _464_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input398_A la_oenb_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__571__A _571_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input565_A mprj_dat_i_user[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[3\] _467_/Y la_buf\[3\]/TE vssd vssd vccd vccd output688/A sky130_fd_sc_hd__einvp_8
XFILLER_49_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_gates\[0\]_A input621/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[0\] _400_/Y mprj_adr_buf\[0\]/TE vssd vssd vccd vccd output1012/A sky130_fd_sc_hd__einvp_4
XFILLER_7_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[51\] user_to_mprj_in_gates\[51\]/Y vssd vssd vccd vccd output829/A
+ sky130_fd_sc_hd__clkinv_4
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output784_A output784/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output951_A output951/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__481__A _481_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_73 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[10\]_TE mprj_adr_buf\[10\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__656__A _656_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[7\]_A _407_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__391__A _391_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[91\] input378/X mprj_logic_high_inst/HI[421] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[91\]/B sky130_fd_sc_hd__and2_1
XFILLER_49_517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input146_A la_data_out_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_622_ _622_/A vssd vssd vccd vccd _622_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_1809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__566__A _566_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input313_A la_iena_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_553_ _553_/A vssd vssd vccd vccd _553_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_53_2308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[55\] _519_/Y la_buf\[55\]/TE vssd vssd vccd vccd output705/A sky130_fd_sc_hd__einvp_8
XFILLER_44_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_484_ _484_/A vssd vssd vccd vccd _484_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1618 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1738 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[127\] input290/X mprj_logic_high_inst/HI[457] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[127\]/B sky130_fd_sc_hd__and2_1
XFILLER_51_2054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[7\]_B mprj_logic_high_inst/HI[337] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[19\] _419_/Y mprj_adr_buf\[19\]/TE vssd vssd vccd vccd output1022/A
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[111\] _575_/Y la_buf\[111\]/TE vssd vssd vccd vccd output640/A sky130_fd_sc_hd__einvp_2
XFILLER_29_1823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[99\] user_to_mprj_in_gates\[99\]/Y vssd vssd vccd vccd output881/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_7_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput480 la_oenb_mprj[68] vssd vssd vccd vccd _331_/A sky130_fd_sc_hd__clkbuf_2
Xinput491 la_oenb_mprj[78] vssd vssd vccd vccd _341_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[54\]_A_N _646_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__476__A _476_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output999_A output999/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[9\] user_wb_dat_gates\[9\]/Y vssd vssd vccd vccd output1076/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_35_255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[44\] input70/X user_to_mprj_in_gates\[44\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[44\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[69\]_A_N _332_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput910 output910/A vssd vssd vccd vccd la_oenb_core[124] sky130_fd_sc_hd__buf_2
Xoutput921 output921/A vssd vssd vccd vccd la_oenb_core[19] sky130_fd_sc_hd__buf_2
XFILLER_28_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput943 output943/A vssd vssd vccd vccd la_oenb_core[39] sky130_fd_sc_hd__buf_2
Xoutput932 output932/A vssd vssd vccd vccd la_oenb_core[29] sky130_fd_sc_hd__buf_2
Xoutput954 output954/A vssd vssd vccd vccd la_oenb_core[49] sky130_fd_sc_hd__buf_2
XFILLER_28_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[6\] input98/X user_to_mprj_in_gates\[6\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[6\]/Y sky130_fd_sc_hd__nand2_2
Xoutput987 output987/A vssd vssd vccd vccd la_oenb_core[79] sky130_fd_sc_hd__buf_2
Xoutput976 output976/A vssd vssd vccd vccd la_oenb_core[69] sky130_fd_sc_hd__buf_2
Xoutput965 output965/A vssd vssd vccd vccd la_oenb_core[59] sky130_fd_sc_hd__buf_2
XFILLER_28_1333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[30\]_A input55/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput998 output998/A vssd vssd vccd vccd la_oenb_core[89] sky130_fd_sc_hd__buf_2
XTAP_450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__386__A _386_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1096_A output1096/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_A input128/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1684 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[95\] _358_/Y mprj_logic_high_inst/HI[297] vssd vssd vccd
+ vccd output1005/A sky130_fd_sc_hd__einvp_4
XFILLER_5_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_822 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input263_A la_iena_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[21\]_A input45/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[119\]_B la_buf_enable\[119\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input430_A la_oenb_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input528_A mprj_adr_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[8\] input376/X mprj_logic_high_inst/HI[338] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[8\]/B sky130_fd_sc_hd__and2_1
Xla_buf_enable\[118\] _381_/A la_buf_enable\[118\]/B vssd vssd vccd vccd la_buf\[118\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_24_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_605_ _605_/A vssd vssd vccd vccd _605_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_70 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_536_ _536_/A vssd vssd vccd vccd _536_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_33_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[88\]_A input118/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_467_ _467_/A vssd vssd vccd vccd _467_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_18_1579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_398_ _398_/A vssd vssd vccd vccd _398_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1768 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[27\]_TE la_buf\[27\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[14\] user_to_mprj_in_gates\[14\]/Y vssd vssd vccd vccd output788/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output747_A output747/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output914_A output914/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[12\]_A input35/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[79\]_A input108/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[7\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput751 output751/A vssd vssd vccd vccd la_data_in_core[97] sky130_fd_sc_hd__buf_2
Xoutput740 output740/A vssd vssd vccd vccd la_data_in_core[87] sky130_fd_sc_hd__buf_2
Xoutput762 output762/A vssd vssd vccd vccd la_data_in_mprj[106] sky130_fd_sc_hd__buf_2
Xoutput795 output795/A vssd vssd vccd vccd la_data_in_mprj[20] sky130_fd_sc_hd__buf_2
Xoutput773 output773/A vssd vssd vccd vccd la_data_in_mprj[116] sky130_fd_sc_hd__buf_2
Xoutput784 output784/A vssd vssd vccd vccd la_data_in_mprj[126] sky130_fd_sc_hd__buf_2
XFILLER_43_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output1011_A output1011/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1109_A output1109/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[7\]_B user_to_mprj_in_gates\[7\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[54\] input337/X mprj_logic_high_inst/HI[384] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[54\]/B sky130_fd_sc_hd__and2_1
XFILLER_41_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input109_A la_data_out_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[10\] _602_/Y mprj_logic_high_inst/HI[212] vssd vssd vccd
+ vccd output894/A sky130_fd_sc_hd__einvp_4
XTAP_1435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[32\] _624_/A la_buf_enable\[32\]/B vssd vssd vccd vccd la_buf\[32\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_in_buffers\[6\] user_to_mprj_in_gates\[6\]/Y vssd vssd vccd vccd output849/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_35_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input478_A la_oenb_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input380_A la_iena_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input74_A la_data_out_core[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[18\] _482_/Y la_buf\[18\]/TE vssd vssd vccd vccd output664/A sky130_fd_sc_hd__einvp_8
XFILLER_6_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output697_A output697/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_519_ _519_/A vssd vssd vccd vccd _519_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_33_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output864_A output864/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_buffers\[17\] user_wb_dat_gates\[17\]/Y vssd vssd vccd vccd output1053/A
+ sky130_fd_sc_hd__inv_6
XFILLER_25_2037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[118\] input24/X user_to_mprj_in_gates\[118\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[118\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1059_A output1059/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[58\] _650_/Y mprj_logic_high_inst/HI[260] vssd vssd vccd
+ vccd output964/A sky130_fd_sc_hd__einvp_8
XFILLER_43_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input226_A la_data_out_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__574__A _574_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[127\]_A input34/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[100\]_A input261/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input595_A mprj_dat_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[115\] user_to_mprj_in_gates\[115\]/Y vssd vssd vccd vccd
+ output772/A sky130_fd_sc_hd__clkinv_4
XFILLER_26_1667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[81\] user_to_mprj_in_gates\[81\]/Y vssd vssd vccd vccd output862/A
+ sky130_fd_sc_hd__inv_2
XFILLER_37_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_97 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_75 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output981_A output981/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[100\]_TE mprj_logic_high_inst/HI[302] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__484__A _484_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_A input24/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput309 la_iena_mprj[29] vssd vssd vccd vccd input309/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[109\]_A input14/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__394__A _394_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[17\] input296/X mprj_logic_high_inst/HI[347] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[17\]/B sky130_fd_sc_hd__and2_1
XFILLER_16_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input176_A la_data_out_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input343_A la_iena_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input37_A la_data_out_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__569__A _569_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[123\]_TE mprj_logic_high_inst/HI[325] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[85\] _549_/Y la_buf\[85\]/TE vssd vssd vccd vccd output738/A sky130_fd_sc_hd__einvp_4
XANTENNA_input510_A la_oenb_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input608_A mprj_dat_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[100\] _363_/A la_buf_enable\[100\]/B vssd vssd vccd vccd la_buf\[100\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_21_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[80\]_A input366/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output827_A output827/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__479__A _479_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[74\] input103/X user_to_mprj_in_gates\[74\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[74\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[22\]_TE mprj_logic_high_inst/HI[224] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[71\]_A input356/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[7\]_B la_buf_enable\[7\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput1050 output1050/A vssd vssd vccd vccd mprj_dat_i_core[14] sky130_fd_sc_hd__buf_2
Xinput117 la_data_out_core[87] vssd vssd vccd vccd input117/X sky130_fd_sc_hd__buf_4
Xinput106 la_data_out_core[77] vssd vssd vccd vccd input106/X sky130_fd_sc_hd__buf_4
Xoutput1094 output1094/A vssd vssd vccd vccd mprj_dat_o_user[25] sky130_fd_sc_hd__buf_2
Xoutput1083 output1083/A vssd vssd vccd vccd mprj_dat_o_user[15] sky130_fd_sc_hd__buf_2
XANTENNA__389__A _389_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput1072 output1072/A vssd vssd vccd vccd mprj_dat_i_core[5] sky130_fd_sc_hd__buf_2
Xoutput1061 output1061/A vssd vssd vccd vccd mprj_dat_i_core[24] sky130_fd_sc_hd__buf_2
Xinput128 la_data_out_core[97] vssd vssd vccd vccd input128/X sky130_fd_sc_hd__buf_4
XFILLER_44_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput139 la_data_out_mprj[106] vssd vssd vccd vccd _570_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[62\]_A input346/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_828 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input293_A la_iena_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input558_A mprj_dat_i_user[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input460_A la_oenb_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[60\]_TE la_buf\[60\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_irq_ena_buf\[0\] input624/X user_irq_ena_buf\[0\]/B vssd vssd vccd vccd user_irq_gates\[0\]/B
+ sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[45\]_TE mprj_logic_high_inst/HI[247] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_gates\[0\]_B user_irq_gates\[0\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[53\]_A input336/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1488 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[44\] user_to_mprj_in_gates\[44\]/Y vssd vssd vccd vccd output821/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output777_A output777/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output944_A output944/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_96 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1344 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_sel_buf\[1\]_A _397_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[100\] input5/X user_to_mprj_in_gates\[100\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[100\]/Y sky130_fd_sc_hd__nand2_1
XTAP_1809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[44\]_A input326/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[83\]_TE la_buf\[83\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[68\]_TE mprj_logic_high_inst/HI[270] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1041_A output1041/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[84\] input370/X mprj_logic_high_inst/HI[414] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[84\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[110\] _373_/Y mprj_logic_high_inst/HI[312] vssd vssd vccd
+ vccd output895/A sky130_fd_sc_hd__einvp_2
XFILLER_40_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[40\] _632_/Y mprj_logic_high_inst/HI[242] vssd vssd vccd
+ vccd output945/A sky130_fd_sc_hd__einvp_2
Xla_buf_enable\[62\] _654_/A la_buf_enable\[62\]/B vssd vssd vccd vccd la_buf\[62\]/TE
+ sky130_fd_sc_hd__and2b_1
X_621_ _621_/A vssd vssd vccd vccd _621_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input139_A la_data_out_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_552_ _552_/A vssd vssd vccd vccd _552_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[35\]_A input316/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input306_A la_iena_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_483_ _483_/A vssd vssd vccd vccd _483_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__582__A _582_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[48\] _512_/Y la_buf\[48\]/TE vssd vssd vccd vccd output697/A sky130_fd_sc_hd__einvp_8
XFILLER_51_2077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_82 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[2\]_A _434_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[104\] _568_/Y la_buf\[104\]/TE vssd vssd vccd vccd output632/A sky130_fd_sc_hd__einvp_8
XFILLER_7_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput470 la_oenb_mprj[59] vssd vssd vccd vccd _651_/A sky130_fd_sc_hd__buf_2
Xinput481 la_oenb_mprj[69] vssd vssd vccd vccd _332_/A sky130_fd_sc_hd__buf_2
XFILLER_3_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput492 la_oenb_mprj[79] vssd vssd vccd vccd _342_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_output894_A output894/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[26\]_A input306/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[37\] input62/X user_to_mprj_in_gates\[37\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[37\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__492__A _492_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[8\]_A_N _600_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput911 output911/A vssd vssd vccd vccd la_oenb_core[125] sky130_fd_sc_hd__buf_2
Xoutput900 output900/A vssd vssd vccd vccd la_oenb_core[115] sky130_fd_sc_hd__buf_2
XFILLER_28_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput955 output955/A vssd vssd vccd vccd la_oenb_core[4] sky130_fd_sc_hd__buf_2
Xoutput933 output933/A vssd vssd vccd vccd la_oenb_core[2] sky130_fd_sc_hd__buf_2
Xoutput944 output944/A vssd vssd vccd vccd la_oenb_core[3] sky130_fd_sc_hd__buf_2
Xoutput922 output922/A vssd vssd vccd vccd la_oenb_core[1] sky130_fd_sc_hd__buf_2
Xoutput988 output988/A vssd vssd vccd vccd la_oenb_core[7] sky130_fd_sc_hd__buf_2
Xoutput977 output977/A vssd vssd vccd vccd la_oenb_core[6] sky130_fd_sc_hd__buf_2
Xoutput966 output966/A vssd vssd vccd vccd la_oenb_core[5] sky130_fd_sc_hd__buf_2
XFILLER_28_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[30\]_B user_to_mprj_in_gates\[30\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[91\]_A user_to_mprj_in_gates\[91\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xoutput999 output999/A vssd vssd vccd vccd la_oenb_core[8] sky130_fd_sc_hd__buf_2
XTAP_440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[17\]_A input296/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_B user_to_mprj_in_gates\[97\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1089_A output1089/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[88\] _351_/Y mprj_logic_high_inst/HI[290] vssd vssd vccd
+ vccd output997/A sky130_fd_sc_hd__einvp_2
XFILLER_11_1371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[21\]_B user_to_mprj_in_gates\[21\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input256_A la_data_out_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[82\]_A user_to_mprj_in_gates\[82\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_49_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__577__A _577_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input423_A la_oenb_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_604_ _604_/A vssd vssd vccd vccd _604_/Y sky130_fd_sc_hd__clkinv_2
X_535_ _535_/A vssd vssd vccd vccd _535_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_716 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[88\]_B user_to_mprj_in_gates\[88\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_466_ _466_/A vssd vssd vccd vccd _466_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_43_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_397_ _397_/A vssd vssd vccd vccd _397_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[31\] _431_/Y mprj_adr_buf\[31\]/TE vssd vssd vccd vccd output1036/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[120\]_A user_to_mprj_in_gates\[120\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output642_A output642/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[12\]_B user_to_mprj_in_gates\[12\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[73\]_A user_to_mprj_in_gates\[73\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output907_A output907/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__487__A _487_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[79\]_B user_to_mprj_in_gates\[79\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[111\]_A user_to_mprj_in_gates\[111\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xoutput730 output730/A vssd vssd vccd vccd la_data_in_core[78] sky130_fd_sc_hd__buf_2
XFILLER_30_1279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[100\]_A _564_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput752 output752/A vssd vssd vccd vccd la_data_in_core[98] sky130_fd_sc_hd__buf_2
Xoutput741 output741/A vssd vssd vccd vccd la_data_in_core[88] sky130_fd_sc_hd__buf_2
Xoutput763 output763/A vssd vssd vccd vccd la_data_in_mprj[107] sky130_fd_sc_hd__buf_2
XFILLER_48_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput796 output796/A vssd vssd vccd vccd la_data_in_mprj[21] sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_buffers\[64\]_A user_to_mprj_in_gates\[64\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput774 output774/A vssd vssd vccd vccd la_data_in_mprj[117] sky130_fd_sc_hd__buf_2
Xoutput785 output785/A vssd vssd vccd vccd la_data_in_mprj[127] sky130_fd_sc_hd__buf_2
XFILLER_46_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__397__A _397_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1004_A output1004/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[47\] input329/X mprj_logic_high_inst/HI[377] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[47\]/B sky130_fd_sc_hd__and2_1
XTAP_2126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[23\]_TE mprj_adr_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[25\] _617_/A la_buf_enable\[25\]/B vssd vssd vccd vccd la_buf\[25\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_35_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[53\]_A_N _645_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input373_A la_iena_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[102\]_A user_to_mprj_in_gates\[102\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input67_A la_data_out_core[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input540_A mprj_adr_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[55\]_A user_to_mprj_in_gates\[55\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[68\]_A_N _331_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_518_ _518_/A vssd vssd vccd vccd _518_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[95\]_A _559_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_449_ _449_/A vssd vssd vccd vccd _449_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_31_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output857_A output857/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[46\]_A user_to_mprj_in_gates\[46\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_822 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[86\]_A _550_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1606 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output1121_A output1121/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[37\]_A user_to_mprj_in_gates\[37\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[10\]_A _474_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input121_A la_data_out_core[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[17\]_TE la_buf\[17\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input219_A la_data_out_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[77\]_A _541_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[127\]_B user_to_mprj_in_gates\[127\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_42_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input490_A la_oenb_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[100\]_B mprj_logic_high_inst/HI[430] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[95\]_B la_buf_enable\[95\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input588_A mprj_dat_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__590__A _590_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[30\] _494_/Y la_buf\[30\]/TE vssd vssd vccd vccd output678/A sky130_fd_sc_hd__einvp_8
XFILLER_7_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[102\] input263/X mprj_logic_high_inst/HI[432] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[102\]/B sky130_fd_sc_hd__and2_1
Xuser_wb_dat_gates\[2\] input572/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[2\]/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_32_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[28\]_A user_to_mprj_in_gates\[28\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[108\] user_to_mprj_in_gates\[108\]/Y vssd vssd vccd vccd
+ output764/A sky130_fd_sc_hd__inv_2
XFILLER_6_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_43 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[74\] user_to_mprj_in_gates\[74\]/Y vssd vssd vccd vccd output854/A
+ sky130_fd_sc_hd__clkinv_2
XFILLER_4_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[118\]_B user_to_mprj_in_gates\[118\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output974_A output974/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[68\]_A _532_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[86\]_B la_buf_enable\[86\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[19\]_A user_to_mprj_in_gates\[19\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[7\] _439_/Y mprj_dat_buf\[7\]/TE vssd vssd vccd vccd output1106/A sky130_fd_sc_hd__einvp_8
XANTENNA_user_wb_dat_gates\[27\]_A input569/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[10\]_B la_buf_enable\[10\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[109\]_B user_to_mprj_in_gates\[109\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_51_173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[59\]_A _523_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[77\]_B la_buf_enable\[77\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1071_A output1071/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input169_A la_data_out_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[70\] _333_/Y mprj_logic_high_inst/HI[272] vssd vssd vccd
+ vccd output978/A sky130_fd_sc_hd__einvp_4
XFILLER_27_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[92\] _355_/A la_buf_enable\[92\]/B vssd vssd vccd vccd la_buf\[92\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_47_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[18\]_A input559/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input336_A la_iena_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[78\] _542_/Y la_buf\[78\]/TE vssd vssd vccd vccd output730/A sky130_fd_sc_hd__einvp_4
XANTENNA_input503_A la_oenb_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__585__A _585_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[8\]_TE la_buf\[8\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[80\]_B mprj_logic_high_inst/HI[410] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_43_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[68\]_B la_buf_enable\[68\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[70\]_A _333_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output722_A output722/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[67\] input95/X user_to_mprj_in_gates\[67\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[67\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__495__A _495_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[71\]_B mprj_logic_high_inst/HI[401] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[59\]_B la_buf_enable\[59\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[126\]_A _389_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[61\]_A _653_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput1040 output1040/A vssd vssd vccd vccd mprj_adr_o_user[6] sky130_fd_sc_hd__buf_2
XFILLER_46_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput1051 output1051/A vssd vssd vccd vccd mprj_dat_i_core[15] sky130_fd_sc_hd__buf_2
Xinput118 la_data_out_core[88] vssd vssd vccd vccd input118/X sky130_fd_sc_hd__buf_4
Xinput107 la_data_out_core[78] vssd vssd vccd vccd input107/X sky130_fd_sc_hd__buf_4
Xoutput1084 output1084/A vssd vssd vccd vccd mprj_dat_o_user[16] sky130_fd_sc_hd__buf_2
XFILLER_44_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput1073 output1073/A vssd vssd vccd vccd mprj_dat_i_core[6] sky130_fd_sc_hd__buf_2
Xoutput1062 output1062/A vssd vssd vccd vccd mprj_dat_i_core[25] sky130_fd_sc_hd__buf_2
Xinput129 la_data_out_core[98] vssd vssd vccd vccd input129/X sky130_fd_sc_hd__buf_4
Xoutput1095 output1095/A vssd vssd vccd vccd mprj_dat_o_user[26] sky130_fd_sc_hd__buf_2
XFILLER_44_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[62\]_B mprj_logic_high_inst/HI[392] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_53_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input286_A la_iena_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[117\]_A _380_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[52\]_A _644_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input453_A la_oenb_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input620_A mprj_we_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[53\]_B mprj_logic_high_inst/HI[383] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[37\] user_to_mprj_in_gates\[37\]/Y vssd vssd vccd vccd output813/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output672_A output672/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output937_A output937/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[43\]_A _635_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[108\]_A _371_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[44\]_B mprj_logic_high_inst/HI[374] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_53_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[113\]_TE mprj_logic_high_inst/HI[315] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[34\]_A _626_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1034_A output1034/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_clk_buf_TE mprj_clk_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[77\] input362/X mprj_logic_high_inst/HI[407] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[77\]/B sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[103\] _366_/Y mprj_logic_high_inst/HI[305] vssd vssd vccd
+ vccd output887/A sky130_fd_sc_hd__einvp_4
XFILLER_44_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_620_ _620_/A vssd vssd vccd vccd _620_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_551_ _551_/A vssd vssd vccd vccd _551_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[33\] _625_/Y mprj_logic_high_inst/HI[235] vssd vssd vccd
+ vccd output937/A sky130_fd_sc_hd__einvp_2
XANTENNA_mprj_adr_buf\[30\]_A _430_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[55\] _647_/A la_buf_enable\[55\]/B vssd vssd vccd vccd la_buf\[55\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_33_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[35\]_B mprj_logic_high_inst/HI[365] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_482_ _482_/A vssd vssd vccd vccd _482_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input201_A la_data_out_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_290 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input97_A la_data_out_core[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input570_A mprj_dat_i_user[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[12\]_TE mprj_logic_high_inst/HI[214] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[25\]_A _617_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput482 la_oenb_mprj[6] vssd vssd vccd vccd _598_/A sky130_fd_sc_hd__clkbuf_2
Xinput471 la_oenb_mprj[5] vssd vssd vccd vccd _597_/A sky130_fd_sc_hd__clkbuf_2
Xinput460 la_oenb_mprj[4] vssd vssd vccd vccd _596_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput493 la_oenb_mprj[7] vssd vssd vccd vccd _599_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_mprj_adr_buf\[21\]_A _421_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[26\]_B mprj_logic_high_inst/HI[356] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_51_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output887_A output887/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj2_vdd_pwrgood_A mprj2_vdd_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[16\]_A _608_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput912 output912/A vssd vssd vccd vccd la_oenb_core[126] sky130_fd_sc_hd__buf_2
Xoutput901 output901/A vssd vssd vccd vccd la_oenb_core[116] sky130_fd_sc_hd__buf_2
XFILLER_12_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput945 output945/A vssd vssd vccd vccd la_oenb_core[40] sky130_fd_sc_hd__buf_2
Xoutput934 output934/A vssd vssd vccd vccd la_oenb_core[30] sky130_fd_sc_hd__buf_2
Xoutput923 output923/A vssd vssd vccd vccd la_oenb_core[20] sky130_fd_sc_hd__buf_2
XFILLER_47_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput978 output978/A vssd vssd vccd vccd la_oenb_core[70] sky130_fd_sc_hd__buf_2
Xoutput956 output956/A vssd vssd vccd vccd la_oenb_core[50] sky130_fd_sc_hd__buf_2
Xoutput967 output967/A vssd vssd vccd vccd la_oenb_core[60] sky130_fd_sc_hd__buf_2
XFILLER_28_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput989 output989/A vssd vssd vccd vccd la_oenb_core[80] sky130_fd_sc_hd__buf_2
XFILLER_45_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[12\]_A _412_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[17\]_B mprj_logic_high_inst/HI[347] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_42_717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[50\]_TE la_buf\[50\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[35\]_TE mprj_logic_high_inst/HI[237] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[109\]_A_N _372_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[29\] _461_/Y mprj_dat_buf\[29\]/TE vssd vssd vccd vccd output1098/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input151_A la_data_out_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input249_A la_data_out_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_603_ _603_/A vssd vssd vccd vccd _603_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input416_A la_oenb_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input12_A la_data_out_core[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[60\] _524_/Y la_buf\[60\]/TE vssd vssd vccd vccd output711/A sky130_fd_sc_hd__einvp_8
X_534_ _534_/A vssd vssd vccd vccd _534_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__593__A _593_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_465_ _465_/A vssd vssd vccd vccd _465_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_396_ _396_/A vssd vssd vccd vccd _396_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[24\] _424_/Y mprj_adr_buf\[24\]/TE vssd vssd vccd vccd output1028/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_2334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output635_A output635/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output802_A output802/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[73\]_TE la_buf\[73\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput290 la_iena_mprj[127] vssd vssd vccd vccd input290/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[58\]_TE mprj_logic_high_inst/HI[260] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[9\] _601_/A la_buf_enable\[9\]/B vssd vssd vccd vccd la_buf\[9\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput720 output720/A vssd vssd vccd vccd la_data_in_core[69] sky130_fd_sc_hd__buf_2
XFILLER_2_109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput753 output753/A vssd vssd vccd vccd la_data_in_core[99] sky130_fd_sc_hd__buf_2
Xoutput742 output742/A vssd vssd vccd vccd la_data_in_core[89] sky130_fd_sc_hd__buf_2
Xoutput731 output731/A vssd vssd vccd vccd la_data_in_core[79] sky130_fd_sc_hd__buf_2
XFILLER_43_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput786 output786/A vssd vssd vccd vccd la_data_in_mprj[12] sky130_fd_sc_hd__buf_2
Xoutput797 output797/A vssd vssd vccd vccd la_data_in_mprj[22] sky130_fd_sc_hd__buf_2
Xoutput764 output764/A vssd vssd vccd vccd la_data_in_mprj[108] sky130_fd_sc_hd__buf_2
Xoutput775 output775/A vssd vssd vccd vccd la_data_in_mprj[118] sky130_fd_sc_hd__buf_2
XANTENNA_input4_A la_data_out_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_dat_buf\[22\]_TE mprj_dat_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_400 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[18\] _610_/A la_buf_enable\[18\]/B vssd vssd vccd vccd la_buf\[18\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_22_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[1\]_TE mprj_logic_high_inst/HI[203] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input199_A la_data_out_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input366_A la_iena_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_irq_gates\[1\] input622/X user_irq_gates\[1\]/B vssd vssd vccd vccd user_irq_gates\[1\]/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_2_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input533_A mprj_adr_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__588__A _588_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[96\]_TE la_buf\[96\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[123\] _386_/A la_buf_enable\[123\]/B vssd vssd vccd vccd la_buf\[123\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_24_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[25\]_A _457_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[7\]_A_N _599_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_517_ _517_/A vssd vssd vccd vccd _517_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_448_ _448_/A vssd vssd vccd vccd _448_/Y sky130_fd_sc_hd__inv_6
X_379_ _379_/A vssd vssd vccd vccd _379_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output752_A output752/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[97\] input128/X user_to_mprj_in_gates\[97\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[97\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__498__A _498_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[16\]_A _448_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[23\]_A user_wb_dat_gates\[23\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_3_1156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_ack_buffer_A user_wb_ack_gate/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output1114_A output1114/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_buffers\[14\]_A user_wb_dat_gates\[14\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_27_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input114_A la_data_out_core[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input483_A la_oenb_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[23\] _487_/Y la_buf\[23\]/TE vssd vssd vccd vccd output670/A sky130_fd_sc_hd__einvp_8
XFILLER_7_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_11 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[67\] user_to_mprj_in_gates\[67\]/Y vssd vssd vccd vccd output846/A
+ sky130_fd_sc_hd__clkinv_2
XFILLER_45_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output967_A output967/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[25\] input567/X repeater1125/X vssd vssd vccd vccd user_wb_dat_gates\[25\]/Y
+ sky130_fd_sc_hd__nand2_8
XTAP_1790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[12\] input35/X user_to_mprj_in_gates\[12\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[12\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_31_2021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_wb_dat_buffers\[22\] user_wb_dat_gates\[22\]/Y vssd vssd vccd vccd output1059/A
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_mprj_adr_buf\[13\]_TE mprj_adr_buf\[13\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[27\]_B repeater1125/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[123\] input30/X user_to_mprj_in_gates\[123\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[123\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[52\]_A_N _644_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[67\]_A_N _330_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output1064_A output1064/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[0\]_A user_wb_dat_gates\[0\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[63\] _655_/Y mprj_logic_high_inst/HI[265] vssd vssd vccd
+ vccd output970/A sky130_fd_sc_hd__einvp_4
Xla_buf_enable\[85\] _348_/A la_buf_enable\[85\]/B vssd vssd vccd vccd la_buf\[85\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_27_1967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[18\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[11\] _443_/Y mprj_dat_buf\[11\]/TE vssd vssd vccd vccd output1079/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input231_A la_data_out_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[1\]_TE mprj_dat_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input329_A la_iena_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[3\]_A _467_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[100\]_B la_buf_enable\[100\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[121\]_TE la_buf\[121\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[127\] _591_/Y la_buf\[127\]/TE vssd vssd vccd vccd output657/A sky130_fd_sc_hd__einvp_4
XFILLER_10_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[120\] user_to_mprj_in_gates\[120\]/Y vssd vssd vccd vccd
+ output778/A sky130_fd_sc_hd__inv_6
XTAP_826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output715_A output715/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[60\]_A input88/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput1030 output1030/A vssd vssd vccd vccd mprj_adr_o_user[26] sky130_fd_sc_hd__buf_2
Xoutput1041 output1041/A vssd vssd vccd vccd mprj_adr_o_user[7] sky130_fd_sc_hd__buf_2
Xinput108 la_data_out_core[79] vssd vssd vccd vccd input108/X sky130_fd_sc_hd__buf_4
Xoutput1085 output1085/A vssd vssd vccd vccd mprj_dat_o_user[17] sky130_fd_sc_hd__buf_2
XFILLER_44_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput1074 output1074/A vssd vssd vccd vccd mprj_dat_i_core[7] sky130_fd_sc_hd__buf_2
Xoutput1052 output1052/A vssd vssd vccd vccd mprj_dat_i_core[16] sky130_fd_sc_hd__buf_2
Xoutput1063 output1063/A vssd vssd vccd vccd mprj_dat_i_core[26] sky130_fd_sc_hd__buf_2
Xinput119 la_data_out_core[89] vssd vssd vccd vccd input119/X sky130_fd_sc_hd__buf_4
Xoutput1096 output1096/A vssd vssd vccd vccd mprj_dat_o_user[27] sky130_fd_sc_hd__buf_2
XFILLER_44_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2016 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[22\] input302/X mprj_logic_high_inst/HI[352] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[22\]/B sky130_fd_sc_hd__and2_1
XFILLER_12_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input181_A la_data_out_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input279_A la_iena_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[51\]_A input78/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input446_A la_oenb_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input42_A la_data_out_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput620 mprj_we_o_core vssd vssd vccd vccd _395_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__596__A _596_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[90\] _554_/Y la_buf\[90\]/TE vssd vssd vccd vccd output744/A sky130_fd_sc_hd__einvp_4
XANTENNA_input613_A mprj_dat_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[91\]_TE mprj_logic_high_inst/HI[293] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[1\]_A user_to_mprj_in_gates\[1\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output665_A output665/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_54 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[42\]_A input68/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output832_A output832/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput90 la_data_out_core[62] vssd vssd vccd vccd input90/X sky130_fd_sc_hd__buf_4
XANTENNA_user_to_mprj_in_gates\[33\]_A input58/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_516 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output1027_A output1027/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_550_ _550_/A vssd vssd vccd vccd _550_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[26\] _618_/Y mprj_logic_high_inst/HI[228] vssd vssd vccd
+ vccd output929/A sky130_fd_sc_hd__einvp_4
Xuser_to_mprj_oen_buffers\[8\] _600_/Y mprj_logic_high_inst/HI[210] vssd vssd vccd
+ vccd output999/A sky130_fd_sc_hd__einvp_2
Xla_buf_enable\[48\] _640_/A la_buf_enable\[48\]/B vssd vssd vccd vccd la_buf\[48\]/TE
+ sky130_fd_sc_hd__and2b_1
X_481_ _481_/A vssd vssd vccd vccd _481_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input396_A la_oenb_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input563_A mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[1\] _465_/Y la_buf\[1\]/TE vssd vssd vccd vccd output666/A sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[24\]_A input48/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput461 la_oenb_mprj[50] vssd vssd vccd vccd _642_/A sky130_fd_sc_hd__clkbuf_2
Xinput450 la_oenb_mprj[40] vssd vssd vccd vccd _632_/A sky130_fd_sc_hd__buf_4
Xinput472 la_oenb_mprj[60] vssd vssd vccd vccd _652_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput483 la_oenb_mprj[70] vssd vssd vccd vccd _333_/A sky130_fd_sc_hd__buf_2
Xinput494 la_oenb_mprj[80] vssd vssd vccd vccd _343_/A sky130_fd_sc_hd__buf_4
XFILLER_35_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output782_A output782/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput902 output902/A vssd vssd vccd vccd la_oenb_core[117] sky130_fd_sc_hd__buf_2
Xoutput913 output913/A vssd vssd vccd vccd la_oenb_core[127] sky130_fd_sc_hd__buf_2
Xoutput924 output924/A vssd vssd vccd vccd la_oenb_core[21] sky130_fd_sc_hd__buf_2
Xoutput946 output946/A vssd vssd vccd vccd la_oenb_core[41] sky130_fd_sc_hd__buf_2
Xoutput935 output935/A vssd vssd vccd vccd la_oenb_core[31] sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_gates\[15\]_A input38/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput979 output979/A vssd vssd vccd vccd la_oenb_core[71] sky130_fd_sc_hd__buf_2
Xoutput968 output968/A vssd vssd vccd vccd la_oenb_core[61] sky130_fd_sc_hd__buf_2
Xoutput957 output957/A vssd vssd vccd vccd la_oenb_core[51] sky130_fd_sc_hd__buf_2
XFILLER_45_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input144_A la_data_out_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_602_ _602_/A vssd vssd vccd vccd _602_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input311_A la_iena_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input409_A la_oenb_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_533_ _533_/A vssd vssd vccd vccd _533_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_464_ _464_/A vssd vssd vccd vccd _464_/Y sky130_fd_sc_hd__clkinv_2
Xla_buf\[53\] _517_/Y la_buf\[53\]/TE vssd vssd vccd vccd output703/A sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[125\] input288/X mprj_logic_high_inst/HI[455] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[125\]/B sky130_fd_sc_hd__and2_1
XFILLER_13_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_395_ _395_/A vssd vssd vccd vccd _395_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_13_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[17\] _417_/Y mprj_adr_buf\[17\]/TE vssd vssd vccd vccd output1020/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output628_A output628/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[97\] user_to_mprj_in_gates\[97\]/Y vssd vssd vccd vccd output879/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_7_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput280 la_iena_mprj[118] vssd vssd vccd vccd input280/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_oen_buffers\[103\]_TE mprj_logic_high_inst/HI[305] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput291 la_iena_mprj[12] vssd vssd vccd vccd input291/X sky130_fd_sc_hd__buf_2
XFILLER_3_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output997_A output997/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[42\] input68/X user_to_mprj_in_gates\[42\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[42\]/Y sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_buffers\[7\] user_wb_dat_gates\[7\]/Y vssd vssd vccd vccd output1074/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_24_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[121\]_A input284/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput721 output721/A vssd vssd vccd vccd la_data_in_core[6] sky130_fd_sc_hd__buf_2
Xoutput710 output710/A vssd vssd vccd vccd la_data_in_core[5] sky130_fd_sc_hd__buf_2
XFILLER_12_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput754 output754/A vssd vssd vccd vccd la_data_in_core[9] sky130_fd_sc_hd__buf_2
Xoutput732 output732/A vssd vssd vccd vccd la_data_in_core[7] sky130_fd_sc_hd__buf_2
Xoutput743 output743/A vssd vssd vccd vccd la_data_in_core[8] sky130_fd_sc_hd__buf_2
XFILLER_28_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[4\] input76/X user_to_mprj_in_gates\[4\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[4\]/Y sky130_fd_sc_hd__nand2_2
Xoutput787 output787/A vssd vssd vccd vccd la_data_in_mprj[13] sky130_fd_sc_hd__buf_2
XFILLER_8_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput765 output765/A vssd vssd vccd vccd la_data_in_mprj[109] sky130_fd_sc_hd__buf_2
Xoutput776 output776/A vssd vssd vccd vccd la_data_in_mprj[119] sky130_fd_sc_hd__buf_2
XFILLER_28_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput798 output798/A vssd vssd vccd vccd la_data_in_mprj[23] sky130_fd_sc_hd__buf_2
XTAP_250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output1094_A output1094/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[112\]_A input274/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_2152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[93\] _356_/Y mprj_logic_high_inst/HI[295] vssd vssd vccd
+ vccd output1003/A sky130_fd_sc_hd__einvp_4
XFILLER_2_633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input261_A la_iena_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input359_A la_iena_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[126\]_TE mprj_logic_high_inst/HI[328] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[6\] input354/X mprj_logic_high_inst/HI[336] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[6\]/B sky130_fd_sc_hd__and2_1
XANTENNA_input526_A mprj_adr_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[116\] _379_/A la_buf_enable\[116\]/B vssd vssd vccd vccd la_buf\[116\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_18_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_516_ _516_/A vssd vssd vccd vccd _516_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[103\]_A input264/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_447_ _447_/A vssd vssd vccd vccd _447_/Y sky130_fd_sc_hd__inv_4
XFILLER_20_209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_378_ _378_/A vssd vssd vccd vccd _378_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[12\] user_to_mprj_in_gates\[12\]/Y vssd vssd vccd vccd output786/A
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_output745_A output745/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[40\]_TE la_buf\[40\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output912_A output912/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[25\]_TE mprj_logic_high_inst/HI[227] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[108\]_A_N _371_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1107_A output1107/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[52\] input335/X mprj_logic_high_inst/HI[382] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[52\]/B sky130_fd_sc_hd__and2_1
XFILLER_46_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[92\]_A input379/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input107_A la_data_out_core[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[30\] _622_/A la_buf_enable\[30\]/B vssd vssd vccd vccd la_buf\[30\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_24_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[4\] user_to_mprj_in_gates\[4\]/Y vssd vssd vccd vccd output827/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_32_1800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input476_A la_oenb_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input72_A la_data_out_core[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[63\]_TE la_buf\[63\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[16\] _480_/Y la_buf\[16\]/TE vssd vssd vccd vccd output662/A sky130_fd_sc_hd__einvp_8
XFILLER_48_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[48\]_TE mprj_logic_high_inst/HI[250] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__599__A _599_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[9\] _409_/Y mprj_adr_buf\[9\]/TE vssd vssd vccd vccd output1043/A sky130_fd_sc_hd__einvp_8
XFILLER_43_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_89 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[83\]_A input369/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output695_A output695/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output862_A output862/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[18\] input559/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[18\]/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_50_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_buffers\[15\] user_wb_dat_gates\[15\]/Y vssd vssd vccd vccd output1051/A
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_mprj_dat_buf\[12\]_TE mprj_dat_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[116\] input22/X user_to_mprj_in_gates\[116\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[116\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[74\]_A input359/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[86\]_TE la_buf\[86\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1057_A output1057/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[6\]_A_N _598_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[126\] _389_/Y mprj_logic_high_inst/HI[328] vssd vssd vccd
+ vccd output912/A sky130_fd_sc_hd__einvp_2
XFILLER_48_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[78\] _341_/A la_buf_enable\[78\]/B vssd vssd vccd vccd la_buf\[78\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[56\] _648_/Y mprj_logic_high_inst/HI[258] vssd vssd vccd
+ vccd output962/A sky130_fd_sc_hd__einvp_8
XFILLER_48_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input224_A la_data_out_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[65\]_A input349/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input593_A mprj_dat_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_61 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[113\] user_to_mprj_in_gates\[113\]/Y vssd vssd vccd vccd
+ output770/A sky130_fd_sc_hd__clkinv_4
XFILLER_39_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output708_A output708/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[56\]_A input339/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[60\]_B user_to_mprj_in_gates\[60\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xoutput1031 output1031/A vssd vssd vccd vccd mprj_adr_o_user[27] sky130_fd_sc_hd__buf_2
Xoutput1042 output1042/A vssd vssd vccd vccd mprj_adr_o_user[8] sky130_fd_sc_hd__buf_2
Xoutput1020 output1020/A vssd vssd vccd vccd mprj_adr_o_user[17] sky130_fd_sc_hd__buf_2
XFILLER_44_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput109 la_data_out_core[7] vssd vssd vccd vccd input109/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_1670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput1075 output1075/A vssd vssd vccd vccd mprj_dat_i_core[8] sky130_fd_sc_hd__buf_2
Xoutput1053 output1053/A vssd vssd vccd vccd mprj_dat_i_core[17] sky130_fd_sc_hd__buf_2
Xoutput1064 output1064/A vssd vssd vccd vccd mprj_dat_i_core[27] sky130_fd_sc_hd__buf_2
Xoutput1097 output1097/A vssd vssd vccd vccd mprj_dat_o_user[28] sky130_fd_sc_hd__buf_2
Xoutput1086 output1086/A vssd vssd vccd vccd mprj_dat_o_user[18] sky130_fd_sc_hd__buf_2
XFILLER_5_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[47\]_A input329/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[15\] input294/X mprj_logic_high_inst/HI[345] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[15\]/B sky130_fd_sc_hd__and2_1
XFILLER_16_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input174_A la_data_out_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[51\]_B user_to_mprj_in_gates\[51\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input341_A la_iena_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput621 user_irq_core[0] vssd vssd vccd vccd input621/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input439_A la_oenb_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput610 mprj_dat_o_core[6] vssd vssd vccd vccd _438_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_input35_A la_data_out_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[83\] _547_/Y la_buf\[83\]/TE vssd vssd vccd vccd output736/A sky130_fd_sc_hd__einvp_4
XANTENNA_user_to_mprj_in_ena_buf\[38\]_A input319/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input606_A mprj_dat_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[5\]_A _437_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output658_A output658/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_88 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[51\]_A_N _643_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[42\]_B user_to_mprj_in_gates\[42\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output825_A output825/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[72\] input101/X user_to_mprj_in_gates\[72\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[72\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[66\]_A_N _329_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[29\]_A input309/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput91 la_data_out_core[63] vssd vssd vccd vccd input91/X sky130_fd_sc_hd__buf_4
Xinput80 la_data_out_core[53] vssd vssd vccd vccd input80/X sky130_fd_sc_hd__buf_4
XANTENNA_la_buf_enable\[19\]_A_N _611_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[94\]_A user_to_mprj_in_gates\[94\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[33\]_B user_to_mprj_in_gates\[33\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[111\]_TE la_buf\[111\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[26\]_TE mprj_adr_buf\[26\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_480_ _480_/A vssd vssd vccd vccd _480_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[19\] _611_/Y mprj_logic_high_inst/HI[221] vssd vssd vccd
+ vccd output921/A sky130_fd_sc_hd__einvp_2
XFILLER_38_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input291_A la_iena_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input389_A la_oenb_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[121\]_A _585_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input556_A mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[24\]_B user_to_mprj_in_gates\[24\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[85\]_A user_to_mprj_in_gates\[85\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__400__A _400_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput462 la_oenb_mprj[51] vssd vssd vccd vccd _643_/A sky130_fd_sc_hd__clkbuf_2
Xinput451 la_oenb_mprj[41] vssd vssd vccd vccd _633_/A sky130_fd_sc_hd__clkbuf_2
Xinput440 la_oenb_mprj[31] vssd vssd vccd vccd _623_/A sky130_fd_sc_hd__buf_2
Xinput473 la_oenb_mprj[61] vssd vssd vccd vccd _653_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput484 la_oenb_mprj[71] vssd vssd vccd vccd _334_/A sky130_fd_sc_hd__clkbuf_2
Xinput495 la_oenb_mprj[81] vssd vssd vccd vccd _344_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[42\] user_to_mprj_in_gates\[42\]/Y vssd vssd vccd vccd output819/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_16_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output775_A output775/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[123\]_A user_to_mprj_in_gates\[123\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output942_A output942/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput903 output903/A vssd vssd vccd vccd la_oenb_core[118] sky130_fd_sc_hd__buf_2
XANTENNA_la_buf\[112\]_A _576_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput936 output936/A vssd vssd vccd vccd la_oenb_core[32] sky130_fd_sc_hd__buf_2
Xoutput925 output925/A vssd vssd vccd vccd la_oenb_core[22] sky130_fd_sc_hd__buf_2
Xoutput914 output914/A vssd vssd vccd vccd la_oenb_core[12] sky130_fd_sc_hd__buf_2
XFILLER_47_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[15\]_B user_to_mprj_in_gates\[15\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[76\]_A user_to_mprj_in_gates\[76\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xoutput969 output969/A vssd vssd vccd vccd la_oenb_core[62] sky130_fd_sc_hd__buf_2
Xoutput958 output958/A vssd vssd vccd vccd la_oenb_core[52] sky130_fd_sc_hd__buf_2
Xoutput947 output947/A vssd vssd vccd vccd la_oenb_core[42] sky130_fd_sc_hd__buf_2
XTAP_410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[114\]_A user_to_mprj_in_gates\[114\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[103\]_A _567_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[67\]_A user_to_mprj_in_gates\[67\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[40\]_A _504_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[82\] input368/X mprj_logic_high_inst/HI[412] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[82\]/B sky130_fd_sc_hd__and2_1
XFILLER_11_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[81\]_TE mprj_logic_high_inst/HI[283] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[60\] _652_/A la_buf_enable\[60\]/B vssd vssd vccd vccd la_buf\[60\]/TE
+ sky130_fd_sc_hd__and2b_1
X_601_ _601_/A vssd vssd vccd vccd _601_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input137_A la_data_out_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_532_ _532_/A vssd vssd vccd vccd _532_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_27_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input304_A la_iena_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_463_ _463_/A vssd vssd vccd vccd _463_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_2_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[46\] _510_/Y la_buf\[46\]/TE vssd vssd vccd vccd output695/A sky130_fd_sc_hd__einvp_8
X_394_ _394_/A vssd vssd vccd vccd _394_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_51_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[118\] input280/X mprj_logic_high_inst/HI[448] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[118\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_buffers\[105\]_A user_to_mprj_in_gates\[105\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[58\]_A user_to_mprj_in_gates\[58\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[31\]_A _495_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[102\] _566_/Y la_buf\[102\]/TE vssd vssd vccd vccd output630/A sky130_fd_sc_hd__einvp_2
XFILLER_4_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_870 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput270 la_iena_mprj[109] vssd vssd vccd vccd input270/X sky130_fd_sc_hd__clkbuf_1
Xinput281 la_iena_mprj[119] vssd vssd vccd vccd input281/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput292 la_iena_mprj[13] vssd vssd vccd vccd input292/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output892_A output892/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[98\]_A _562_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[121\]_B mprj_logic_high_inst/HI[451] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[35\] input60/X user_to_mprj_in_gates\[35\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[35\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput711 output711/A vssd vssd vccd vccd la_data_in_core[60] sky130_fd_sc_hd__buf_2
Xoutput700 output700/A vssd vssd vccd vccd la_data_in_core[50] sky130_fd_sc_hd__buf_2
XFILLER_12_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[49\]_A user_to_mprj_in_gates\[49\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xoutput744 output744/A vssd vssd vccd vccd la_data_in_core[90] sky130_fd_sc_hd__buf_2
Xoutput733 output733/A vssd vssd vccd vccd la_data_in_core[80] sky130_fd_sc_hd__buf_2
Xoutput722 output722/A vssd vssd vccd vccd la_data_in_core[70] sky130_fd_sc_hd__buf_2
XFILLER_47_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[22\]_A _486_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput777 output777/A vssd vssd vccd vccd la_data_in_mprj[11] sky130_fd_sc_hd__buf_2
Xoutput766 output766/A vssd vssd vccd vccd la_data_in_mprj[10] sky130_fd_sc_hd__buf_2
Xoutput755 output755/A vssd vssd vccd vccd la_data_in_mprj[0] sky130_fd_sc_hd__buf_2
Xoutput788 output788/A vssd vssd vccd vccd la_data_in_mprj[14] sky130_fd_sc_hd__buf_2
XFILLER_48_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[40\]_B la_buf_enable\[40\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput799 output799/A vssd vssd vccd vccd la_data_in_mprj[24] sky130_fd_sc_hd__buf_2
XTAP_240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[89\]_A _553_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[112\]_B mprj_logic_high_inst/HI[442] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output1087_A output1087/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[86\] _349_/Y mprj_logic_high_inst/HI[288] vssd vssd vccd
+ vccd output995/A sky130_fd_sc_hd__einvp_2
XANTENNA_la_buf\[13\]_A _477_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input254_A la_data_out_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[31\]_B la_buf_enable\[31\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[0\]_A input260/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input421_A la_oenb_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input519_A mprj_adr_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[109\] _372_/A la_buf_enable\[109\]/B vssd vssd vccd vccd la_buf\[109\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_18_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_515_ _515_/A vssd vssd vccd vccd _515_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[103\]_B mprj_logic_high_inst/HI[433] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_1951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_446_ _446_/A vssd vssd vccd vccd _446_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf_enable\[98\]_B la_buf_enable\[98\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_377_ _377_/A vssd vssd vccd vccd _377_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output640_A output640/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output738_A output738/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[22\]_B la_buf_enable\[22\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output905_A output905/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[89\]_B la_buf_enable\[89\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[91\]_A _354_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[13\]_B la_buf_enable\[13\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output1002_A output1002/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[45\] input327/X mprj_logic_high_inst/HI[375] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[45\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_ena_buf\[92\]_B mprj_logic_high_inst/HI[422] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_1214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[23\] _615_/A la_buf_enable\[23\]/B vssd vssd vccd vccd la_buf\[23\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_24_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[82\]_A _345_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input469_A la_oenb_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input371_A la_iena_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input65_A la_data_out_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[83\]_B mprj_logic_high_inst/HI[413] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_34_836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1712 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output688_A output688/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_429_ _429_/A vssd vssd vccd vccd _429_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_31_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[73\]_A _336_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output855_A output855/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[0\]_A input550/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput1 caravel_clk vssd vssd vccd vccd _391_/A sky130_fd_sc_hd__clkbuf_1
Xuser_to_mprj_in_gates\[109\] input14/X user_to_mprj_in_gates\[109\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[109\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[74\]_B mprj_logic_high_inst/HI[404] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_52_633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[0\]_A input4/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[116\]_TE mprj_logic_high_inst/HI[318] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[64\]_A _656_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[119\] _382_/Y mprj_logic_high_inst/HI[321] vssd vssd vccd
+ vccd output904/A sky130_fd_sc_hd__einvp_4
XFILLER_0_946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[49\] _641_/Y mprj_logic_high_inst/HI[251] vssd vssd vccd
+ vccd output954/A sky130_fd_sc_hd__einvp_2
XFILLER_47_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[65\]_B mprj_logic_high_inst/HI[395] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input217_A la_data_out_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[30\]_TE la_buf\[30\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[15\]_TE mprj_logic_high_inst/HI[217] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input586_A mprj_dat_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[55\]_A _647_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[100\] input261/X mprj_logic_high_inst/HI[430] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[100\]/B sky130_fd_sc_hd__and2_1
Xuser_wb_dat_gates\[0\] input550/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[0\]/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_7_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__403__A _403_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[107\]_A_N _370_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[106\] user_to_mprj_in_gates\[106\]/Y vssd vssd vccd vccd
+ output762/A sky130_fd_sc_hd__inv_2
XFILLER_43_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[56\]_B mprj_logic_high_inst/HI[386] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[72\] user_to_mprj_in_gates\[72\]/Y vssd vssd vccd vccd output852/A
+ sky130_fd_sc_hd__inv_2
XFILLER_4_1275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output972_A output972/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[30\] input573/X repeater1125/X vssd vssd vccd vccd user_wb_dat_gates\[30\]/Y
+ sky130_fd_sc_hd__nand2_8
XFILLER_33_2118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[46\]_A _638_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput1010 output1010/A vssd vssd vccd vccd la_oenb_core[9] sky130_fd_sc_hd__buf_2
Xoutput1032 output1032/A vssd vssd vccd vccd mprj_adr_o_user[28] sky130_fd_sc_hd__buf_2
Xoutput1021 output1021/A vssd vssd vccd vccd mprj_adr_o_user[18] sky130_fd_sc_hd__buf_2
XFILLER_44_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput1043 output1043/A vssd vssd vccd vccd mprj_adr_o_user[9] sky130_fd_sc_hd__buf_2
XFILLER_48_1682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[5\] _437_/Y mprj_dat_buf\[5\]/TE vssd vssd vccd vccd output1104/A sky130_fd_sc_hd__einvp_8
Xoutput1076 output1076/A vssd vssd vccd vccd mprj_dat_i_core[9] sky130_fd_sc_hd__buf_2
Xoutput1054 output1054/A vssd vssd vccd vccd mprj_dat_i_core[18] sky130_fd_sc_hd__buf_2
Xoutput1065 output1065/A vssd vssd vccd vccd mprj_dat_i_core[28] sky130_fd_sc_hd__buf_2
Xoutput1098 output1098/A vssd vssd vccd vccd mprj_dat_o_user[29] sky130_fd_sc_hd__buf_2
Xoutput1087 output1087/A vssd vssd vccd vccd mprj_dat_o_user[19] sky130_fd_sc_hd__buf_2
XFILLER_44_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[47\]_B mprj_logic_high_inst/HI[377] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[53\]_TE la_buf\[53\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[38\]_TE mprj_logic_high_inst/HI[240] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[37\]_A _629_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input167_A la_data_out_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[90\] _353_/A la_buf_enable\[90\]/B vssd vssd vccd vccd la_buf\[90\]/TE
+ sky130_fd_sc_hd__and2b_1
Xinput622 user_irq_core[1] vssd vssd vccd vccd input622/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput611 mprj_dat_o_core[7] vssd vssd vccd vccd _439_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput600 mprj_dat_o_core[26] vssd vssd vccd vccd _458_/A sky130_fd_sc_hd__buf_2
XFILLER_43_1045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input334_A la_iena_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input28_A la_data_out_core[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[38\]_B mprj_logic_high_inst/HI[368] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_47_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input501_A la_oenb_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[76\] _540_/Y la_buf\[76\]/TE vssd vssd vccd vccd output728/A sky130_fd_sc_hd__einvp_4
XFILLER_1_1448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[28\]_A _620_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output720_A output720/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output818_A output818/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[76\]_TE la_buf\[76\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[24\]_A _424_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[29\]_B mprj_logic_high_inst/HI[359] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[65\] input93/X user_to_mprj_in_gates\[65\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[65\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[5\]_A_N _597_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[19\]_A _611_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[1\]_A _593_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput81 la_data_out_core[54] vssd vssd vccd vccd input81/X sky130_fd_sc_hd__clkbuf_4
Xinput70 la_data_out_core[44] vssd vssd vccd vccd input70/X sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput92 la_data_out_core[64] vssd vssd vccd vccd input92/X sky130_fd_sc_hd__buf_4
XFILLER_44_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[15\]_A _415_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[25\]_TE mprj_dat_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2026 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[4\]_TE mprj_logic_high_inst/HI[206] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input284_A la_iena_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input451_A la_oenb_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input549_A mprj_cyc_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[99\]_TE la_buf\[99\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput430 la_oenb_mprj[22] vssd vssd vccd vccd _614_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput463 la_oenb_mprj[52] vssd vssd vccd vccd _644_/A sky130_fd_sc_hd__clkbuf_2
Xinput452 la_oenb_mprj[42] vssd vssd vccd vccd _634_/A sky130_fd_sc_hd__buf_4
Xinput441 la_oenb_mprj[32] vssd vssd vccd vccd _624_/A sky130_fd_sc_hd__buf_2
XFILLER_5_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput474 la_oenb_mprj[62] vssd vssd vccd vccd _654_/A sky130_fd_sc_hd__clkbuf_2
Xinput485 la_oenb_mprj[72] vssd vssd vccd vccd _335_/A sky130_fd_sc_hd__buf_2
Xinput496 la_oenb_mprj[82] vssd vssd vccd vccd _345_/A sky130_fd_sc_hd__buf_4
XFILLER_40_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[35\] user_to_mprj_in_gates\[35\]/Y vssd vssd vccd vccd output811/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output670_A output670/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output768_A output768/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output935_A output935/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput904 output904/A vssd vssd vccd vccd la_oenb_core[119] sky130_fd_sc_hd__buf_2
Xoutput926 output926/A vssd vssd vccd vccd la_oenb_core[23] sky130_fd_sc_hd__buf_2
Xoutput937 output937/A vssd vssd vccd vccd la_oenb_core[33] sky130_fd_sc_hd__buf_2
Xoutput915 output915/A vssd vssd vccd vccd la_oenb_core[13] sky130_fd_sc_hd__buf_2
XFILLER_28_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput959 output959/A vssd vssd vccd vccd la_oenb_core[53] sky130_fd_sc_hd__buf_2
Xoutput948 output948/A vssd vssd vccd vccd la_oenb_core[43] sky130_fd_sc_hd__buf_2
XFILLER_45_2320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_19 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2346 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1032_A output1032/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__501__A _501_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[75\] input360/X mprj_logic_high_inst/HI[405] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[75\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[101\] _364_/Y mprj_logic_high_inst/HI[303] vssd vssd vccd
+ vccd output885/A sky130_fd_sc_hd__einvp_2
XFILLER_24_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_600_ _600_/A vssd vssd vccd vccd _600_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_2244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[31\] _623_/Y mprj_logic_high_inst/HI[233] vssd vssd vccd
+ vccd output935/A sky130_fd_sc_hd__einvp_2
X_531_ _531_/A vssd vssd vccd vccd _531_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[53\] _645_/A la_buf_enable\[53\]/B vssd vssd vccd vccd la_buf\[53\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_27_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_462_ _462_/A vssd vssd vccd vccd _462_/Y sky130_fd_sc_hd__inv_4
XANTENNA_la_buf_enable\[50\]_A_N _642_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_393_ _393_/A vssd vssd vccd vccd _393_/Y sky130_fd_sc_hd__inv_6
XFILLER_13_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input499_A la_oenb_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input95_A la_data_out_core[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[65\]_A_N _657_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[39\] _503_/Y la_buf\[39\]/TE vssd vssd vccd vccd output687/A sky130_fd_sc_hd__einvp_8
XFILLER_51_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__411__A _411_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[28\]_A _460_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput260 la_iena_mprj[0] vssd vssd vccd vccd input260/X sky130_fd_sc_hd__clkbuf_1
Xinput271 la_iena_mprj[10] vssd vssd vccd vccd input271/X sky130_fd_sc_hd__buf_2
XFILLER_49_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput282 la_iena_mprj[11] vssd vssd vccd vccd input282/X sky130_fd_sc_hd__clkbuf_2
Xinput293 la_iena_mprj[14] vssd vssd vccd vccd input293/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[18\]_A_N _610_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output885_A output885/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[28\] input52/X user_to_mprj_in_gates\[28\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[28\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_34_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[101\]_TE la_buf\[101\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[0\]_A _400_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[16\]_TE mprj_adr_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput712 output712/A vssd vssd vccd vccd la_data_in_core[61] sky130_fd_sc_hd__buf_2
Xoutput701 output701/A vssd vssd vccd vccd la_data_in_core[51] sky130_fd_sc_hd__buf_2
Xoutput734 output734/A vssd vssd vccd vccd la_data_in_core[81] sky130_fd_sc_hd__buf_2
Xoutput723 output723/A vssd vssd vccd vccd la_data_in_core[71] sky130_fd_sc_hd__buf_2
Xoutput745 output745/A vssd vssd vccd vccd la_data_in_core[91] sky130_fd_sc_hd__buf_2
Xoutput756 output756/A vssd vssd vccd vccd la_data_in_mprj[100] sky130_fd_sc_hd__buf_2
Xoutput767 output767/A vssd vssd vccd vccd la_data_in_mprj[110] sky130_fd_sc_hd__buf_2
Xoutput778 output778/A vssd vssd vccd vccd la_data_in_mprj[120] sky130_fd_sc_hd__buf_2
XFILLER_45_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[0\]_TE mprj_adr_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput789 output789/A vssd vssd vccd vccd la_data_in_mprj[15] sky130_fd_sc_hd__buf_2
XTAP_230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[19\]_A _451_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_buffers\[26\]_A user_wb_dat_gates\[26\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_45_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[79\] _342_/Y mprj_logic_high_inst/HI[281] vssd vssd vccd
+ vccd output987/A sky130_fd_sc_hd__einvp_2
XFILLER_1_101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[27\] _459_/Y mprj_dat_buf\[27\]/TE vssd vssd vccd vccd output1096/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_2223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[4\]_TE mprj_dat_buf\[4\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input247_A la_data_out_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[0\]_B mprj_logic_high_inst/HI[330] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_buffers\[17\]_A user_wb_dat_gates\[17\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input414_A la_oenb_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input10_A la_data_out_core[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_514_ _514_/A vssd vssd vccd vccd _514_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[124\]_TE la_buf\[124\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_445_ _445_/A vssd vssd vccd vccd _445_/Y sky130_fd_sc_hd__inv_2
XTAP_1996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_376_ _376_/A vssd vssd vccd vccd _376_/Y sky130_fd_sc_hd__inv_2
XANTENNA__406__A _406_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[22\] _422_/Y mprj_adr_buf\[22\]/TE vssd vssd vccd vccd output1026/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output633_A output633/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1516 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output800_A output800/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[121\]_B la_buf_enable\[121\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[71\]_TE mprj_logic_high_inst/HI[273] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[7\] _599_/A la_buf_enable\[7\]/B vssd vssd vccd vccd la_buf\[7\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_gates\[90\]_A input121/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input2_A caravel_clk2 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[112\]_B la_buf_enable\[112\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[38\] input319/X mprj_logic_high_inst/HI[368] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[38\]/B sky130_fd_sc_hd__and2_1
XTAP_1215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[16\] _608_/A la_buf_enable\[16\]/B vssd vssd vccd vccd la_buf\[16\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_11_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input197_A la_data_out_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[3\]_A user_wb_dat_gates\[3\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[81\]_A input111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input364_A la_iena_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input58_A la_data_out_core[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input531_A mprj_adr_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[121\] _384_/A la_buf_enable\[121\]/B vssd vssd vccd vccd la_buf\[121\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_24_2053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_47 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[6\]_A _470_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[103\]_B la_buf_enable\[103\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[94\]_TE mprj_logic_high_inst/HI[296] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_428_ _428_/A vssd vssd vccd vccd _428_/Y sky130_fd_sc_hd__inv_8
XFILLER_14_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_359_ _359_/A vssd vssd vccd vccd _359_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output750_A output750/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output848_A output848/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[72\]_A input101/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[95\] input126/X user_to_mprj_in_gates\[95\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[95\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[0\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput2 caravel_clk2 vssd vssd vccd vccd _392_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[0\]_B user_to_mprj_in_gates\[0\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_51_188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1234 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[63\]_A input91/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1112_A output1112/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input112_A la_data_out_core[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_75 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input579_A mprj_dat_i_user[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_52 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input481_A la_oenb_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[21\] _485_/Y la_buf\[21\]/TE vssd vssd vccd vccd output668/A sky130_fd_sc_hd__einvp_8
XFILLER_7_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[54\]_A input81/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[4\]_A user_to_mprj_in_gates\[4\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[65\] user_to_mprj_in_gates\[65\]/Y vssd vssd vccd vccd output844/A
+ sky130_fd_sc_hd__inv_2
XFILLER_37_2233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output798_A output798/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output965_A output965/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[23\] input565/X repeater1125/X vssd vssd vccd vccd user_wb_dat_gates\[23\]/Y
+ sky130_fd_sc_hd__nand2_8
XTAP_1590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[10\] input15/X user_to_mprj_in_gates\[10\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[10\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_14_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[45\]_A input71/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput1000 output1000/A vssd vssd vccd vccd la_oenb_core[90] sky130_fd_sc_hd__buf_2
Xuser_wb_dat_buffers\[20\] user_wb_dat_gates\[20\]/Y vssd vssd vccd vccd output1057/A
+ sky130_fd_sc_hd__clkinv_8
Xoutput1033 output1033/A vssd vssd vccd vccd mprj_adr_o_user[29] sky130_fd_sc_hd__buf_2
Xoutput1022 output1022/A vssd vssd vccd vccd mprj_adr_o_user[19] sky130_fd_sc_hd__buf_2
Xoutput1011 output1011/A vssd vssd vccd vccd mprj_ack_i_core sky130_fd_sc_hd__buf_2
Xoutput1044 output1044/A vssd vssd vccd vccd mprj_cyc_o_user sky130_fd_sc_hd__buf_2
XFILLER_44_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput1055 output1055/A vssd vssd vccd vccd mprj_dat_i_core[19] sky130_fd_sc_hd__buf_2
Xoutput1066 output1066/A vssd vssd vccd vccd mprj_dat_i_core[29] sky130_fd_sc_hd__buf_2
Xoutput1088 output1088/A vssd vssd vccd vccd mprj_dat_o_user[1] sky130_fd_sc_hd__buf_2
Xoutput1077 output1077/A vssd vssd vccd vccd mprj_dat_o_user[0] sky130_fd_sc_hd__buf_2
Xoutput1099 output1099/A vssd vssd vccd vccd mprj_dat_o_user[2] sky130_fd_sc_hd__buf_2
XFILLER_48_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[121\] input28/X user_to_mprj_in_gates\[121\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[121\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output1062_A output1062/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__504__A _504_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[120\]_A input27/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[36\]_A input61/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[61\] _653_/Y mprj_logic_high_inst/HI[263] vssd vssd vccd
+ vccd output968/A sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[83\] _346_/A la_buf_enable\[83\]/B vssd vssd vccd vccd la_buf\[83\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_27_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput612 mprj_dat_o_core[8] vssd vssd vccd vccd _440_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput601 mprj_dat_o_core[27] vssd vssd vccd vccd _459_/A sky130_fd_sc_hd__clkbuf_2
Xinput623 user_irq_core[2] vssd vssd vccd vccd input623/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input327_A la_iena_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1438 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[69\] _533_/Y la_buf\[69\]/TE vssd vssd vccd vccd output720/A sky130_fd_sc_hd__einvp_8
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[27\]_A input51/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__414__A _414_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[111\]_A input17/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[125\] _589_/Y la_buf\[125\]/TE vssd vssd vccd vccd output655/A sky130_fd_sc_hd__einvp_2
XFILLER_10_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output713_A output713/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[106\]_TE mprj_logic_high_inst/HI[308] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[58\] input85/X user_to_mprj_in_gates\[58\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[58\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[18\]_A input41/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_A input7/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput82 la_data_out_core[55] vssd vssd vccd vccd input82/X sky130_fd_sc_hd__buf_4
Xinput71 la_data_out_core[45] vssd vssd vccd vccd input71/X sky130_fd_sc_hd__buf_4
Xinput60 la_data_out_core[35] vssd vssd vccd vccd input60/X sky130_fd_sc_hd__clkbuf_4
Xinput93 la_data_out_core[65] vssd vssd vccd vccd input93/X sky130_fd_sc_hd__buf_4
XFILLER_11_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[20\]_TE la_buf\[20\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[20\] input300/X mprj_logic_high_inst/HI[350] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[20\]/B sky130_fd_sc_hd__and2_1
XFILLER_40_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[106\]_A_N _369_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_54 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input277_A la_iena_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input40_A la_data_out_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input444_A la_oenb_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput420 la_oenb_mprj[13] vssd vssd vccd vccd _605_/A sky130_fd_sc_hd__buf_2
XFILLER_7_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput464 la_oenb_mprj[53] vssd vssd vccd vccd _645_/A sky130_fd_sc_hd__buf_2
Xinput453 la_oenb_mprj[43] vssd vssd vccd vccd _635_/A sky130_fd_sc_hd__buf_4
Xinput431 la_oenb_mprj[23] vssd vssd vccd vccd _615_/A sky130_fd_sc_hd__buf_2
Xinput442 la_oenb_mprj[33] vssd vssd vccd vccd _625_/A sky130_fd_sc_hd__buf_2
XANTENNA_input611_A mprj_dat_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput475 la_oenb_mprj[63] vssd vssd vccd vccd _655_/A sky130_fd_sc_hd__buf_2
Xinput486 la_oenb_mprj[73] vssd vssd vccd vccd _336_/A sky130_fd_sc_hd__buf_2
Xinput497 la_oenb_mprj[83] vssd vssd vccd vccd _346_/A sky130_fd_sc_hd__buf_4
XFILLER_48_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__409__A _409_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[28\] user_to_mprj_in_gates\[28\]/Y vssd vssd vccd vccd output803/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output663_A output663/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput927 output927/A vssd vssd vccd vccd la_oenb_core[24] sky130_fd_sc_hd__buf_2
Xoutput905 output905/A vssd vssd vccd vccd la_oenb_core[11] sky130_fd_sc_hd__buf_2
Xoutput916 output916/A vssd vssd vccd vccd la_oenb_core[14] sky130_fd_sc_hd__buf_2
XANTENNA_la_buf\[43\]_TE la_buf\[43\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output830_A output830/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput949 output949/A vssd vssd vccd vccd la_oenb_core[44] sky130_fd_sc_hd__buf_2
Xoutput938 output938/A vssd vssd vccd vccd la_oenb_core[34] sky130_fd_sc_hd__buf_2
XANTENNA_output928_A output928/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[28\]_TE mprj_logic_high_inst/HI[230] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[0\]_B la_buf_enable\[0\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[124\]_A input287/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output1025_A output1025/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[68\] input352/X mprj_logic_high_inst/HI[398] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[68\]/B sky130_fd_sc_hd__and2_1
XFILLER_40_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_530_ _530_/A vssd vssd vccd vccd _530_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[115\]_A input277/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_65 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[24\] _616_/Y mprj_logic_high_inst/HI[226] vssd vssd vccd
+ vccd output927/A sky130_fd_sc_hd__einvp_2
Xla_buf_enable\[46\] _638_/A la_buf_enable\[46\]/B vssd vssd vccd vccd la_buf\[46\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[6\] _598_/Y mprj_logic_high_inst/HI[208] vssd vssd vccd
+ vccd output977/A sky130_fd_sc_hd__einvp_2
X_461_ _461_/A vssd vssd vccd vccd _461_/Y sky130_fd_sc_hd__inv_4
XFILLER_32_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_392_ _392_/A vssd vssd vccd vccd _392_/Y sky130_fd_sc_hd__inv_4
XFILLER_41_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[66\]_TE la_buf\[66\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input394_A la_oenb_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input88_A la_data_out_core[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input561_A mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1590 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[4\]_A_N _596_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput250 la_data_out_mprj[91] vssd vssd vccd vccd _555_/A sky130_fd_sc_hd__clkbuf_1
Xinput261 la_iena_mprj[100] vssd vssd vccd vccd input261/X sky130_fd_sc_hd__clkbuf_1
Xinput272 la_iena_mprj[110] vssd vssd vccd vccd input272/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput294 la_iena_mprj[15] vssd vssd vccd vccd input294/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput283 la_iena_mprj[120] vssd vssd vccd vccd input283/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_in_ena_buf\[106\]_A input267/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output878_A output878/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output780_A output780/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput702 output702/A vssd vssd vccd vccd la_data_in_core[52] sky130_fd_sc_hd__buf_2
Xoutput735 output735/A vssd vssd vccd vccd la_data_in_core[82] sky130_fd_sc_hd__buf_2
Xoutput724 output724/A vssd vssd vccd vccd la_data_in_core[72] sky130_fd_sc_hd__buf_2
Xoutput713 output713/A vssd vssd vccd vccd la_data_in_core[62] sky130_fd_sc_hd__buf_2
XANTENNA_mprj_dat_buf\[15\]_TE mprj_dat_buf\[15\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__602__A _602_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput746 output746/A vssd vssd vccd vccd la_data_in_core[92] sky130_fd_sc_hd__buf_2
XFILLER_47_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput757 output757/A vssd vssd vccd vccd la_data_in_mprj[101] sky130_fd_sc_hd__buf_2
Xoutput768 output768/A vssd vssd vccd vccd la_data_in_mprj[111] sky130_fd_sc_hd__buf_2
Xoutput779 output779/A vssd vssd vccd vccd la_data_in_mprj[121] sky130_fd_sc_hd__buf_2
XFILLER_41_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[89\]_TE la_buf\[89\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__512__A _512_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[95\]_A input382/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input142_A la_data_out_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2020 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input407_A la_oenb_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_513_ _513_/A vssd vssd vccd vccd _513_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_444_ _444_/A vssd vssd vccd vccd _444_/Y sky130_fd_sc_hd__inv_4
XTAP_1975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[51\] _515_/Y la_buf\[51\]/TE vssd vssd vccd vccd output701/A sky130_fd_sc_hd__einvp_8
XTAP_1997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_375_ _375_/A vssd vssd vccd vccd _375_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[123\] input286/X mprj_logic_high_inst/HI[453] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[123\]/B sky130_fd_sc_hd__and2_1
XFILLER_13_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__422__A _422_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[15\] _415_/Y mprj_adr_buf\[15\]/TE vssd vssd vccd vccd output1018/A
+ sky130_fd_sc_hd__einvp_4
XFILLER_5_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[95\] user_to_mprj_in_gates\[95\]/Y vssd vssd vccd vccd output877/A
+ sky130_fd_sc_hd__inv_2
XFILLER_42_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[86\]_A input372/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output995_A output995/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[40\] input66/X user_to_mprj_in_gates\[40\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[40\]/Y sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_buffers\[5\] user_wb_dat_gates\[5\]/Y vssd vssd vccd vccd output1072/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_51_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[10\]_A input271/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[90\]_B user_to_mprj_in_gates\[90\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__332__A _332_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[2\] input54/X user_to_mprj_in_gates\[2\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[2\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_90 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[77\]_A input362/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[64\]_A_N _656_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output1092_A output1092/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[79\]_A_N _342_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__507__A _507_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[81\]_B user_to_mprj_in_gates\[81\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[91\] _354_/Y mprj_logic_high_inst/HI[293] vssd vssd vccd
+ vccd output1001/A sky130_fd_sc_hd__einvp_4
XANTENNA_la_buf_enable\[17\]_A_N _609_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input357_A la_iena_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[4\] input332/X mprj_logic_high_inst/HI[334] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[4\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_ena_buf\[68\]_A input352/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input524_A mprj_adr_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[99\] _563_/Y la_buf\[99\]/TE vssd vssd vccd vccd output753/A sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[114\] _377_/A la_buf_enable\[114\]/B vssd vssd vccd vccd la_buf\[114\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_1_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_427_ _427_/A vssd vssd vccd vccd _427_/Y sky130_fd_sc_hd__inv_8
XANTENNA__417__A _417_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_358_ _358_/A vssd vssd vccd vccd _358_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[10\] user_to_mprj_in_gates\[10\]/Y vssd vssd vccd vccd output766/A
+ sky130_fd_sc_hd__inv_6
XANTENNA_user_to_mprj_in_gates\[72\]_B user_to_mprj_in_gates\[72\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output743_A output743/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output910_A output910/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[88\] input118/X user_to_mprj_in_gates\[88\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[88\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[59\]_A input342/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput3 caravel_rstn vssd vssd vccd vccd input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[63\]_B user_to_mprj_in_gates\[63\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[114\]_TE la_buf\[114\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1105_A output1105/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[29\]_TE mprj_adr_buf\[29\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[50\] input333/X mprj_logic_high_inst/HI[380] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[50\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input105_A la_data_out_core[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_87 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[2\] user_to_mprj_in_gates\[2\]/Y vssd vssd vccd vccd output805/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_42_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input474_A la_oenb_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input70_A la_data_out_core[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[14\] _478_/Y la_buf\[14\]/TE vssd vssd vccd vccd output660/A sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[54\]_B user_to_mprj_in_gates\[54\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[61\]_TE mprj_logic_high_inst/HI[263] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[7\] _407_/Y mprj_adr_buf\[7\]/TE vssd vssd vccd vccd output1041/A sky130_fd_sc_hd__einvp_4
XFILLER_43_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[58\] user_to_mprj_in_gates\[58\]/Y vssd vssd vccd vccd output836/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output693_A output693/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[8\]_A _440_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output958_A output958/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output860_A output860/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[16\] input557/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[16\]/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_31_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[45\]_B user_to_mprj_in_gates\[45\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xoutput1001 output1001/A vssd vssd vccd vccd la_oenb_core[91] sky130_fd_sc_hd__buf_2
Xuser_wb_dat_buffers\[13\] user_wb_dat_gates\[13\]/Y vssd vssd vccd vccd output1049/A
+ sky130_fd_sc_hd__clkinv_8
Xoutput1023 output1023/A vssd vssd vccd vccd mprj_adr_o_user[1] sky130_fd_sc_hd__buf_2
Xoutput1012 output1012/A vssd vssd vccd vccd mprj_adr_o_user[0] sky130_fd_sc_hd__buf_2
XFILLER_44_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput1034 output1034/A vssd vssd vccd vccd mprj_adr_o_user[2] sky130_fd_sc_hd__buf_2
XFILLER_44_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput1045 output1045/A vssd vssd vccd vccd mprj_dat_i_core[0] sky130_fd_sc_hd__buf_2
Xoutput1067 output1067/A vssd vssd vccd vccd mprj_dat_i_core[2] sky130_fd_sc_hd__buf_2
Xoutput1056 output1056/A vssd vssd vccd vccd mprj_dat_i_core[1] sky130_fd_sc_hd__buf_2
Xoutput1089 output1089/A vssd vssd vccd vccd mprj_dat_o_user[20] sky130_fd_sc_hd__buf_2
Xoutput1078 output1078/A vssd vssd vccd vccd mprj_dat_o_user[10] sky130_fd_sc_hd__buf_2
XANTENNA__610__A _610_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[114\] input20/X user_to_mprj_in_gates\[114\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[114\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_1907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[30\]_A user_to_mprj_in_gates\[30\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[120\]_B user_to_mprj_in_gates\[120\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[36\]_B user_to_mprj_in_gates\[36\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[97\]_A user_to_mprj_in_gates\[97\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1055_A output1055/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[70\]_A _534_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[98\] input385/X mprj_logic_high_inst/HI[428] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[98\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[84\]_TE mprj_logic_high_inst/HI[286] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1150 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[124\] _387_/Y mprj_logic_high_inst/HI[326] vssd vssd vccd
+ vccd output910/A sky130_fd_sc_hd__einvp_2
XANTENNA__520__A _520_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput613 mprj_dat_o_core[9] vssd vssd vccd vccd _441_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput602 mprj_dat_o_core[28] vssd vssd vccd vccd _460_/A sky130_fd_sc_hd__clkbuf_2
Xinput624 user_irq_ena[0] vssd vssd vccd vccd input624/X sky130_fd_sc_hd__clkbuf_1
Xuser_to_mprj_oen_buffers\[54\] _646_/Y mprj_logic_high_inst/HI[256] vssd vssd vccd
+ vccd output960/A sky130_fd_sc_hd__einvp_4
XFILLER_48_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[76\] _339_/A la_buf_enable\[76\]/B vssd vssd vccd vccd la_buf\[76\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_5_2276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[21\]_A user_to_mprj_in_gates\[21\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_input222_A la_data_out_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input591_A mprj_dat_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[124\]_A _588_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[27\]_B user_to_mprj_in_gates\[27\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_69 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[88\]_A user_to_mprj_in_gates\[88\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[111\]_B user_to_mprj_in_gates\[111\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[61\]_A _525_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[118\] _582_/Y la_buf\[118\]/TE vssd vssd vccd vccd output647/A sky130_fd_sc_hd__einvp_2
XFILLER_10_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__430__A _430_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[111\] user_to_mprj_in_gates\[111\]/Y vssd vssd vccd vccd
+ output768/A sky130_fd_sc_hd__inv_2
XTAP_627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output706_A output706/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[12\]_A user_to_mprj_in_gates\[12\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_34_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[20\]_A input562/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[126\]_A user_to_mprj_in_gates\[126\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[115\]_A _579_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__605__A _605_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[18\]_B user_to_mprj_in_gates\[18\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[79\]_A user_to_mprj_in_gates\[79\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_B user_to_mprj_in_gates\[102\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xinput72 la_data_out_core[46] vssd vssd vccd vccd input72/X sky130_fd_sc_hd__buf_4
Xinput61 la_data_out_core[36] vssd vssd vccd vccd input61/X sky130_fd_sc_hd__clkbuf_4
Xinput50 la_data_out_core[26] vssd vssd vccd vccd input50/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_la_buf\[52\]_A _516_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput94 la_data_out_core[66] vssd vssd vccd vccd input94/X sky130_fd_sc_hd__buf_4
Xinput83 la_data_out_core[56] vssd vssd vccd vccd input83/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[70\]_B la_buf_enable\[70\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__340__A _340_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_432 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[11\]_A input552/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[13\] input292/X mprj_logic_high_inst/HI[343] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[13\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_buffers\[117\]_A user_to_mprj_in_gates\[117\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__515__A _515_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[106\]_A _570_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[43\]_A _507_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input172_A la_data_out_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[61\]_B la_buf_enable\[61\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input437_A la_oenb_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput410 la_oenb_mprj[11] vssd vssd vccd vccd _603_/A sky130_fd_sc_hd__clkbuf_2
Xinput421 la_oenb_mprj[14] vssd vssd vccd vccd _606_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input33_A la_data_out_core[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput454 la_oenb_mprj[44] vssd vssd vccd vccd _636_/A sky130_fd_sc_hd__clkbuf_2
Xinput432 la_oenb_mprj[24] vssd vssd vccd vccd _616_/A sky130_fd_sc_hd__buf_2
Xinput443 la_oenb_mprj[34] vssd vssd vccd vccd _626_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[81\] _545_/Y la_buf\[81\]/TE vssd vssd vccd vccd output734/A sky130_fd_sc_hd__einvp_4
Xinput465 la_oenb_mprj[54] vssd vssd vccd vccd _646_/A sky130_fd_sc_hd__clkbuf_2
Xinput476 la_oenb_mprj[64] vssd vssd vccd vccd _656_/A sky130_fd_sc_hd__buf_2
Xinput487 la_oenb_mprj[74] vssd vssd vccd vccd _337_/A sky130_fd_sc_hd__buf_2
XANTENNA_input604_A mprj_dat_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput498 la_oenb_mprj[84] vssd vssd vccd vccd _347_/A sky130_fd_sc_hd__buf_4
XFILLER_5_1361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[108\]_A user_to_mprj_in_gates\[108\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__425__A _425_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output656_A output656/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[34\]_A _498_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput906 output906/A vssd vssd vccd vccd la_oenb_core[120] sky130_fd_sc_hd__buf_2
Xoutput928 output928/A vssd vssd vccd vccd la_oenb_core[25] sky130_fd_sc_hd__buf_2
Xoutput917 output917/A vssd vssd vccd vccd la_oenb_core[15] sky130_fd_sc_hd__buf_2
Xoutput939 output939/A vssd vssd vccd vccd la_oenb_core[35] sky130_fd_sc_hd__buf_2
XANTENNA_la_buf_enable\[52\]_B la_buf_enable\[52\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output823_A output823/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[70\] input99/X user_to_mprj_in_gates\[70\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[70\]/Y sky130_fd_sc_hd__nand2_1
XTAP_457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[124\]_B mprj_logic_high_inst/HI[454] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_35_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_clk_buf _391_/Y mprj_clk_buf/TE vssd vssd vccd vccd output1119/A sky130_fd_sc_hd__einvp_4
XFILLER_50_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__335__A _335_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[25\]_A _489_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[43\]_B la_buf_enable\[43\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output1018_A output1018/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[110\]_A _373_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[115\]_B mprj_logic_high_inst/HI[445] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_460_ _460_/A vssd vssd vccd vccd _460_/Y sky130_fd_sc_hd__inv_4
XFILLER_2_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[17\] _609_/Y mprj_logic_high_inst/HI[219] vssd vssd vccd
+ vccd output919/A sky130_fd_sc_hd__einvp_4
X_391_ _391_/A vssd vssd vccd vccd _391_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[39\] _631_/A la_buf_enable\[39\]/B vssd vssd vccd vccd la_buf\[39\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_41_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input387_A la_iena_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[16\]_A _480_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input554_A mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[34\]_B la_buf_enable\[34\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2052 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[3\]_A input321/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[101\]_A _364_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput240 la_data_out_mprj[82] vssd vssd vccd vccd _546_/A sky130_fd_sc_hd__buf_4
Xinput251 la_data_out_mprj[92] vssd vssd vccd vccd _556_/A sky130_fd_sc_hd__clkbuf_2
Xinput262 la_iena_mprj[101] vssd vssd vccd vccd input262/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput295 la_iena_mprj[16] vssd vssd vccd vccd input295/X sky130_fd_sc_hd__clkbuf_1
Xinput273 la_iena_mprj[111] vssd vssd vccd vccd input273/X sky130_fd_sc_hd__clkbuf_1
Xinput284 la_iena_mprj[121] vssd vssd vccd vccd input284/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_in_ena_buf\[106\]_B mprj_logic_high_inst/HI[436] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_589_ _589_/A vssd vssd vccd vccd _589_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_1_1077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[10\]_TE la_buf\[10\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[40\] user_to_mprj_in_gates\[40\]/Y vssd vssd vccd vccd output817/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_53_1945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output773_A output773/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output940_A output940/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput703 output703/A vssd vssd vccd vccd la_data_in_core[53] sky130_fd_sc_hd__buf_2
XFILLER_32_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput736 output736/A vssd vssd vccd vccd la_data_in_core[83] sky130_fd_sc_hd__buf_2
Xoutput725 output725/A vssd vssd vccd vccd la_data_in_core[73] sky130_fd_sc_hd__buf_2
Xoutput714 output714/A vssd vssd vccd vccd la_data_in_core[63] sky130_fd_sc_hd__buf_2
XFILLER_47_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[25\]_B la_buf_enable\[25\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput747 output747/A vssd vssd vccd vccd la_data_in_core[93] sky130_fd_sc_hd__buf_2
XFILLER_47_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput758 output758/A vssd vssd vccd vccd la_data_in_mprj[102] sky130_fd_sc_hd__buf_2
Xoutput769 output769/A vssd vssd vccd vccd la_data_in_mprj[112] sky130_fd_sc_hd__buf_2
XANTENNA_la_buf_enable\[105\]_A_N _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[119\]_TE mprj_logic_high_inst/HI[321] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[94\]_A _357_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[16\]_B la_buf_enable\[16\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[80\] input366/X mprj_logic_high_inst/HI[410] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[80\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[95\]_B mprj_logic_high_inst/HI[425] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input135_A la_data_out_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[33\]_TE la_buf\[33\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_512_ _512_/A vssd vssd vccd vccd _512_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input302_A la_iena_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_443_ _443_/A vssd vssd vccd vccd _443_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_14_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[18\]_TE mprj_logic_high_inst/HI[220] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[85\]_A _348_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[44\] _508_/Y la_buf\[44\]/TE vssd vssd vccd vccd output693/A sky130_fd_sc_hd__einvp_8
X_374_ _374_/A vssd vssd vccd vccd _374_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[116\] input278/X mprj_logic_high_inst/HI[446] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[116\]/B sky130_fd_sc_hd__and2_1
XFILLER_29_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[100\] _564_/Y la_buf\[100\]/TE vssd vssd vccd vccd output628/A sky130_fd_sc_hd__einvp_4
XFILLER_29_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[86\]_B mprj_logic_high_inst/HI[416] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_49_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[88\] user_to_mprj_in_gates\[88\]/Y vssd vssd vccd vccd output869/A
+ sky130_fd_sc_hd__inv_2
XFILLER_48_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output890_A output890/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output988_A output988/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[33\] input58/X user_to_mprj_in_gates\[33\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[33\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[76\]_A _339_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[1\]_TE la_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[10\]_B mprj_logic_high_inst/HI[340] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__613__A _613_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[3\]_A input575/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[77\]_B mprj_logic_high_inst/HI[407] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[56\]_TE la_buf\[56\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[3\]_A input65/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[3\]_A_N _595_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output1085_A output1085/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[67\]_A _330_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__523__A _523_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[84\] _347_/Y mprj_logic_high_inst/HI[286] vssd vssd vccd
+ vccd output993/A sky130_fd_sc_hd__einvp_2
XFILLER_3_935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input252_A la_data_out_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[68\]_B mprj_logic_high_inst/HI[398] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_16 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input517_A mprj_adr_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[107\] _370_/A la_buf_enable\[107\]/B vssd vssd vccd vccd la_buf\[107\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_18_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1016 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[58\]_A _650_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_426_ _426_/A vssd vssd vccd vccd _426_/Y sky130_fd_sc_hd__inv_8
XTAP_1795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_357_ _357_/A vssd vssd vccd vccd _357_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__433__A _433_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output736_A output736/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[79\]_TE la_buf\[79\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output903_A output903/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[59\]_B mprj_logic_high_inst/HI[389] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput4 la_data_out_core[0] vssd vssd vccd vccd input4/X sky130_fd_sc_hd__buf_4
XFILLER_37_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__608__A _608_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[49\]_A _641_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__343__A _343_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2044 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1000_A output1000/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[28\]_TE mprj_dat_buf\[28\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[43\] input325/X mprj_logic_high_inst/HI[373] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[43\]/B sky130_fd_sc_hd__and2_1
XFILLER_3_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__518__A _518_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[7\]_TE mprj_logic_high_inst/HI[209] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_1069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[21\] _613_/A la_buf_enable\[21\]/B vssd vssd vccd vccd la_buf\[21\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_23_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_87 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input63_A la_data_out_core[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input467_A la_oenb_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_ack_buffer user_wb_ack_gate/Y vssd vssd vccd vccd output1011/A sky130_fd_sc_hd__clkinv_8
XFILLER_34_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__428__A _428_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output686_A output686/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_409_ _409_/A vssd vssd vccd vccd _409_/Y sky130_fd_sc_hd__inv_6
XFILLER_14_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output853_A output853/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[63\]_A_N _655_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput1002 output1002/A vssd vssd vccd vccd la_oenb_core[92] sky130_fd_sc_hd__buf_2
Xoutput1024 output1024/A vssd vssd vccd vccd mprj_adr_o_user[20] sky130_fd_sc_hd__buf_2
Xoutput1013 output1013/A vssd vssd vccd vccd mprj_adr_o_user[10] sky130_fd_sc_hd__buf_2
Xoutput1035 output1035/A vssd vssd vccd vccd mprj_adr_o_user[30] sky130_fd_sc_hd__buf_2
XANTENNA_la_buf_enable\[78\]_A_N _341_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[27\]_A _427_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput1046 output1046/A vssd vssd vccd vccd mprj_dat_i_core[10] sky130_fd_sc_hd__buf_2
Xoutput1057 output1057/A vssd vssd vccd vccd mprj_dat_i_core[20] sky130_fd_sc_hd__buf_2
Xoutput1079 output1079/A vssd vssd vccd vccd mprj_dat_o_user[11] sky130_fd_sc_hd__buf_2
Xoutput1068 output1068/A vssd vssd vccd vccd mprj_dat_i_core[30] sky130_fd_sc_hd__buf_2
XFILLER_9_1123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_sel_buf\[2\]_TE mprj_sel_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[107\] input12/X user_to_mprj_in_gates\[107\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[107\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__338__A _338_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[16\]_A_N _608_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[4\]_A _596_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output1048_A output1048/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[18\]_A _418_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[117\] _380_/Y mprj_logic_high_inst/HI[319] vssd vssd vccd
+ vccd output902/A sky130_fd_sc_hd__einvp_2
Xinput603 mprj_dat_o_core[29] vssd vssd vccd vccd _461_/A sky130_fd_sc_hd__clkbuf_2
Xinput625 user_irq_ena[1] vssd vssd vccd vccd input625/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_2003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput614 mprj_iena_wb vssd vssd vccd vccd input614/X sky130_fd_sc_hd__buf_6
XFILLER_47_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[47\] _639_/Y mprj_logic_high_inst/HI[249] vssd vssd vccd
+ vccd output952/A sky130_fd_sc_hd__einvp_2
XFILLER_47_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[69\] _332_/A la_buf_enable\[69\]/B vssd vssd vccd vccd la_buf\[69\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_29_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input215_A la_data_out_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input584_A mprj_dat_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_buffers\[1\]_A user_irq_gates\[1\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[104\] user_to_mprj_in_gates\[104\]/Y vssd vssd vccd vccd
+ output760/A sky130_fd_sc_hd__clkinv_4
XFILLER_43_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[70\] user_to_mprj_in_gates\[70\]/Y vssd vssd vccd vccd output850/A
+ sky130_fd_sc_hd__inv_2
XFILLER_4_1042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[20\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output970_A output970/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[104\]_TE la_buf\[104\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[19\]_TE mprj_adr_buf\[19\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput40 la_data_out_core[17] vssd vssd vccd vccd input40/X sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput73 la_data_out_core[47] vssd vssd vccd vccd input73/X sky130_fd_sc_hd__buf_4
Xinput62 la_data_out_core[37] vssd vssd vccd vccd input62/X sky130_fd_sc_hd__clkbuf_4
Xinput51 la_data_out_core[27] vssd vssd vccd vccd input51/X sky130_fd_sc_hd__clkbuf_4
Xinput95 la_data_out_core[67] vssd vssd vccd vccd input95/X sky130_fd_sc_hd__buf_4
Xinput84 la_data_out_core[57] vssd vssd vccd vccd input84/X sky130_fd_sc_hd__buf_4
XANTENNA__621__A _621_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[3\]_TE mprj_adr_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[3\] _435_/Y mprj_dat_buf\[3\]/TE vssd vssd vccd vccd output1102/A sky130_fd_sc_hd__einvp_8
XFILLER_26_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[11\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[51\]_TE mprj_logic_high_inst/HI[253] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_89 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__531__A _531_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input165_A la_data_out_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[7\]_TE mprj_dat_buf\[7\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput400 la_oenb_mprj[110] vssd vssd vccd vccd _373_/A sky130_fd_sc_hd__clkbuf_4
Xinput411 la_oenb_mprj[120] vssd vssd vccd vccd _383_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input332_A la_iena_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput455 la_oenb_mprj[45] vssd vssd vccd vccd _637_/A sky130_fd_sc_hd__clkbuf_2
Xinput422 la_oenb_mprj[15] vssd vssd vccd vccd _607_/A sky130_fd_sc_hd__buf_2
Xinput433 la_oenb_mprj[25] vssd vssd vccd vccd _617_/A sky130_fd_sc_hd__buf_2
Xinput444 la_oenb_mprj[35] vssd vssd vccd vccd _627_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input26_A la_data_out_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput466 la_oenb_mprj[55] vssd vssd vccd vccd _647_/A sky130_fd_sc_hd__buf_2
Xinput477 la_oenb_mprj[65] vssd vssd vccd vccd _657_/A sky130_fd_sc_hd__buf_2
Xinput488 la_oenb_mprj[75] vssd vssd vccd vccd _338_/A sky130_fd_sc_hd__buf_2
XFILLER_5_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput499 la_oenb_mprj[85] vssd vssd vccd vccd _348_/A sky130_fd_sc_hd__buf_4
Xla_buf\[74\] _538_/Y la_buf\[74\]/TE vssd vssd vccd vccd output726/A sky130_fd_sc_hd__einvp_8
XFILLER_28_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[127\]_TE la_buf\[127\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput907 output907/A vssd vssd vccd vccd la_oenb_core[121] sky130_fd_sc_hd__buf_2
Xoutput918 output918/A vssd vssd vccd vccd la_oenb_core[16] sky130_fd_sc_hd__buf_2
Xoutput929 output929/A vssd vssd vccd vccd la_oenb_core[26] sky130_fd_sc_hd__buf_2
XANTENNA_output649_A output649/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__441__A _441_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output816_A output816/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[63\] input91/X user_to_mprj_in_gates\[63\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[63\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[74\]_TE mprj_logic_high_inst/HI[276] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__616__A _616_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[3\]_A _403_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__351__A _351_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[29\]_A user_wb_dat_gates\[29\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_44_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_390_ _390_/A vssd vssd vccd vccd _390_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1270 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__526__A _526_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input282_A la_iena_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input547_A mprj_adr_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[3\]_B mprj_logic_high_inst/HI[333] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput230 la_data_out_mprj[73] vssd vssd vccd vccd _537_/A sky130_fd_sc_hd__buf_2
Xinput241 la_data_out_mprj[83] vssd vssd vccd vccd _547_/A sky130_fd_sc_hd__buf_4
Xinput252 la_data_out_mprj[93] vssd vssd vccd vccd _557_/A sky130_fd_sc_hd__buf_2
XFILLER_7_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput263 la_iena_mprj[102] vssd vssd vccd vccd input263/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[97\]_TE mprj_logic_high_inst/HI[299] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xinput296 la_iena_mprj[17] vssd vssd vccd vccd input296/X sky130_fd_sc_hd__clkbuf_1
Xinput274 la_iena_mprj[112] vssd vssd vccd vccd input274/X sky130_fd_sc_hd__clkbuf_1
Xinput285 la_iena_mprj[122] vssd vssd vccd vccd input285/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_657_ _657_/A vssd vssd vccd vccd _657_/Y sky130_fd_sc_hd__inv_2
X_588_ _588_/A vssd vssd vccd vccd _588_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__436__A _436_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[33\] user_to_mprj_in_gates\[33\]/Y vssd vssd vccd vccd output809/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output766_A output766/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput726 output726/A vssd vssd vccd vccd la_data_in_core[74] sky130_fd_sc_hd__buf_2
Xoutput704 output704/A vssd vssd vccd vccd la_data_in_core[54] sky130_fd_sc_hd__buf_2
Xoutput715 output715/A vssd vssd vccd vccd la_data_in_core[64] sky130_fd_sc_hd__buf_2
XANTENNA_output933_A output933/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput748 output748/A vssd vssd vccd vccd la_data_in_core[94] sky130_fd_sc_hd__buf_2
Xoutput737 output737/A vssd vssd vccd vccd la_data_in_core[84] sky130_fd_sc_hd__buf_2
XFILLER_47_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput759 output759/A vssd vssd vccd vccd la_data_in_mprj[103] sky130_fd_sc_hd__buf_2
XFILLER_45_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[124\]_B la_buf_enable\[124\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_542 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__346__A _346_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1590 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[93\]_A input124/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output1030_A output1030/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[73\] input358/X mprj_logic_high_inst/HI[403] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[73\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[115\]_B la_buf_enable\[115\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input128_A la_data_out_core[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_511_ _511_/A vssd vssd vccd vccd _511_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_33_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[51\] _643_/A la_buf_enable\[51\]/B vssd vssd vccd vccd la_buf\[51\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_1933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_442_ _442_/A vssd vssd vccd vccd _442_/Y sky130_fd_sc_hd__inv_4
XFILLER_14_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_373_ _373_/A vssd vssd vccd vccd _373_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input497_A la_oenb_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[6\]_A user_wb_dat_gates\[6\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input93_A la_data_out_core[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_A input114/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[37\] _501_/Y la_buf\[37\]/TE vssd vssd vccd vccd output685/A sky130_fd_sc_hd__einvp_8
XFILLER_13_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[109\] input270/X mprj_logic_high_inst/HI[439] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[109\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[9\] input581/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[9\]/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_13_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[9\]_A _473_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_682 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[106\]_B la_buf_enable\[106\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output883_A output883/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[26\] input50/X user_to_mprj_in_gates\[26\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[26\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_53_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[75\]_A input104/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[3\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_81 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[3\]_B user_to_mprj_in_gates\[3\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1078_A output1078/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[66\]_A input94/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[77\] _340_/Y mprj_logic_high_inst/HI[279] vssd vssd vccd
+ vccd output985/A sky130_fd_sc_hd__einvp_4
Xla_buf_enable\[99\] _362_/A la_buf_enable\[99\]/B vssd vssd vccd vccd la_buf\[99\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_46_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[25\] _457_/Y mprj_dat_buf\[25\]/TE vssd vssd vccd vccd output1094/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_28_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input245_A la_data_out_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input412_A la_oenb_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_425_ _425_/A vssd vssd vccd vccd _425_/Y sky130_fd_sc_hd__clkinv_8
XTAP_1796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[104\]_A_N _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_356_ _356_/A vssd vssd vccd vccd _356_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[57\]_A input84/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[20\] _420_/Y mprj_adr_buf\[20\]/TE vssd vssd vccd vccd output1024/A
+ sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[119\]_A_N _382_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output631_A output631/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output729_A output729/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[109\]_TE mprj_logic_high_inst/HI[311] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput5 la_data_out_core[100] vssd vssd vccd vccd input5/X sky130_fd_sc_hd__buf_4
XFILLER_49_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[7\]_A user_to_mprj_in_gates\[7\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_52_604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__624__A _624_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[48\]_A input74/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[5\] _597_/A la_buf_enable\[5\]/B vssd vssd vccd vccd la_buf\[5\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_20_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_578 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[23\]_TE la_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[36\] input317/X mprj_logic_high_inst/HI[366] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[36\]/B sky130_fd_sc_hd__and2_1
XFILLER_3_1482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_11 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__534__A _534_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[14\] _606_/A la_buf_enable\[14\]/B vssd vssd vccd vccd la_buf\[14\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_gates\[123\]_A input30/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[39\]_A input64/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1646 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input195_A la_data_out_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input362_A la_iena_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input56_A la_data_out_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_408_ _408_/A vssd vssd vccd vccd _408_/Y sky130_fd_sc_hd__inv_12
XFILLER_14_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output679_A output679/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__444__A _444_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[114\]_A input20/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_339_ _339_/A vssd vssd vccd vccd _339_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[46\]_TE la_buf\[46\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output846_A output846/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput1003 output1003/A vssd vssd vccd vccd la_oenb_core[93] sky130_fd_sc_hd__buf_2
Xoutput1014 output1014/A vssd vssd vccd vccd mprj_adr_o_user[11] sky130_fd_sc_hd__buf_2
Xuser_to_mprj_in_gates\[93\] input124/X user_to_mprj_in_gates\[93\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[93\]/Y sky130_fd_sc_hd__nand2_1
Xoutput1036 output1036/A vssd vssd vccd vccd mprj_adr_o_user[31] sky130_fd_sc_hd__buf_2
Xoutput1025 output1025/A vssd vssd vccd vccd mprj_adr_o_user[21] sky130_fd_sc_hd__buf_2
XANTENNA_la_buf_enable\[2\]_A_N _594_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput1047 output1047/A vssd vssd vccd vccd mprj_dat_i_core[11] sky130_fd_sc_hd__buf_2
Xoutput1058 output1058/A vssd vssd vccd vccd mprj_dat_i_core[21] sky130_fd_sc_hd__buf_2
XFILLER_44_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput1069 output1069/A vssd vssd vccd vccd mprj_dat_i_core[31] sky130_fd_sc_hd__buf_2
XFILLER_26_1962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__619__A _619_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_82 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__354__A _354_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[105\]_A input10/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_736 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput604 mprj_dat_o_core[2] vssd vssd vccd vccd _434_/A sky130_fd_sc_hd__clkbuf_2
Xinput626 user_irq_ena[2] vssd vssd vccd vccd input626/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_output1110_A output1110/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput615 mprj_sel_o_core[0] vssd vssd vccd vccd _396_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__529__A _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input110_A la_data_out_core[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input208_A la_data_out_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[69\]_TE la_buf\[69\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input577_A mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_49 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__439__A _439_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[63\] user_to_mprj_in_gates\[63\]/Y vssd vssd vccd vccd output842/A
+ sky130_fd_sc_hd__inv_2
XFILLER_1_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output796_A output796/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output963_A output963/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[21\] input563/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[21\]/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_50_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput30 la_data_out_core[123] vssd vssd vccd vccd input30/X sky130_fd_sc_hd__clkbuf_4
XFILLER_15_1663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput63 la_data_out_core[38] vssd vssd vccd vccd input63/X sky130_fd_sc_hd__clkbuf_4
Xinput52 la_data_out_core[28] vssd vssd vccd vccd input52/X sky130_fd_sc_hd__clkbuf_4
Xinput41 la_data_out_core[18] vssd vssd vccd vccd input41/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_mprj_dat_buf\[18\]_TE mprj_dat_buf\[18\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput96 la_data_out_core[68] vssd vssd vccd vccd input96/X sky130_fd_sc_hd__buf_4
Xinput85 la_data_out_core[58] vssd vssd vccd vccd input85/X sky130_fd_sc_hd__buf_4
Xinput74 la_data_out_core[48] vssd vssd vccd vccd input74/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_la_buf_enable\[3\]_B la_buf_enable\[3\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[127\]_A input290/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__349__A _349_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1060_A output1060/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[81\] _344_/A la_buf_enable\[81\]/B vssd vssd vccd vccd la_buf\[81\]/TE
+ sky130_fd_sc_hd__and2b_1
Xinput401 la_oenb_mprj[111] vssd vssd vccd vccd _374_/A sky130_fd_sc_hd__clkbuf_4
Xinput412 la_oenb_mprj[121] vssd vssd vccd vccd _384_/A sky130_fd_sc_hd__buf_2
XANTENNA_input158_A la_data_out_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[118\]_A input280/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput423 la_oenb_mprj[16] vssd vssd vccd vccd _608_/A sky130_fd_sc_hd__clkbuf_2
Xinput434 la_oenb_mprj[26] vssd vssd vccd vccd _618_/A sky130_fd_sc_hd__buf_2
Xinput445 la_oenb_mprj[36] vssd vssd vccd vccd _628_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput467 la_oenb_mprj[56] vssd vssd vccd vccd _648_/A sky130_fd_sc_hd__clkbuf_2
Xinput456 la_oenb_mprj[46] vssd vssd vccd vccd _638_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_input325_A la_iena_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput478 la_oenb_mprj[66] vssd vssd vccd vccd _329_/A sky130_fd_sc_hd__buf_4
XANTENNA_input19_A la_data_out_core[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[62\]_A_N _654_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput489 la_oenb_mprj[76] vssd vssd vccd vccd _339_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[67\] _531_/Y la_buf\[67\]/TE vssd vssd vccd vccd output718/A sky130_fd_sc_hd__einvp_8
XFILLER_16_445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[77\]_A_N _340_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput908 output908/A vssd vssd vccd vccd la_oenb_core[122] sky130_fd_sc_hd__buf_2
Xoutput919 output919/A vssd vssd vccd vccd la_oenb_core[17] sky130_fd_sc_hd__buf_2
Xla_buf\[123\] _587_/Y la_buf\[123\]/TE vssd vssd vccd vccd output653/A sky130_fd_sc_hd__einvp_2
XFILLER_45_2324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[15\]_A_N _607_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output711_A output711/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[109\]_A input270/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output809_A output809/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[56\] input83/X user_to_mprj_in_gates\[56\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[56\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_26_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[40\]_A input322/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_2063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__632__A _632_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_319 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[31\]_A input312/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__542__A _542_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input275_A la_iena_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input442_A la_oenb_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[98\]_A input385/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput220 la_data_out_mprj[64] vssd vssd vccd vccd _528_/A sky130_fd_sc_hd__buf_2
Xinput231 la_data_out_mprj[74] vssd vssd vccd vccd _538_/A sky130_fd_sc_hd__clkbuf_2
Xinput242 la_data_out_mprj[84] vssd vssd vccd vccd _548_/A sky130_fd_sc_hd__buf_4
Xinput253 la_data_out_mprj[94] vssd vssd vccd vccd _558_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput297 la_iena_mprj[18] vssd vssd vccd vccd input297/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput264 la_iena_mprj[103] vssd vssd vccd vccd input264/X sky130_fd_sc_hd__clkbuf_1
Xinput275 la_iena_mprj[113] vssd vssd vccd vccd input275/X sky130_fd_sc_hd__clkbuf_1
Xinput286 la_iena_mprj[123] vssd vssd vccd vccd input286/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1024 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_656_ _656_/A vssd vssd vccd vccd _656_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_587_ _587_/A vssd vssd vccd vccd _587_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[22\]_A input302/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output661_A output661/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[26\] user_to_mprj_in_gates\[26\]/Y vssd vssd vccd vccd output801/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA__452__A _452_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output759_A output759/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput727 output727/A vssd vssd vccd vccd la_data_in_core[75] sky130_fd_sc_hd__buf_2
Xoutput716 output716/A vssd vssd vccd vccd la_data_in_core[65] sky130_fd_sc_hd__buf_2
Xoutput705 output705/A vssd vssd vccd vccd la_data_in_core[55] sky130_fd_sc_hd__buf_2
Xoutput749 output749/A vssd vssd vccd vccd la_data_in_core[95] sky130_fd_sc_hd__buf_2
Xoutput738 output738/A vssd vssd vccd vccd la_data_in_core[85] sky130_fd_sc_hd__buf_2
XANTENNA_output926_A output926/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[89\]_A input375/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[41\]_TE mprj_logic_high_inst/HI[243] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XTAP_278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__627__A _627_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[13\]_A input292/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[93\]_B user_to_mprj_in_gates\[93\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__362__A _362_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[117\]_TE la_buf\[117\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output1023_A output1023/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[66\] input350/X mprj_logic_high_inst/HI[396] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[66\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2012 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_510_ _510_/A vssd vssd vccd vccd _510_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[0\]_A input624/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[22\] _614_/Y mprj_logic_high_inst/HI[224] vssd vssd vccd
+ vccd output925/A sky130_fd_sc_hd__einvp_4
XANTENNA__537__A _537_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[44\] _636_/A la_buf_enable\[44\]/B vssd vssd vccd vccd la_buf\[44\]/TE
+ sky130_fd_sc_hd__and2b_1
X_441_ _441_/A vssd vssd vccd vccd _441_/Y sky130_fd_sc_hd__inv_6
Xuser_to_mprj_oen_buffers\[4\] _596_/Y mprj_logic_high_inst/HI[206] vssd vssd vccd
+ vccd output955/A sky130_fd_sc_hd__einvp_4
XFILLER_2_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_372_ _372_/A vssd vssd vccd vccd _372_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_B user_to_mprj_in_gates\[84\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_input392_A la_oenb_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input86_A la_data_out_core[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[64\]_TE mprj_logic_high_inst/HI[266] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_639_ _639_/A vssd vssd vccd vccd _639_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__447__A _447_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output876_A output876/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[19\] input42/X user_to_mprj_in_gates\[19\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[19\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_gates\[75\]_B user_to_mprj_in_gates\[75\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[29\] user_wb_dat_gates\[29\]/Y vssd vssd vccd vccd output1066/A
+ sky130_fd_sc_hd__inv_6
XFILLER_47_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[60\]_A user_to_mprj_in_gates\[60\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__357__A _357_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[66\]_B user_to_mprj_in_gates\[66\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[87\]_TE mprj_logic_high_inst/HI[289] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[18\] _450_/Y mprj_dat_buf\[18\]/TE vssd vssd vccd vccd output1086/A
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input238_A la_data_out_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[51\]_A user_to_mprj_in_gates\[51\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_input140_A la_data_out_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input405_A la_oenb_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_424_ _424_/A vssd vssd vccd vccd _424_/Y sky130_fd_sc_hd__inv_12
XTAP_1764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_355_ _355_/A vssd vssd vccd vccd _355_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[121\] input284/X mprj_logic_high_inst/HI[451] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[121\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[57\]_B user_to_mprj_in_gates\[57\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[91\]_A _555_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[13\] _413_/Y mprj_adr_buf\[13\]/TE vssd vssd vccd vccd output1016/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_48_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[127\] user_to_mprj_in_gates\[127\]/Y vssd vssd vccd vccd
+ output785/A sky130_fd_sc_hd__clkinv_4
XFILLER_9_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[93\] user_to_mprj_in_gates\[93\]/Y vssd vssd vccd vccd output875/A
+ sky130_fd_sc_hd__inv_2
XFILLER_42_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[42\]_A user_to_mprj_in_gates\[42\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xinput6 la_data_out_core[101] vssd vssd vccd vccd input6/X sky130_fd_sc_hd__buf_4
XFILLER_42_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output993_A output993/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_buffers\[3\] user_wb_dat_gates\[3\]/Y vssd vssd vccd vccd output1070/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_33_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[48\]_B user_to_mprj_in_gates\[48\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[82\]_A _546_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__640__A _640_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[0\] input4/X user_to_mprj_in_gates\[0\]/B vssd vssd vccd vccd
+ user_to_mprj_in_gates\[0\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[33\]_A user_to_mprj_in_gates\[33\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[29\] input309/X mprj_logic_high_inst/HI[359] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[29\]/B sky130_fd_sc_hd__and2_1
XFILLER_3_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1090_A output1090/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_79 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_45 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_23 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[123\]_B user_to_mprj_in_gates\[123\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[39\]_B user_to_mprj_in_gates\[39\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[73\]_A _537_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input188_A la_data_out_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[91\]_B la_buf_enable\[91\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__550__A _550_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input355_A la_iena_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input49_A la_data_out_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[24\]_A user_to_mprj_in_gates\[24\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_input522_A mprj_adr_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[97\] _561_/Y la_buf\[97\]/TE vssd vssd vccd vccd output751/A sky130_fd_sc_hd__einvp_2
Xla_buf_enable\[112\] _375_/A la_buf_enable\[112\]/B vssd vssd vccd vccd la_buf\[112\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_19_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[2\] input310/X mprj_logic_high_inst/HI[332] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[2\]/B sky130_fd_sc_hd__and2_1
XFILLER_4_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[127\]_A _591_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_407_ _407_/A vssd vssd vccd vccd _407_/Y sky130_fd_sc_hd__inv_12
X_338_ _338_/A vssd vssd vccd vccd _338_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[114\]_B user_to_mprj_in_gates\[114\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[64\]_A _528_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output741_A output741/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[82\]_B la_buf_enable\[82\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput1004 output1004/A vssd vssd vccd vccd la_oenb_core[94] sky130_fd_sc_hd__buf_2
Xoutput1015 output1015/A vssd vssd vccd vccd mprj_adr_o_user[12] sky130_fd_sc_hd__buf_2
XFILLER_48_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__460__A _460_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output839_A output839/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput1026 output1026/A vssd vssd vccd vccd mprj_adr_o_user[22] sky130_fd_sc_hd__buf_2
Xoutput1037 output1037/A vssd vssd vccd vccd mprj_adr_o_user[3] sky130_fd_sc_hd__buf_2
XFILLER_44_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput1048 output1048/A vssd vssd vccd vccd mprj_dat_i_core[12] sky130_fd_sc_hd__buf_2
XFILLER_9_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[86\] input116/X user_to_mprj_in_gates\[86\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[86\]/Y sky130_fd_sc_hd__nand2_1
Xoutput1059 output1059/A vssd vssd vccd vccd mprj_dat_i_core[22] sky130_fd_sc_hd__buf_2
XFILLER_9_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[15\]_A user_to_mprj_in_gates\[15\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_49_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_72 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[23\]_A input565/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2346 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__635__A _635_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[118\]_A _582_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[105\]_B user_to_mprj_in_gates\[105\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[55\]_A _519_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[73\]_B la_buf_enable\[73\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__370__A _370_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1738 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput616 mprj_sel_o_core[1] vssd vssd vccd vccd _397_/A sky130_fd_sc_hd__clkbuf_2
Xinput605 mprj_dat_o_core[30] vssd vssd vccd vccd _462_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_output1103_A output1103/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[103\]_A_N _366_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[14\]_A input555/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_936 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[118\]_A_N _381_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input103_A la_data_out_core[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[109\]_A _573_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__545__A _545_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[0\] user_to_mprj_in_gates\[0\]/Y vssd vssd vccd vccd output755/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_36_2281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[46\]_A _510_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input472_A la_oenb_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[64\]_B la_buf_enable\[64\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[12\] _476_/Y la_buf\[12\]/TE vssd vssd vccd vccd output658/A sky130_fd_sc_hd__einvp_8
Xla_buf\[8\] _472_/Y la_buf\[8\]/TE vssd vssd vccd vccd output743/A sky130_fd_sc_hd__einvp_8
XFILLER_10_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[5\] _405_/Y mprj_adr_buf\[5\]/TE vssd vssd vccd vccd output1039/A sky130_fd_sc_hd__einvp_8
XFILLER_47_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[13\]_TE la_buf\[13\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[56\] user_to_mprj_in_gates\[56\]/Y vssd vssd vccd vccd output834/A
+ sky130_fd_sc_hd__clkinv_4
XTAP_2092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output691_A output691/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__455__A _455_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output789_A output789/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[37\]_A _501_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput31 la_data_out_core[124] vssd vssd vccd vccd input31/X sky130_fd_sc_hd__clkbuf_4
XFILLER_50_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput20 la_data_out_core[114] vssd vssd vccd vccd input20/X sky130_fd_sc_hd__clkbuf_4
Xuser_wb_dat_gates\[14\] input555/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[14\]/Y
+ sky130_fd_sc_hd__nand2_2
XANTENNA_output956_A output956/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput64 la_data_out_core[39] vssd vssd vccd vccd input64/X sky130_fd_sc_hd__clkbuf_4
Xinput53 la_data_out_core[29] vssd vssd vccd vccd input53/X sky130_fd_sc_hd__clkbuf_4
Xinput42 la_data_out_core[19] vssd vssd vccd vccd input42/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_la_buf_enable\[55\]_B la_buf_enable\[55\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput97 la_data_out_core[69] vssd vssd vccd vccd input97/X sky130_fd_sc_hd__buf_4
Xinput86 la_data_out_core[59] vssd vssd vccd vccd input86/X sky130_fd_sc_hd__buf_4
Xinput75 la_data_out_core[49] vssd vssd vccd vccd input75/X sky130_fd_sc_hd__buf_4
XFILLER_48_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[11\] user_wb_dat_gates\[11\]/Y vssd vssd vccd vccd output1047/A
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_user_to_mprj_oen_buffers\[122\]_A _385_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[127\]_B mprj_logic_high_inst/HI[457] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[112\] input18/X user_to_mprj_in_gates\[112\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[112\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__365__A _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[28\]_A _492_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[46\]_B la_buf_enable\[46\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output1053_A output1053/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[96\] input383/X mprj_logic_high_inst/HI[426] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[96\]/B sky130_fd_sc_hd__and2_1
XFILLER_27_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[113\]_A _376_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[122\] _385_/Y mprj_logic_high_inst/HI[324] vssd vssd vccd
+ vccd output908/A sky130_fd_sc_hd__einvp_4
Xmprj_sel_buf\[3\] _399_/Y mprj_sel_buf\[3\]/TE vssd vssd vccd vccd output1112/A sky130_fd_sc_hd__einvp_8
Xinput402 la_oenb_mprj[112] vssd vssd vccd vccd _375_/A sky130_fd_sc_hd__buf_2
XFILLER_7_1618 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[52\] _644_/Y mprj_logic_high_inst/HI[254] vssd vssd vccd
+ vccd output958/A sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[118\]_B mprj_logic_high_inst/HI[448] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xinput424 la_oenb_mprj[17] vssd vssd vccd vccd _609_/A sky130_fd_sc_hd__buf_2
Xinput435 la_oenb_mprj[27] vssd vssd vccd vccd _619_/A sky130_fd_sc_hd__buf_2
Xinput446 la_oenb_mprj[37] vssd vssd vccd vccd _629_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput413 la_oenb_mprj[122] vssd vssd vccd vccd _385_/A sky130_fd_sc_hd__buf_2
XFILLER_7_1629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[74\] _337_/A la_buf_enable\[74\]/B vssd vssd vccd vccd la_buf\[74\]/TE
+ sky130_fd_sc_hd__and2b_1
Xinput468 la_oenb_mprj[57] vssd vssd vccd vccd _649_/A sky130_fd_sc_hd__buf_2
Xinput457 la_oenb_mprj[47] vssd vssd vccd vccd _639_/A sky130_fd_sc_hd__buf_4
Xinput479 la_oenb_mprj[67] vssd vssd vccd vccd _330_/A sky130_fd_sc_hd__buf_2
XFILLER_5_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input318_A la_iena_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input220_A la_data_out_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[36\]_TE la_buf\[36\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[1\]_A_N _593_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[19\]_A _483_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[37\]_B la_buf_enable\[37\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput909 output909/A vssd vssd vccd vccd la_oenb_core[123] sky130_fd_sc_hd__buf_2
XFILLER_32_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[116\] _580_/Y la_buf\[116\]/TE vssd vssd vccd vccd output645/A sky130_fd_sc_hd__einvp_4
XANTENNA_user_to_mprj_in_ena_buf\[6\]_A input354/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[104\]_A _367_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_clk2_buf_A _392_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[109\]_B mprj_logic_high_inst/HI[439] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output704_A output704/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[49\] input75/X user_to_mprj_in_gates\[49\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[49\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[40\]_B mprj_logic_high_inst/HI[370] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2020 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[4\]_TE la_buf\[4\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[28\]_B la_buf_enable\[28\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[30\]_A _622_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[59\]_TE la_buf\[59\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[97\]_A _360_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[11\] input282/X mprj_logic_high_inst/HI[341] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[11\]/B sky130_fd_sc_hd__and2_1
XFILLER_43_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[31\]_B mprj_logic_high_inst/HI[361] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[19\]_B la_buf_enable\[19\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input170_A la_data_out_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[21\]_A _613_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input268_A la_iena_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[98\]_B mprj_logic_high_inst/HI[428] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput210 la_data_out_mprj[55] vssd vssd vccd vccd _519_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_input435_A la_oenb_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input31_A la_data_out_core[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput221 la_data_out_mprj[65] vssd vssd vccd vccd _529_/A sky130_fd_sc_hd__clkbuf_2
Xinput232 la_data_out_mprj[75] vssd vssd vccd vccd _539_/A sky130_fd_sc_hd__buf_2
Xinput243 la_data_out_mprj[85] vssd vssd vccd vccd _549_/A sky130_fd_sc_hd__buf_4
Xinput254 la_data_out_mprj[95] vssd vssd vccd vccd _559_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput265 la_iena_mprj[104] vssd vssd vccd vccd input265/X sky130_fd_sc_hd__clkbuf_1
Xinput276 la_iena_mprj[114] vssd vssd vccd vccd input276/X sky130_fd_sc_hd__clkbuf_1
Xinput287 la_iena_mprj[124] vssd vssd vccd vccd input287/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input602_A mprj_dat_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput298 la_iena_mprj[19] vssd vssd vccd vccd input298/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_1014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_655_ _655_/A vssd vssd vccd vccd _655_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_1_1047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[88\]_A _351_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_586_ _586_/A vssd vssd vccd vccd _586_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[22\]_B mprj_logic_high_inst/HI[352] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_31_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output654_A output654/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[19\] user_to_mprj_in_gates\[19\]/Y vssd vssd vccd vccd output793/A
+ sky130_fd_sc_hd__clkinv_4
Xoutput717 output717/A vssd vssd vccd vccd la_data_in_core[66] sky130_fd_sc_hd__buf_2
Xoutput706 output706/A vssd vssd vccd vccd la_data_in_core[56] sky130_fd_sc_hd__buf_2
XFILLER_32_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput739 output739/A vssd vssd vccd vccd la_data_in_core[86] sky130_fd_sc_hd__buf_2
Xoutput728 output728/A vssd vssd vccd vccd la_data_in_core[76] sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_oen_buffers\[12\]_A _604_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output919_A output919/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output821_A output821/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[89\]_B mprj_logic_high_inst/HI[419] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[79\]_A _342_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_repeater1125_A repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[13\]_B mprj_logic_high_inst/HI[343] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__643__A _643_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[6\]_A input578/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[61\]_A_N _653_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[76\]_A_N _339_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1016_A output1016/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[6\]_A input98/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[59\] input342/X mprj_logic_high_inst/HI[389] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[59\]/B sky130_fd_sc_hd__and2_1
XFILLER_2_2024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_irq_ena_buf\[0\]_B user_irq_ena_buf\[0\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_440_ _440_/A vssd vssd vccd vccd _440_/Y sky130_fd_sc_hd__clkinv_4
XTAP_1968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[15\] _607_/Y mprj_logic_high_inst/HI[217] vssd vssd vccd
+ vccd output917/A sky130_fd_sc_hd__einvp_4
X_371_ _371_/A vssd vssd vccd vccd _371_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[37\] _629_/A la_buf_enable\[37\]/B vssd vssd vccd vccd la_buf\[37\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_1979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[14\]_A_N _606_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__553__A _553_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input385_A la_iena_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[29\]_A_N _621_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input79_A la_data_out_core[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input552_A mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1936 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_638_ _638_/A vssd vssd vccd vccd _638_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_569_ _569_/A vssd vssd vccd vccd _569_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__463__A _463_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output771_A output771/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output869_A output869/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__638__A _638_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[30\]_A _462_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__373__A _373_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input133_A la_data_out_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__548__A _548_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input300_A la_iena_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_423_ _423_/A vssd vssd vccd vccd _423_/Y sky130_fd_sc_hd__inv_8
XTAP_1765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_dat_buf\[21\]_A _453_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[42\] _506_/Y la_buf\[42\]/TE vssd vssd vccd vccd output691/A sky130_fd_sc_hd__einvp_8
XFILLER_41_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_354_ _354_/A vssd vssd vccd vccd _354_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[114\] input276/X mprj_logic_high_inst/HI[444] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[114\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[31\]_TE mprj_logic_high_inst/HI[233] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput7 la_data_out_core[102] vssd vssd vccd vccd input7/X sky130_fd_sc_hd__buf_4
XFILLER_37_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[86\] user_to_mprj_in_gates\[86\]/Y vssd vssd vccd vccd output867/A
+ sky130_fd_sc_hd__inv_2
XFILLER_42_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__458__A _458_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output986_A output986/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[107\]_TE la_buf\[107\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[31\] input56/X user_to_mprj_in_gates\[31\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[31\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[12\]_A _444_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[6\]_TE mprj_adr_buf\[6\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__368__A _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[7\]_A _599_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_buffers\[10\]_A user_wb_dat_gates\[10\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_output1083_A output1083/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[54\]_TE mprj_logic_high_inst/HI[256] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[82\] _345_/Y mprj_logic_high_inst/HI[284] vssd vssd vccd
+ vccd output991/A sky130_fd_sc_hd__einvp_2
XFILLER_10_1957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[30\] _462_/Y mprj_dat_buf\[30\]/TE vssd vssd vccd vccd output1100/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input348_A la_iena_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input250_A la_data_out_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input515_A la_oenb_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[105\] _368_/A la_buf_enable\[105\]/B vssd vssd vccd vccd la_buf\[105\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_2252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_406_ _406_/A vssd vssd vccd vccd _406_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_41_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_337_ _337_/A vssd vssd vccd vccd _337_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput1005 output1005/A vssd vssd vccd vccd la_oenb_core[95] sky130_fd_sc_hd__buf_2
XANTENNA_output734_A output734/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput1038 output1038/A vssd vssd vccd vccd mprj_adr_o_user[4] sky130_fd_sc_hd__buf_2
Xoutput1027 output1027/A vssd vssd vccd vccd mprj_adr_o_user[23] sky130_fd_sc_hd__buf_2
Xoutput1016 output1016/A vssd vssd vccd vccd mprj_adr_o_user[13] sky130_fd_sc_hd__buf_2
XFILLER_48_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput1049 output1049/A vssd vssd vccd vccd mprj_dat_i_core[13] sky130_fd_sc_hd__buf_2
XFILLER_48_1666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output901_A output901/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[79\] input108/X user_to_mprj_in_gates\[79\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[79\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[92\]_TE la_buf\[92\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[23\]_B repeater1125/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[77\]_TE mprj_logic_high_inst/HI[279] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__651__A _651_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput617 mprj_sel_o_core[2] vssd vssd vccd vccd _398_/A sky130_fd_sc_hd__buf_2
Xinput606 mprj_dat_o_core[31] vssd vssd vccd vccd _463_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_1660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[14\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[41\] input323/X mprj_logic_high_inst/HI[371] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[41\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_cyc_buf_TE mprj_cyc_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input298_A la_iena_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__561__A _561_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input61_A la_data_out_core[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input465_A la_oenb_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[49\] user_to_mprj_in_gates\[49\]/Y vssd vssd vccd vccd output826/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_50_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output684_A output684/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput21 la_data_out_core[115] vssd vssd vccd vccd input21/X sky130_fd_sc_hd__clkbuf_4
Xinput10 la_data_out_core[105] vssd vssd vccd vccd input10/X sky130_fd_sc_hd__buf_4
XFILLER_35_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output851_A output851/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput32 la_data_out_core[125] vssd vssd vccd vccd input32/X sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output949_A output949/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput43 la_data_out_core[1] vssd vssd vccd vccd input43/X sky130_fd_sc_hd__buf_4
Xinput54 la_data_out_core[2] vssd vssd vccd vccd input54/X sky130_fd_sc_hd__buf_4
XANTENNA__471__A _471_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput98 la_data_out_core[6] vssd vssd vccd vccd input98/X sky130_fd_sc_hd__buf_4
Xinput76 la_data_out_core[4] vssd vssd vccd vccd input76/X sky130_fd_sc_hd__buf_4
Xinput87 la_data_out_core[5] vssd vssd vccd vccd input87/X sky130_fd_sc_hd__buf_4
Xinput65 la_data_out_core[3] vssd vssd vccd vccd input65/X sky130_fd_sc_hd__buf_4
XFILLER_7_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[105\] input10/X user_to_mprj_in_gates\[105\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[105\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA__646__A _646_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj2_logic_high_inst mprj2_pwrgood/A vccd2_uq6 vssd2_uq5 mprj2_logic_high
XANTENNA_mprj_adr_buf\[6\]_A _406_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__381__A _381_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[89\] input375/X mprj_logic_high_inst/HI[419] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[89\]/B sky130_fd_sc_hd__and2_1
XANTENNA_output1046_A output1046/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[115\] _378_/Y mprj_logic_high_inst/HI[317] vssd vssd vccd
+ vccd output900/A sky130_fd_sc_hd__einvp_4
Xinput403 la_oenb_mprj[113] vssd vssd vccd vccd _376_/A sky130_fd_sc_hd__clkbuf_4
Xinput425 la_oenb_mprj[18] vssd vssd vccd vccd _610_/A sky130_fd_sc_hd__clkbuf_2
Xinput436 la_oenb_mprj[28] vssd vssd vccd vccd _620_/A sky130_fd_sc_hd__buf_2
Xinput414 la_oenb_mprj[123] vssd vssd vccd vccd _386_/A sky130_fd_sc_hd__clkbuf_4
Xinput458 la_oenb_mprj[48] vssd vssd vccd vccd _640_/A sky130_fd_sc_hd__clkbuf_2
Xinput447 la_oenb_mprj[38] vssd vssd vccd vccd _630_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput469 la_oenb_mprj[58] vssd vssd vccd vccd _650_/A sky130_fd_sc_hd__clkbuf_2
Xuser_to_mprj_oen_buffers\[45\] _637_/Y mprj_logic_high_inst/HI[247] vssd vssd vccd
+ vccd output950/A sky130_fd_sc_hd__einvp_4
Xla_buf_enable\[67\] _330_/A la_buf_enable\[67\]/B vssd vssd vccd vccd la_buf\[67\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_5_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1354 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input213_A la_data_out_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__556__A _556_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input582_A mprj_dat_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_rstn_buf_TE mprj_rstn_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[6\]_B mprj_logic_high_inst/HI[336] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[109\] _573_/Y la_buf\[109\]/TE vssd vssd vccd vccd output637/A sky130_fd_sc_hd__einvp_2
XTAP_439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[102\] user_to_mprj_in_gates\[102\]/Y vssd vssd vccd vccd
+ output758/A sky130_fd_sc_hd__clkinv_4
XFILLER_23_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output899_A output899/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__466__A _466_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[102\]_A_N _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[117\]_A_N _380_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[127\]_B la_buf_enable\[127\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_dat_buf\[1\] _433_/Y mprj_dat_buf\[1\]/TE vssd vssd vccd vccd output1088/A sky130_fd_sc_hd__einvp_8
XTAP_951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_logic_high_inst mprj_rstn_buf/TE la_buf_enable\[26\]/B la_buf_enable\[27\]/B
+ la_buf_enable\[28\]/B la_buf_enable\[29\]/B la_buf_enable\[30\]/B la_buf_enable\[31\]/B
+ la_buf_enable\[32\]/B la_buf_enable\[33\]/B la_buf_enable\[34\]/B la_buf_enable\[35\]/B
+ mprj_adr_buf\[0\]/TE la_buf_enable\[36\]/B la_buf_enable\[37\]/B la_buf_enable\[38\]/B
+ la_buf_enable\[39\]/B la_buf_enable\[40\]/B la_buf_enable\[41\]/B la_buf_enable\[42\]/B
+ la_buf_enable\[43\]/B la_buf_enable\[44\]/B la_buf_enable\[45\]/B mprj_adr_buf\[1\]/TE
+ la_buf_enable\[46\]/B la_buf_enable\[47\]/B la_buf_enable\[48\]/B la_buf_enable\[49\]/B
+ la_buf_enable\[50\]/B la_buf_enable\[51\]/B la_buf_enable\[52\]/B la_buf_enable\[53\]/B
+ la_buf_enable\[54\]/B la_buf_enable\[55\]/B mprj_adr_buf\[2\]/TE la_buf_enable\[56\]/B
+ la_buf_enable\[57\]/B la_buf_enable\[58\]/B la_buf_enable\[59\]/B la_buf_enable\[60\]/B
+ la_buf_enable\[61\]/B la_buf_enable\[62\]/B la_buf_enable\[63\]/B la_buf_enable\[64\]/B
+ la_buf_enable\[65\]/B mprj_adr_buf\[3\]/TE la_buf_enable\[66\]/B la_buf_enable\[67\]/B
+ la_buf_enable\[68\]/B la_buf_enable\[69\]/B la_buf_enable\[70\]/B la_buf_enable\[71\]/B
+ la_buf_enable\[72\]/B la_buf_enable\[73\]/B la_buf_enable\[74\]/B la_buf_enable\[75\]/B
+ mprj_adr_buf\[4\]/TE la_buf_enable\[76\]/B la_buf_enable\[77\]/B la_buf_enable\[78\]/B
+ la_buf_enable\[79\]/B la_buf_enable\[80\]/B la_buf_enable\[81\]/B la_buf_enable\[82\]/B
+ la_buf_enable\[83\]/B la_buf_enable\[84\]/B la_buf_enable\[85\]/B mprj_adr_buf\[5\]/TE
+ la_buf_enable\[86\]/B la_buf_enable\[87\]/B la_buf_enable\[88\]/B la_buf_enable\[89\]/B
+ la_buf_enable\[90\]/B la_buf_enable\[91\]/B la_buf_enable\[92\]/B la_buf_enable\[93\]/B
+ la_buf_enable\[94\]/B la_buf_enable\[95\]/B mprj_adr_buf\[6\]/TE la_buf_enable\[96\]/B
+ la_buf_enable\[97\]/B la_buf_enable\[98\]/B la_buf_enable\[99\]/B la_buf_enable\[100\]/B
+ la_buf_enable\[101\]/B la_buf_enable\[102\]/B la_buf_enable\[103\]/B la_buf_enable\[104\]/B
+ la_buf_enable\[105\]/B mprj_adr_buf\[7\]/TE la_buf_enable\[106\]/B la_buf_enable\[107\]/B
+ la_buf_enable\[108\]/B la_buf_enable\[109\]/B la_buf_enable\[110\]/B la_buf_enable\[111\]/B
+ la_buf_enable\[112\]/B la_buf_enable\[113\]/B la_buf_enable\[114\]/B la_buf_enable\[115\]/B
+ mprj_adr_buf\[8\]/TE la_buf_enable\[116\]/B la_buf_enable\[117\]/B la_buf_enable\[118\]/B
+ la_buf_enable\[119\]/B la_buf_enable\[120\]/B la_buf_enable\[121\]/B la_buf_enable\[122\]/B
+ la_buf_enable\[123\]/B la_buf_enable\[124\]/B la_buf_enable\[125\]/B mprj_adr_buf\[9\]/TE
+ mprj_clk_buf/TE la_buf_enable\[126\]/B la_buf_enable\[127\]/B mprj_logic_high_inst/HI[202]
+ mprj_logic_high_inst/HI[203] mprj_logic_high_inst/HI[204] mprj_logic_high_inst/HI[205]
+ mprj_logic_high_inst/HI[206] mprj_logic_high_inst/HI[207] mprj_logic_high_inst/HI[208]
+ mprj_logic_high_inst/HI[209] mprj_adr_buf\[10\]/TE mprj_logic_high_inst/HI[210]
+ mprj_logic_high_inst/HI[211] mprj_logic_high_inst/HI[212] mprj_logic_high_inst/HI[213]
+ mprj_logic_high_inst/HI[214] mprj_logic_high_inst/HI[215] mprj_logic_high_inst/HI[216]
+ mprj_logic_high_inst/HI[217] mprj_logic_high_inst/HI[218] mprj_logic_high_inst/HI[219]
+ mprj_adr_buf\[11\]/TE mprj_logic_high_inst/HI[220] mprj_logic_high_inst/HI[221]
+ mprj_logic_high_inst/HI[222] mprj_logic_high_inst/HI[223] mprj_logic_high_inst/HI[224]
+ mprj_logic_high_inst/HI[225] mprj_logic_high_inst/HI[226] mprj_logic_high_inst/HI[227]
+ mprj_logic_high_inst/HI[228] mprj_logic_high_inst/HI[229] mprj_adr_buf\[12\]/TE
+ mprj_logic_high_inst/HI[230] mprj_logic_high_inst/HI[231] mprj_logic_high_inst/HI[232]
+ mprj_logic_high_inst/HI[233] mprj_logic_high_inst/HI[234] mprj_logic_high_inst/HI[235]
+ mprj_logic_high_inst/HI[236] mprj_logic_high_inst/HI[237] mprj_logic_high_inst/HI[238]
+ mprj_logic_high_inst/HI[239] mprj_adr_buf\[13\]/TE mprj_logic_high_inst/HI[240]
+ mprj_logic_high_inst/HI[241] mprj_logic_high_inst/HI[242] mprj_logic_high_inst/HI[243]
+ mprj_logic_high_inst/HI[244] mprj_logic_high_inst/HI[245] mprj_logic_high_inst/HI[246]
+ mprj_logic_high_inst/HI[247] mprj_logic_high_inst/HI[248] mprj_logic_high_inst/HI[249]
+ mprj_adr_buf\[14\]/TE mprj_logic_high_inst/HI[250] mprj_logic_high_inst/HI[251]
+ mprj_logic_high_inst/HI[252] mprj_logic_high_inst/HI[253] mprj_logic_high_inst/HI[254]
+ mprj_logic_high_inst/HI[255] mprj_logic_high_inst/HI[256] mprj_logic_high_inst/HI[257]
+ mprj_logic_high_inst/HI[258] mprj_logic_high_inst/HI[259] mprj_adr_buf\[15\]/TE
+ mprj_logic_high_inst/HI[260] mprj_logic_high_inst/HI[261] mprj_logic_high_inst/HI[262]
+ mprj_logic_high_inst/HI[263] mprj_logic_high_inst/HI[264] mprj_logic_high_inst/HI[265]
+ mprj_logic_high_inst/HI[266] mprj_logic_high_inst/HI[267] mprj_logic_high_inst/HI[268]
+ mprj_logic_high_inst/HI[269] mprj_adr_buf\[16\]/TE mprj_logic_high_inst/HI[270]
+ mprj_logic_high_inst/HI[271] mprj_logic_high_inst/HI[272] mprj_logic_high_inst/HI[273]
+ mprj_logic_high_inst/HI[274] mprj_logic_high_inst/HI[275] mprj_logic_high_inst/HI[276]
+ mprj_logic_high_inst/HI[277] mprj_logic_high_inst/HI[278] mprj_logic_high_inst/HI[279]
+ mprj_adr_buf\[17\]/TE mprj_logic_high_inst/HI[280] mprj_logic_high_inst/HI[281]
+ mprj_logic_high_inst/HI[282] mprj_logic_high_inst/HI[283] mprj_logic_high_inst/HI[284]
+ mprj_logic_high_inst/HI[285] mprj_logic_high_inst/HI[286] mprj_logic_high_inst/HI[287]
+ mprj_logic_high_inst/HI[288] mprj_logic_high_inst/HI[289] mprj_adr_buf\[18\]/TE
+ mprj_logic_high_inst/HI[290] mprj_logic_high_inst/HI[291] mprj_logic_high_inst/HI[292]
+ mprj_logic_high_inst/HI[293] mprj_logic_high_inst/HI[294] mprj_logic_high_inst/HI[295]
+ mprj_logic_high_inst/HI[296] mprj_logic_high_inst/HI[297] mprj_logic_high_inst/HI[298]
+ mprj_logic_high_inst/HI[299] mprj_adr_buf\[19\]/TE mprj_clk2_buf/TE mprj_logic_high_inst/HI[300]
+ mprj_logic_high_inst/HI[301] mprj_logic_high_inst/HI[302] mprj_logic_high_inst/HI[303]
+ mprj_logic_high_inst/HI[304] mprj_logic_high_inst/HI[305] mprj_logic_high_inst/HI[306]
+ mprj_logic_high_inst/HI[307] mprj_logic_high_inst/HI[308] mprj_logic_high_inst/HI[309]
+ mprj_adr_buf\[20\]/TE mprj_logic_high_inst/HI[310] mprj_logic_high_inst/HI[311]
+ mprj_logic_high_inst/HI[312] mprj_logic_high_inst/HI[313] mprj_logic_high_inst/HI[314]
+ mprj_logic_high_inst/HI[315] mprj_logic_high_inst/HI[316] mprj_logic_high_inst/HI[317]
+ mprj_logic_high_inst/HI[318] mprj_logic_high_inst/HI[319] mprj_adr_buf\[21\]/TE
+ mprj_logic_high_inst/HI[320] mprj_logic_high_inst/HI[321] mprj_logic_high_inst/HI[322]
+ mprj_logic_high_inst/HI[323] mprj_logic_high_inst/HI[324] mprj_logic_high_inst/HI[325]
+ mprj_logic_high_inst/HI[326] mprj_logic_high_inst/HI[327] mprj_logic_high_inst/HI[328]
+ mprj_logic_high_inst/HI[329] mprj_adr_buf\[22\]/TE mprj_logic_high_inst/HI[330]
+ mprj_logic_high_inst/HI[331] mprj_logic_high_inst/HI[332] mprj_logic_high_inst/HI[333]
+ mprj_logic_high_inst/HI[334] mprj_logic_high_inst/HI[335] mprj_logic_high_inst/HI[336]
+ mprj_logic_high_inst/HI[337] mprj_logic_high_inst/HI[338] mprj_logic_high_inst/HI[339]
+ mprj_adr_buf\[23\]/TE mprj_logic_high_inst/HI[340] mprj_logic_high_inst/HI[341]
+ mprj_logic_high_inst/HI[342] mprj_logic_high_inst/HI[343] mprj_logic_high_inst/HI[344]
+ mprj_logic_high_inst/HI[345] mprj_logic_high_inst/HI[346] mprj_logic_high_inst/HI[347]
+ mprj_logic_high_inst/HI[348] mprj_logic_high_inst/HI[349] mprj_adr_buf\[24\]/TE
+ mprj_logic_high_inst/HI[350] mprj_logic_high_inst/HI[351] mprj_logic_high_inst/HI[352]
+ mprj_logic_high_inst/HI[353] mprj_logic_high_inst/HI[354] mprj_logic_high_inst/HI[355]
+ mprj_logic_high_inst/HI[356] mprj_logic_high_inst/HI[357] mprj_logic_high_inst/HI[358]
+ mprj_logic_high_inst/HI[359] mprj_adr_buf\[25\]/TE mprj_logic_high_inst/HI[360]
+ mprj_logic_high_inst/HI[361] mprj_logic_high_inst/HI[362] mprj_logic_high_inst/HI[363]
+ mprj_logic_high_inst/HI[364] mprj_logic_high_inst/HI[365] mprj_logic_high_inst/HI[366]
+ mprj_logic_high_inst/HI[367] mprj_logic_high_inst/HI[368] mprj_logic_high_inst/HI[369]
+ mprj_adr_buf\[26\]/TE mprj_logic_high_inst/HI[370] mprj_logic_high_inst/HI[371]
+ mprj_logic_high_inst/HI[372] mprj_logic_high_inst/HI[373] mprj_logic_high_inst/HI[374]
+ mprj_logic_high_inst/HI[375] mprj_logic_high_inst/HI[376] mprj_logic_high_inst/HI[377]
+ mprj_logic_high_inst/HI[378] mprj_logic_high_inst/HI[379] mprj_adr_buf\[27\]/TE
+ mprj_logic_high_inst/HI[380] mprj_logic_high_inst/HI[381] mprj_logic_high_inst/HI[382]
+ mprj_logic_high_inst/HI[383] mprj_logic_high_inst/HI[384] mprj_logic_high_inst/HI[385]
+ mprj_logic_high_inst/HI[386] mprj_logic_high_inst/HI[387] mprj_logic_high_inst/HI[388]
+ mprj_logic_high_inst/HI[389] mprj_adr_buf\[28\]/TE mprj_logic_high_inst/HI[390]
+ mprj_logic_high_inst/HI[391] mprj_logic_high_inst/HI[392] mprj_logic_high_inst/HI[393]
+ mprj_logic_high_inst/HI[394] mprj_logic_high_inst/HI[395] mprj_logic_high_inst/HI[396]
+ mprj_logic_high_inst/HI[397] mprj_logic_high_inst/HI[398] mprj_logic_high_inst/HI[399]
+ mprj_adr_buf\[29\]/TE mprj_cyc_buf/TE mprj_logic_high_inst/HI[400] mprj_logic_high_inst/HI[401]
+ mprj_logic_high_inst/HI[402] mprj_logic_high_inst/HI[403] mprj_logic_high_inst/HI[404]
+ mprj_logic_high_inst/HI[405] mprj_logic_high_inst/HI[406] mprj_logic_high_inst/HI[407]
+ mprj_logic_high_inst/HI[408] mprj_logic_high_inst/HI[409] mprj_adr_buf\[30\]/TE
+ mprj_logic_high_inst/HI[410] mprj_logic_high_inst/HI[411] mprj_logic_high_inst/HI[412]
+ mprj_logic_high_inst/HI[413] mprj_logic_high_inst/HI[414] mprj_logic_high_inst/HI[415]
+ mprj_logic_high_inst/HI[416] mprj_logic_high_inst/HI[417] mprj_logic_high_inst/HI[418]
+ mprj_logic_high_inst/HI[419] mprj_adr_buf\[31\]/TE mprj_logic_high_inst/HI[420]
+ mprj_logic_high_inst/HI[421] mprj_logic_high_inst/HI[422] mprj_logic_high_inst/HI[423]
+ mprj_logic_high_inst/HI[424] mprj_logic_high_inst/HI[425] mprj_logic_high_inst/HI[426]
+ mprj_logic_high_inst/HI[427] mprj_logic_high_inst/HI[428] mprj_logic_high_inst/HI[429]
+ mprj_dat_buf\[0\]/TE mprj_logic_high_inst/HI[430] mprj_logic_high_inst/HI[431] mprj_logic_high_inst/HI[432]
+ mprj_logic_high_inst/HI[433] mprj_logic_high_inst/HI[434] mprj_logic_high_inst/HI[435]
+ mprj_logic_high_inst/HI[436] mprj_logic_high_inst/HI[437] mprj_logic_high_inst/HI[438]
+ mprj_logic_high_inst/HI[439] mprj_dat_buf\[1\]/TE mprj_logic_high_inst/HI[440] mprj_logic_high_inst/HI[441]
+ mprj_logic_high_inst/HI[442] mprj_logic_high_inst/HI[443] mprj_logic_high_inst/HI[444]
+ mprj_logic_high_inst/HI[445] mprj_logic_high_inst/HI[446] mprj_logic_high_inst/HI[447]
+ mprj_logic_high_inst/HI[448] mprj_logic_high_inst/HI[449] mprj_dat_buf\[2\]/TE mprj_logic_high_inst/HI[450]
+ mprj_logic_high_inst/HI[451] mprj_logic_high_inst/HI[452] mprj_logic_high_inst/HI[453]
+ mprj_logic_high_inst/HI[454] mprj_logic_high_inst/HI[455] mprj_logic_high_inst/HI[456]
+ mprj_logic_high_inst/HI[457] user_irq_ena_buf\[0\]/B user_irq_ena_buf\[1\]/B mprj_dat_buf\[3\]/TE
+ user_irq_ena_buf\[2\]/B mprj_pwrgood/A user_to_mprj_wb_ena_buf/B mprj_dat_buf\[4\]/TE
+ mprj_dat_buf\[5\]/TE mprj_dat_buf\[6\]/TE mprj_dat_buf\[7\]/TE mprj_stb_buf/TE mprj_dat_buf\[8\]/TE
+ mprj_dat_buf\[9\]/TE mprj_dat_buf\[10\]/TE mprj_dat_buf\[11\]/TE mprj_dat_buf\[12\]/TE
+ mprj_dat_buf\[13\]/TE mprj_dat_buf\[14\]/TE mprj_dat_buf\[15\]/TE mprj_dat_buf\[16\]/TE
+ mprj_dat_buf\[17\]/TE mprj_we_buf/TE mprj_dat_buf\[18\]/TE mprj_dat_buf\[19\]/TE
+ mprj_dat_buf\[20\]/TE mprj_dat_buf\[21\]/TE mprj_dat_buf\[22\]/TE mprj_dat_buf\[23\]/TE
+ mprj_dat_buf\[24\]/TE mprj_dat_buf\[25\]/TE mprj_dat_buf\[26\]/TE mprj_dat_buf\[27\]/TE
+ mprj_sel_buf\[0\]/TE mprj_dat_buf\[28\]/TE mprj_dat_buf\[29\]/TE mprj_dat_buf\[30\]/TE
+ mprj_dat_buf\[31\]/TE la_buf_enable\[0\]/B la_buf_enable\[1\]/B la_buf_enable\[2\]/B
+ la_buf_enable\[3\]/B la_buf_enable\[4\]/B la_buf_enable\[5\]/B mprj_sel_buf\[1\]/TE
+ la_buf_enable\[6\]/B la_buf_enable\[7\]/B la_buf_enable\[8\]/B la_buf_enable\[9\]/B
+ la_buf_enable\[10\]/B la_buf_enable\[11\]/B la_buf_enable\[12\]/B la_buf_enable\[13\]/B
+ la_buf_enable\[14\]/B la_buf_enable\[15\]/B mprj_sel_buf\[2\]/TE la_buf_enable\[16\]/B
+ la_buf_enable\[17\]/B la_buf_enable\[18\]/B la_buf_enable\[19\]/B la_buf_enable\[20\]/B
+ la_buf_enable\[21\]/B la_buf_enable\[22\]/B la_buf_enable\[23\]/B la_buf_enable\[24\]/B
+ la_buf_enable\[25\]/B mprj_sel_buf\[3\]/TE vccd1_uq5 vssd1_uq4 mprj_logic_high
XFILLER_26_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__376__A _376_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_A input127/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input163_A la_data_out_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[118\]_B la_buf_enable\[118\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[20\]_A input44/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput211 la_data_out_mprj[56] vssd vssd vccd vccd _520_/A sky130_fd_sc_hd__clkbuf_2
Xinput200 la_data_out_mprj[46] vssd vssd vccd vccd _510_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input330_A la_iena_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input428_A la_oenb_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput222 la_data_out_mprj[66] vssd vssd vccd vccd _530_/A sky130_fd_sc_hd__clkbuf_2
Xinput233 la_data_out_mprj[76] vssd vssd vccd vccd _540_/A sky130_fd_sc_hd__clkbuf_4
Xinput244 la_data_out_mprj[86] vssd vssd vccd vccd _550_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input24_A la_data_out_core[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput255 la_data_out_mprj[96] vssd vssd vccd vccd _560_/A sky130_fd_sc_hd__buf_2
Xinput266 la_iena_mprj[105] vssd vssd vccd vccd input266/X sky130_fd_sc_hd__clkbuf_1
Xinput277 la_iena_mprj[115] vssd vssd vccd vccd input277/X sky130_fd_sc_hd__clkbuf_1
Xinput288 la_iena_mprj[125] vssd vssd vccd vccd input288/X sky130_fd_sc_hd__clkbuf_1
X_654_ _654_/A vssd vssd vccd vccd _654_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput299 la_iena_mprj[1] vssd vssd vccd vccd input299/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_1004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[72\] _536_/Y la_buf\[72\]/TE vssd vssd vccd vccd output724/A sky130_fd_sc_hd__einvp_8
X_585_ _585_/A vssd vssd vccd vccd _585_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_wb_dat_buffers\[9\]_A user_wb_dat_gates\[9\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[87\]_A input117/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput718 output718/A vssd vssd vccd vccd la_data_in_core[67] sky130_fd_sc_hd__buf_2
Xoutput707 output707/A vssd vssd vccd vccd la_data_in_core[57] sky130_fd_sc_hd__buf_2
Xoutput729 output729/A vssd vssd vccd vccd la_data_in_core[77] sky130_fd_sc_hd__buf_2
XANTENNA_output647_A output647/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[109\]_B la_buf_enable\[109\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[11\]_A input26/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output814_A output814/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[61\] input89/X user_to_mprj_in_gates\[61\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[61\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[78\]_A input107/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[6\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[26\]_TE la_buf\[26\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[0\]_A_N _592_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output1009_A output1009/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[6\]_B user_to_mprj_in_gates\[6\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_564 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_370_ _370_/A vssd vssd vccd vccd _370_/Y sky130_fd_sc_hd__inv_2
XTAP_1969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[69\]_A input97/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input280_A la_iena_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input378_A la_iena_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input545_A mprj_adr_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_637_ _637_/A vssd vssd vccd vccd _637_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_568_ _568_/A vssd vssd vccd vccd _568_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[49\]_TE la_buf\[49\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_499_ _499_/A vssd vssd vccd vccd _499_/Y sky130_fd_sc_hd__clkinv_2
Xuser_to_mprj_in_buffers\[31\] user_to_mprj_in_gates\[31\]/Y vssd vssd vccd vccd output807/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_34_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output764_A output764/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output931_A output931/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1056 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__654__A _654_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[71\] input356/X mprj_logic_high_inst/HI[401] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[71\]/B sky130_fd_sc_hd__and2_1
XFILLER_49_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input126_A la_data_out_core[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_422_ _422_/A vssd vssd vccd vccd _422_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_14_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[126\]_A input33/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__564__A _564_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_353_ _353_/A vssd vssd vccd vccd _353_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input495_A la_oenb_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input91_A la_data_out_core[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[35\] _499_/Y la_buf\[35\]/TE vssd vssd vccd vccd output683/A sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[107\] input268/X mprj_logic_high_inst/HI[437] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[107\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_gates\[7\] input579/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[7\]/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_10_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput8 la_data_out_core[103] vssd vssd vccd vccd input8/X sky130_fd_sc_hd__buf_4
XFILLER_42_1447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[79\] user_to_mprj_in_gates\[79\]/Y vssd vssd vccd vccd output859/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf_enable\[60\]_A_N _652_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output979_A output979/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__474__A _474_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output881_A output881/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[117\]_A input23/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[24\] input48/X user_to_mprj_in_gates\[24\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[24\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA_la_buf_enable\[75\]_A_N _338_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_560 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[13\]_A_N _605_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__649__A _649_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[28\]_A_N _620_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__384__A _384_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[108\]_A input13/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output1076_A output1076/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[75\] _338_/Y mprj_logic_high_inst/HI[277] vssd vssd vccd
+ vccd output983/A sky130_fd_sc_hd__einvp_4
XFILLER_3_747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput890 output890/A vssd vssd vccd vccd la_oenb_core[106] sky130_fd_sc_hd__buf_2
Xla_buf_enable\[97\] _360_/A la_buf_enable\[97\]/B vssd vssd vccd vccd la_buf\[97\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_dat_buf\[23\] _455_/Y mprj_dat_buf\[23\]/TE vssd vssd vccd vccd output1092/A
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input243_A la_data_out_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__559__A _559_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input410_A la_oenb_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input508_A la_oenb_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_405_ _405_/A vssd vssd vccd vccd _405_/Y sky130_fd_sc_hd__inv_12
XPHY_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_336_ _336_/A vssd vssd vccd vccd _336_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput1006 output1006/A vssd vssd vccd vccd la_oenb_core[96] sky130_fd_sc_hd__buf_2
XFILLER_48_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput1028 output1028/A vssd vssd vccd vccd mprj_adr_o_user[24] sky130_fd_sc_hd__buf_2
Xoutput1017 output1017/A vssd vssd vccd vccd mprj_adr_o_user[14] sky130_fd_sc_hd__buf_2
Xoutput1039 output1039/A vssd vssd vccd vccd mprj_adr_o_user[5] sky130_fd_sc_hd__buf_2
XFILLER_48_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output727_A output727/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__469__A _469_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[122\]_TE mprj_logic_high_inst/HI[324] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[70\]_A input355/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[6\]_B la_buf_enable\[6\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[3\] _595_/A la_buf_enable\[3\]/B vssd vssd vccd vccd la_buf\[3\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_21_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput607 mprj_dat_o_core[3] vssd vssd vccd vccd _435_/A sky130_fd_sc_hd__clkbuf_2
Xinput618 mprj_sel_o_core[3] vssd vssd vccd vccd _399_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__379__A _379_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[21\]_TE mprj_logic_high_inst/HI[223] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[34\] input315/X mprj_logic_high_inst/HI[364] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[34\]/B sky130_fd_sc_hd__and2_1
XFILLER_3_1282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[61\]_A input345/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[12\] _604_/A la_buf_enable\[12\]/B vssd vssd vccd vccd la_buf\[12\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_input193_A la_data_out_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input360_A la_iena_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input458_A la_oenb_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input54_A la_data_out_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input625_A user_irq_ena[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xpowergood_check mprj2_vdd_pwrgood/A mprj_vdd_pwrgood/A vccd vssd vccd vssd vccd vssd
+ mgmt_protect_hv
XFILLER_4_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_80 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[52\]_A input335/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output677_A output677/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput22 la_data_out_core[116] vssd vssd vccd vccd input22/X sky130_fd_sc_hd__clkbuf_4
Xinput11 la_data_out_core[106] vssd vssd vccd vccd input11/X sky130_fd_sc_hd__buf_4
Xinput33 la_data_out_core[126] vssd vssd vccd vccd input33/X sky130_fd_sc_hd__clkbuf_4
Xinput55 la_data_out_core[30] vssd vssd vccd vccd input55/X sky130_fd_sc_hd__clkbuf_4
Xinput44 la_data_out_core[20] vssd vssd vccd vccd input44/X sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput88 la_data_out_core[60] vssd vssd vccd vccd input88/X sky130_fd_sc_hd__buf_4
Xinput77 la_data_out_core[50] vssd vssd vccd vccd input77/X sky130_fd_sc_hd__buf_4
Xinput66 la_data_out_core[40] vssd vssd vccd vccd input66/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_output844_A output844/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput99 la_data_out_core[70] vssd vssd vccd vccd input99/X sky130_fd_sc_hd__buf_4
XFILLER_6_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[91\] input122/X user_to_mprj_in_gates\[91\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[91\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_48_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[44\]_TE mprj_logic_high_inst/HI[246] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[0\]_A _396_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[43\]_A input325/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_49 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_319 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output1039_A output1039/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput426 la_oenb_mprj[19] vssd vssd vccd vccd _611_/A sky130_fd_sc_hd__clkbuf_4
Xinput437 la_oenb_mprj[29] vssd vssd vccd vccd _621_/A sky130_fd_sc_hd__buf_2
Xinput404 la_oenb_mprj[114] vssd vssd vccd vccd _377_/A sky130_fd_sc_hd__clkbuf_4
Xinput415 la_oenb_mprj[124] vssd vssd vccd vccd _387_/A sky130_fd_sc_hd__clkbuf_4
Xuser_to_mprj_oen_buffers\[108\] _371_/Y mprj_logic_high_inst/HI[310] vssd vssd vccd
+ vccd output892/A sky130_fd_sc_hd__einvp_4
Xinput459 la_oenb_mprj[49] vssd vssd vccd vccd _641_/A sky130_fd_sc_hd__buf_2
Xinput448 la_oenb_mprj[39] vssd vssd vccd vccd _631_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[38\] _630_/Y mprj_logic_high_inst/HI[240] vssd vssd vccd
+ vccd output942/A sky130_fd_sc_hd__einvp_4
XFILLER_44_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[34\]_A input315/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input206_A la_data_out_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__572__A _572_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input575_A mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[82\]_TE la_buf\[82\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[1\]_A _433_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[67\]_TE mprj_logic_high_inst/HI[269] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[61\] user_to_mprj_in_gates\[61\]/Y vssd vssd vccd vccd output840/A
+ sky130_fd_sc_hd__inv_2
XFILLER_34_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[25\]_A input305/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output794_A output794/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output961_A output961/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__482__A _482_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[31\]_TE mprj_dat_buf\[31\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[90\]_A user_to_mprj_in_gates\[90\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__657__A _657_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[16\]_A input295/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_B user_to_mprj_in_gates\[96\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__392__A _392_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1850 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[20\]_B user_to_mprj_in_gates\[20\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xinput201 la_data_out_mprj[47] vssd vssd vccd vccd _511_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_buffers\[81\]_A user_to_mprj_in_gates\[81\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_input156_A la_data_out_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput212 la_data_out_mprj[57] vssd vssd vccd vccd _521_/A sky130_fd_sc_hd__clkbuf_2
Xinput223 la_data_out_mprj[67] vssd vssd vccd vccd _531_/A sky130_fd_sc_hd__clkbuf_2
Xinput234 la_data_out_mprj[77] vssd vssd vccd vccd _541_/A sky130_fd_sc_hd__buf_2
Xinput245 la_data_out_mprj[87] vssd vssd vccd vccd _551_/A sky130_fd_sc_hd__buf_2
XANTENNA_input323_A la_iena_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput256 la_data_out_mprj[97] vssd vssd vccd vccd _561_/A sky130_fd_sc_hd__buf_2
Xinput267 la_iena_mprj[106] vssd vssd vccd vccd input267/X sky130_fd_sc_hd__clkbuf_1
Xinput278 la_iena_mprj[116] vssd vssd vccd vccd input278/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input17_A la_data_out_core[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__567__A _567_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_653_ _653_/A vssd vssd vccd vccd _653_/Y sky130_fd_sc_hd__inv_2
Xinput289 la_iena_mprj[126] vssd vssd vccd vccd input289/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[65\] _529_/Y la_buf\[65\]/TE vssd vssd vccd vccd output716/A sky130_fd_sc_hd__einvp_8
XFILLER_38_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_584_ _584_/A vssd vssd vccd vccd _584_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_44_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[87\]_B user_to_mprj_in_gates\[87\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput708 output708/A vssd vssd vccd vccd la_data_in_core[58] sky130_fd_sc_hd__buf_2
Xla_buf\[121\] _585_/Y la_buf\[121\]/TE vssd vssd vccd vccd output651/A sky130_fd_sc_hd__einvp_4
Xmprj_adr_buf\[29\] _429_/Y mprj_adr_buf\[29\]/TE vssd vssd vccd vccd output1033/A
+ sky130_fd_sc_hd__einvp_8
Xoutput719 output719/A vssd vssd vccd vccd la_data_in_core[68] sky130_fd_sc_hd__buf_2
XFILLER_49_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[11\]_B user_to_mprj_in_gates\[11\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[72\]_A user_to_mprj_in_gates\[72\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output807_A output807/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__477__A _477_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[54\] input81/X user_to_mprj_in_gates\[54\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[54\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[78\]_B user_to_mprj_in_gates\[78\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[110\]_A user_to_mprj_in_gates\[110\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[63\]_A user_to_mprj_in_gates\[63\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_input9_A la_data_out_core[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__387__A _387_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[69\]_B user_to_mprj_in_gates\[69\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input273_A la_iena_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[101\]_A user_to_mprj_in_gates\[101\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input440_A la_oenb_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input538_A mprj_adr_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[54\]_A user_to_mprj_in_gates\[54\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[101\]_A_N _364_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_636_ _636_/A vssd vssd vccd vccd _636_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[116\]_A_N _379_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_567_ _567_/A vssd vssd vccd vccd _567_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[22\]_TE mprj_adr_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_498_ _498_/A vssd vssd vccd vccd _498_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf\[94\]_A _558_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[24\] user_to_mprj_in_gates\[24\]/Y vssd vssd vccd vccd output799/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output757_A output757/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output924_A output924/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[45\]_A user_to_mprj_in_gates\[45\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_354 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[85\]_A _549_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1021_A output1021/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1119_A output1119/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[36\]_A user_to_mprj_in_gates\[36\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[64\] input348/X mprj_logic_high_inst/HI[394] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[64\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input119_A la_data_out_core[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[20\] _612_/Y mprj_logic_high_inst/HI[222] vssd vssd vccd
+ vccd output923/A sky130_fd_sc_hd__einvp_2
XFILLER_42_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[42\] _634_/A la_buf_enable\[42\]/B vssd vssd vccd vccd la_buf\[42\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[2\] _594_/Y mprj_logic_high_inst/HI[204] vssd vssd vccd
+ vccd output933/A sky130_fd_sc_hd__einvp_4
X_421_ _421_/A vssd vssd vccd vccd _421_/Y sky130_fd_sc_hd__inv_12
XTAP_1756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[126\]_B user_to_mprj_in_gates\[126\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_352_ _352_/A vssd vssd vccd vccd _352_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[76\]_A _540_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input390_A la_oenb_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input84_A la_data_out_core[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[94\]_B la_buf_enable\[94\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input488_A la_oenb_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__580__A _580_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[28\] _492_/Y la_buf\[28\]/TE vssd vssd vccd vccd output675/A sky130_fd_sc_hd__einvp_8
XFILLER_6_745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[27\]_A user_to_mprj_in_gates\[27\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput9 la_data_out_core[104] vssd vssd vccd vccd input9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[16\]_TE la_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_619_ _619_/A vssd vssd vccd vccd _619_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[67\]_A _531_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output874_A output874/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[117\]_B user_to_mprj_in_gates\[117\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[17\] input40/X user_to_mprj_in_gates\[17\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[17\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[85\]_B la_buf_enable\[85\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__490__A _490_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[27\] user_wb_dat_gates\[27\]/Y vssd vssd vccd vccd output1064/A
+ sky130_fd_sc_hd__inv_6
XFILLER_25_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[18\]_A user_to_mprj_in_gates\[18\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[26\]_A input568/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[58\]_A _522_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[108\]_B user_to_mprj_in_gates\[108\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_51_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_15 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_48 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[76\]_B la_buf_enable\[76\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output1069_A output1069/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1352 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput891 output891/A vssd vssd vccd vccd la_oenb_core[107] sky130_fd_sc_hd__buf_2
XFILLER_2_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput880 output880/A vssd vssd vccd vccd la_data_in_mprj[98] sky130_fd_sc_hd__buf_2
XFILLER_43_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[68\] _331_/Y mprj_logic_high_inst/HI[270] vssd vssd vccd
+ vccd output975/A sky130_fd_sc_hd__einvp_8
XANTENNA_user_wb_dat_gates\[17\]_A input558/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[16\] _448_/Y mprj_dat_buf\[16\]/TE vssd vssd vccd vccd output1084/A
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input236_A la_data_out_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[39\]_TE la_buf\[39\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input403_A la_oenb_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__575__A _575_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[49\]_A _513_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_404_ _404_/A vssd vssd vccd vccd _404_/Y sky130_fd_sc_hd__inv_2
XTAP_1597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_335_ _335_/A vssd vssd vccd vccd _335_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[67\]_B la_buf_enable\[67\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput1007 output1007/A vssd vssd vccd vccd la_oenb_core[97] sky130_fd_sc_hd__buf_2
Xoutput1029 output1029/A vssd vssd vccd vccd mprj_adr_o_user[25] sky130_fd_sc_hd__buf_2
Xoutput1018 output1018/A vssd vssd vccd vccd mprj_adr_o_user[15] sky130_fd_sc_hd__buf_2
XFILLER_29_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_adr_buf\[11\] _411_/Y mprj_adr_buf\[11\]/TE vssd vssd vccd vccd output1014/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_26_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[125\] user_to_mprj_in_gates\[125\]/Y vssd vssd vccd vccd
+ output783/A sky130_fd_sc_hd__clkinv_4
XFILLER_2_781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_20 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[91\] user_to_mprj_in_gates\[91\]/Y vssd vssd vccd vccd output873/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_49_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output991_A output991/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__485__A _485_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[1\] user_wb_dat_gates\[1\]/Y vssd vssd vccd vccd output1056/A
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_user_to_mprj_in_ena_buf\[70\]_B mprj_logic_high_inst/HI[400] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[7\]_TE la_buf\[7\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[58\]_B la_buf_enable\[58\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[60\]_A _652_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[125\]_A _388_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput619 mprj_stb_o_core vssd vssd vccd vccd _394_/A sky130_fd_sc_hd__clkbuf_4
Xinput608 mprj_dat_o_core[4] vssd vssd vccd vccd _436_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__395__A _395_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[27\] input307/X mprj_logic_high_inst/HI[357] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[27\]/B sky130_fd_sc_hd__and2_1
XFILLER_3_1294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[61\]_B mprj_logic_high_inst/HI[391] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_24_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[49\]_B la_buf_enable\[49\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[116\]_A _379_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[51\]_A _643_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input186_A la_data_out_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input353_A la_iena_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input47_A la_data_out_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input520_A mprj_adr_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[110\] _373_/A la_buf_enable\[110\]/B vssd vssd vccd vccd la_buf\[110\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf_enable\[74\]_A_N _337_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[95\] _559_/Y la_buf\[95\]/TE vssd vssd vccd vccd output749/A sky130_fd_sc_hd__einvp_4
Xuser_to_mprj_in_ena_buf\[0\] input260/X mprj_logic_high_inst/HI[330] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[0\]/B sky130_fd_sc_hd__and2_1
XFILLER_4_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input618_A mprj_sel_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[89\]_A_N _352_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[52\]_B mprj_logic_high_inst/HI[382] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_15_652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[12\]_A_N _604_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput12 la_data_out_core[107] vssd vssd vccd vccd input12/X sky130_fd_sc_hd__buf_4
XFILLER_52_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput34 la_data_out_core[127] vssd vssd vccd vccd input34/X sky130_fd_sc_hd__clkbuf_4
Xinput23 la_data_out_core[117] vssd vssd vccd vccd input23/X sky130_fd_sc_hd__buf_4
Xinput45 la_data_out_core[21] vssd vssd vccd vccd input45/X sky130_fd_sc_hd__clkbuf_4
XFILLER_15_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[9\]_A input387/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput89 la_data_out_core[61] vssd vssd vccd vccd input89/X sky130_fd_sc_hd__buf_4
Xinput78 la_data_out_core[51] vssd vssd vccd vccd input78/X sky130_fd_sc_hd__buf_4
Xinput67 la_data_out_core[41] vssd vssd vccd vccd input67/X sky130_fd_sc_hd__clkbuf_4
Xinput56 la_data_out_core[31] vssd vssd vccd vccd input56/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_oen_buffers\[42\]_A _634_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[107\]_A _370_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[27\]_A_N _619_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output837_A output837/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[84\] input114/X user_to_mprj_in_gates\[84\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[84\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_788 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[43\]_B mprj_logic_high_inst/HI[373] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_40_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[33\]_A _625_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput427 la_oenb_mprj[1] vssd vssd vccd vccd _593_/A sky130_fd_sc_hd__clkbuf_2
Xinput405 la_oenb_mprj[115] vssd vssd vccd vccd _378_/A sky130_fd_sc_hd__clkbuf_4
Xinput416 la_oenb_mprj[125] vssd vssd vccd vccd _388_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_output1101_A output1101/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput449 la_oenb_mprj[3] vssd vssd vccd vccd _595_/A sky130_fd_sc_hd__clkbuf_2
Xinput438 la_oenb_mprj[2] vssd vssd vccd vccd _594_/A sky130_fd_sc_hd__buf_2
XFILLER_5_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input101_A la_data_out_core[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[34\]_B mprj_logic_high_inst/HI[364] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_43_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1878 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input470_A la_oenb_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input568_A mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[24\]_A _616_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[6\] _470_/Y la_buf\[6\]/TE vssd vssd vccd vccd output721/A sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[112\]_TE mprj_logic_high_inst/HI[314] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[10\] _474_/Y la_buf\[10\]/TE vssd vssd vccd vccd output638/A sky130_fd_sc_hd__einvp_8
XFILLER_45_2328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[3\] _403_/Y mprj_adr_buf\[3\]/TE vssd vssd vccd vccd output1037/A sky130_fd_sc_hd__einvp_8
XFILLER_47_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_we_buf_TE mprj_we_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[20\]_A _420_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[25\]_B mprj_logic_high_inst/HI[355] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[54\] user_to_mprj_in_gates\[54\]/Y vssd vssd vccd vccd output832/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_37_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output787_A output787/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_gates\[12\] input553/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[12\]/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_50_2067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output954_A output954/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[11\]_TE mprj_logic_high_inst/HI[213] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[15\]_A _607_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[110\] input16/X user_to_mprj_in_gates\[110\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[110\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA_mprj_adr_buf\[11\]_A _411_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[16\]_B mprj_logic_high_inst/HI[346] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_43_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[9\]_A input581/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1051_A output1051/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[94\] input381/X mprj_logic_high_inst/HI[424] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[94\]/B sky130_fd_sc_hd__and2_1
XFILLER_27_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[120\] _383_/Y mprj_logic_high_inst/HI[322] vssd vssd vccd
+ vccd output906/A sky130_fd_sc_hd__einvp_4
XFILLER_44_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_sel_buf\[1\] _397_/Y mprj_sel_buf\[1\]/TE vssd vssd vccd vccd output1110/A sky130_fd_sc_hd__einvp_8
XFILLER_1_857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput202 la_data_out_mprj[48] vssd vssd vccd vccd _512_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput213 la_data_out_mprj[58] vssd vssd vccd vccd _522_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput224 la_data_out_mprj[68] vssd vssd vccd vccd _532_/A sky130_fd_sc_hd__clkbuf_2
Xinput235 la_data_out_mprj[78] vssd vssd vccd vccd _542_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input149_A la_data_out_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[9\]_A input131/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[72\] _335_/A la_buf_enable\[72\]/B vssd vssd vccd vccd la_buf\[72\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[50\] _642_/Y mprj_logic_high_inst/HI[252] vssd vssd vccd
+ vccd output956/A sky130_fd_sc_hd__einvp_4
Xinput246 la_data_out_mprj[88] vssd vssd vccd vccd _552_/A sky130_fd_sc_hd__clkbuf_4
Xinput257 la_data_out_mprj[98] vssd vssd vccd vccd _562_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput268 la_iena_mprj[107] vssd vssd vccd vccd input268/X sky130_fd_sc_hd__clkbuf_1
Xinput279 la_iena_mprj[117] vssd vssd vccd vccd input279/X sky130_fd_sc_hd__clkbuf_1
X_652_ _652_/A vssd vssd vccd vccd _652_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input316_A la_iena_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_583_ _583_/A vssd vssd vccd vccd _583_/Y sky130_fd_sc_hd__inv_2
XANTENNA__583__A _583_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[58\] _522_/Y la_buf\[58\]/TE vssd vssd vccd vccd output708/A sky130_fd_sc_hd__einvp_8
XFILLER_16_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[34\]_TE mprj_logic_high_inst/HI[236] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput709 output709/A vssd vssd vccd vccd la_data_in_core[59] sky130_fd_sc_hd__buf_2
XFILLER_12_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[114\] _578_/Y la_buf\[114\]/TE vssd vssd vccd vccd output643/A sky130_fd_sc_hd__einvp_4
XFILLER_10_1361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output702_A output702/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[47\] input73/X user_to_mprj_in_gates\[47\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[47\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_514 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__493__A _493_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[9\]_TE mprj_adr_buf\[9\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[9\] input131/X user_to_mprj_in_gates\[9\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[9\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_8_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2016 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[72\]_TE la_buf\[72\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1099_A output1099/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[57\]_TE mprj_logic_high_inst/HI[259] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[98\] _361_/Y mprj_logic_high_inst/HI[300] vssd vssd vccd
+ vccd output1008/A sky130_fd_sc_hd__einvp_8
XFILLER_13_1979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input266_A la_iena_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input433_A la_oenb_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__578__A _578_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input600_A mprj_dat_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_82 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_635_ _635_/A vssd vssd vccd vccd _635_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_dat_buf\[24\]_A _456_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_buffers\[31\]_A user_wb_dat_gates\[31\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_44_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_566_ _566_/A vssd vssd vccd vccd _566_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_dat_buf\[21\]_TE mprj_dat_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1824 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_497_ _497_/A vssd vssd vccd vccd _497_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_51_2162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[0\]_TE mprj_logic_high_inst/HI[202] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[17\] user_to_mprj_in_gates\[17\]/Y vssd vssd vccd vccd output791/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output652_A output652/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output917_A output917/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[95\]_TE la_buf\[95\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__488__A _488_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[15\]_A _447_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[22\]_A user_wb_dat_gates\[22\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_36_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output1014_A output1014/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__398__A _398_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[57\] input340/X mprj_logic_high_inst/HI[387] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[57\]/B sky130_fd_sc_hd__and2_1
XTAP_580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_buffers\[13\]_A user_wb_dat_gates\[13\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XTAP_1713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_420_ _420_/A vssd vssd vccd vccd _420_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_14_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[13\] _605_/Y mprj_logic_high_inst/HI[215] vssd vssd vccd
+ vccd output915/A sky130_fd_sc_hd__einvp_2
X_351_ _351_/A vssd vssd vccd vccd _351_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[35\] _627_/A la_buf_enable\[35\]/B vssd vssd vccd vccd la_buf\[35\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_1779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[9\] user_to_mprj_in_gates\[9\]/Y vssd vssd vccd vccd output882/A
+ sky130_fd_sc_hd__inv_6
XANTENNA_input383_A la_iena_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input77_A la_data_out_core[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input550_A mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_618_ _618_/A vssd vssd vccd vccd _618_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_17_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_549_ _549_/A vssd vssd vccd vccd _549_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output867_A output867/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[26\]_B repeater1125/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[100\]_A_N _363_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[12\]_TE mprj_adr_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[115\]_A_N _378_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput870 output870/A vssd vssd vccd vccd la_data_in_mprj[89] sky130_fd_sc_hd__buf_2
Xoutput881 output881/A vssd vssd vccd vccd la_data_in_mprj[99] sky130_fd_sc_hd__buf_2
Xoutput892 output892/A vssd vssd vccd vccd la_oenb_core[108] sky130_fd_sc_hd__buf_2
XFILLER_8_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[17\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input131_A la_data_out_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input229_A la_data_out_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_403_ _403_/A vssd vssd vccd vccd _403_/Y sky130_fd_sc_hd__inv_12
XTAP_1554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[2\]_A _466_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_50 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input598_A mprj_dat_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_334_ _334_/A vssd vssd vccd vccd _334_/Y sky130_fd_sc_hd__inv_2
XTAP_1587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[40\] _504_/Y la_buf\[40\]/TE vssd vssd vccd vccd output689/A sky130_fd_sc_hd__einvp_4
XTAP_1598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__591__A _591_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[112\] input274/X mprj_logic_high_inst/HI[442] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[112\]/B sky130_fd_sc_hd__and2_1
XFILLER_41_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput1008 output1008/A vssd vssd vccd vccd la_oenb_core[98] sky130_fd_sc_hd__buf_2
Xoutput1019 output1019/A vssd vssd vccd vccd mprj_adr_o_user[16] sky130_fd_sc_hd__buf_2
XFILLER_46_2094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_10 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[118\] user_to_mprj_in_gates\[118\]/Y vssd vssd vccd vccd
+ output775/A sky130_fd_sc_hd__clkinv_4
XANTENNA_user_irq_gates\[2\]_A input623/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_43 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[84\] user_to_mprj_in_gates\[84\]/Y vssd vssd vccd vccd output865/A
+ sky130_fd_sc_hd__clkinv_2
XANTENNA_mprj_dat_buf\[0\]_TE mprj_dat_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output984_A output984/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2010 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[120\]_TE la_buf\[120\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput609 mprj_dat_o_core[5] vssd vssd vccd vccd _437_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[9\]_A _409_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output1081_A output1081/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[80\] _343_/Y mprj_logic_high_inst/HI[282] vssd vssd vccd
+ vccd output989/A sky130_fd_sc_hd__einvp_2
XANTENNA_input179_A la_data_out_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[50\]_A input77/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input346_A la_iena_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input513_A la_oenb_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__586__A _586_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[88\] _552_/Y la_buf\[88\]/TE vssd vssd vccd vccd output741/A sky130_fd_sc_hd__einvp_2
XFILLER_21_1831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[103\] _366_/A la_buf_enable\[103\]/B vssd vssd vccd vccd la_buf\[103\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_35_918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[0\]_A user_to_mprj_in_gates\[0\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput13 la_data_out_core[108] vssd vssd vccd vccd input13/X sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_81 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput24 la_data_out_core[118] vssd vssd vccd vccd input24/X sky130_fd_sc_hd__clkbuf_4
Xinput46 la_data_out_core[22] vssd vssd vccd vccd input46/X sky130_fd_sc_hd__clkbuf_4
Xinput35 la_data_out_core[12] vssd vssd vccd vccd input35/X sky130_fd_sc_hd__buf_2
XFILLER_15_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[9\]_B mprj_logic_high_inst/HI[339] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xinput79 la_data_out_core[52] vssd vssd vccd vccd input79/X sky130_fd_sc_hd__buf_4
Xinput68 la_data_out_core[42] vssd vssd vccd vccd input68/X sky130_fd_sc_hd__clkbuf_4
Xinput57 la_data_out_core[32] vssd vssd vccd vccd input57/X sky130_fd_sc_hd__buf_4
XFILLER_48_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output732_A output732/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[41\]_A input67/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[77\] input106/X user_to_mprj_in_gates\[77\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[77\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__496__A _496_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[90\]_TE mprj_logic_high_inst/HI[292] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[29\]_TE la_buf\[29\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[32\]_A input57/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput428 la_oenb_mprj[20] vssd vssd vccd vccd _612_/A sky130_fd_sc_hd__clkbuf_4
Xinput406 la_oenb_mprj[116] vssd vssd vccd vccd _379_/A sky130_fd_sc_hd__clkbuf_4
Xinput417 la_oenb_mprj[126] vssd vssd vccd vccd _389_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput439 la_oenb_mprj[30] vssd vssd vccd vccd _622_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1460 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[99\]_A input130/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_954 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input296_A la_iena_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input463_A la_oenb_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[23\]_A input47/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output682_A output682/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[47\] user_to_mprj_in_gates\[47\]/Y vssd vssd vccd vccd output824/A
+ sky130_fd_sc_hd__inv_2
XFILLER_37_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output947_A output947/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[14\]_A input37/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[103\] input8/X user_to_mprj_in_gates\[103\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[103\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[9\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[73\]_A_N _336_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output1044_A output1044/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[88\]_A_N _351_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[87\] input373/X mprj_logic_high_inst/HI[417] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[87\]/B sky130_fd_sc_hd__and2_1
Xmprj_clk2_buf _392_/Y mprj_clk2_buf/TE vssd vssd vccd vccd output1120/A sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[113\] _376_/Y mprj_logic_high_inst/HI[315] vssd vssd vccd
+ vccd output898/A sky130_fd_sc_hd__einvp_2
Xinput203 la_data_out_mprj[49] vssd vssd vccd vccd _513_/A sky130_fd_sc_hd__clkbuf_2
Xinput214 la_data_out_mprj[59] vssd vssd vccd vccd _523_/A sky130_fd_sc_hd__clkbuf_2
Xinput225 la_data_out_mprj[69] vssd vssd vccd vccd _533_/A sky130_fd_sc_hd__clkbuf_2
Xinput236 la_data_out_mprj[79] vssd vssd vccd vccd _543_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_gates\[9\]_B user_to_mprj_in_gates\[9\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[11\]_A_N _603_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput247 la_data_out_mprj[89] vssd vssd vccd vccd _553_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput258 la_data_out_mprj[99] vssd vssd vccd vccd _563_/A sky130_fd_sc_hd__clkbuf_1
Xinput269 la_iena_mprj[108] vssd vssd vccd vccd input269/X sky130_fd_sc_hd__clkbuf_1
X_651_ _651_/A vssd vssd vccd vccd _651_/Y sky130_fd_sc_hd__clkinv_2
Xuser_to_mprj_oen_buffers\[43\] _635_/Y mprj_logic_high_inst/HI[245] vssd vssd vccd
+ vccd output948/A sky130_fd_sc_hd__einvp_2
Xla_buf_enable\[65\] _657_/A la_buf_enable\[65\]/B vssd vssd vccd vccd la_buf\[65\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_29_564 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_irq_buffers\[1\] user_irq_gates\[1\]/Y vssd vssd vccd vccd output1122/A sky130_fd_sc_hd__clkinv_4
XFILLER_44_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_582_ _582_/A vssd vssd vccd vccd _582_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input211_A la_data_out_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[26\]_A_N _618_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input309_A la_iena_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2344 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input580_A mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[107\] _571_/Y la_buf\[107\]/TE vssd vssd vccd vccd output635/A sky130_fd_sc_hd__einvp_2
XTAP_228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[100\] user_to_mprj_in_gates\[100\]/Y vssd vssd vccd vccd
+ output756/A sky130_fd_sc_hd__inv_2
XFILLER_23_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output897_A output897/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[120\]_A input283/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[102\]_TE mprj_logic_high_inst/HI[304] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[111\]_A input273/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input259_A la_data_out_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input161_A la_data_out_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input426_A la_oenb_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input22_A la_data_out_core[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_634_ _634_/A vssd vssd vccd vccd _634_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_2089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[70\] _534_/Y la_buf\[70\]/TE vssd vssd vccd vccd output722/A sky130_fd_sc_hd__einvp_8
XANTENNA__594__A _594_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_565_ _565_/A vssd vssd vccd vccd _565_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_53_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_496_ _496_/A vssd vssd vccd vccd _496_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[102\]_A input263/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output645_A output645/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output812_A output812/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[125\]_TE mprj_logic_high_inst/HI[327] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[24\]_TE mprj_logic_high_inst/HI[226] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output1007_A output1007/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[91\]_A input378/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ _350_/A vssd vssd vccd vccd _350_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[28\] _620_/A la_buf_enable\[28\]/B vssd vssd vccd vccd la_buf\[28\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_52_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input376_A la_iena_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input543_A mprj_adr_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__589__A _589_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[82\]_A input368/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_617_ _617_/A vssd vssd vccd vccd _617_/Y sky130_fd_sc_hd__clkinv_2
X_548_ _548_/A vssd vssd vccd vccd _548_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_479_ _479_/A vssd vssd vccd vccd _479_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_20_518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output762_A output762/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[62\]_TE la_buf\[62\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[47\]_TE mprj_logic_high_inst/HI[249] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__499__A _499_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[73\]_A input358/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[9\]_B la_buf_enable\[9\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1124_A output1124/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput882 output882/A vssd vssd vccd vccd la_data_in_mprj[9] sky130_fd_sc_hd__buf_2
Xoutput860 output860/A vssd vssd vccd vccd la_data_in_mprj[7] sky130_fd_sc_hd__buf_2
Xoutput871 output871/A vssd vssd vccd vccd la_data_in_mprj[8] sky130_fd_sc_hd__buf_2
Xoutput893 output893/A vssd vssd vccd vccd la_oenb_core[109] sky130_fd_sc_hd__buf_2
XFILLER_47_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[11\]_TE mprj_dat_buf\[11\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input124_A la_data_out_core[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[64\]_A input348/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_402_ _402_/A vssd vssd vccd vccd _402_/Y sky130_fd_sc_hd__inv_2
XPHY_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_333_ _333_/A vssd vssd vccd vccd _333_/Y sky130_fd_sc_hd__inv_2
XTAP_1599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input493_A la_oenb_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[85\]_TE la_buf\[85\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[33\] _497_/Y la_buf\[33\]/TE vssd vssd vccd vccd output681/A sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[105\] input266/X mprj_logic_high_inst/HI[435] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[105\]/B sky130_fd_sc_hd__and2_1
Xuser_wb_dat_gates\[5\] input577/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[5\]/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_48_2305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput1009 output1009/A vssd vssd vccd vccd la_oenb_core[99] sky130_fd_sc_hd__buf_2
XFILLER_29_1025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_irq_gates\[2\]_B user_irq_gates\[2\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[77\] user_to_mprj_in_gates\[77\]/Y vssd vssd vccd vccd output857/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_in_ena_buf\[55\]_A input338/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output977_A output977/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[22\] input46/X user_to_mprj_in_gates\[22\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[22\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_sel_buf\[3\]_A _399_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[46\]_A input328/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output1074_A output1074/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[50\]_B user_to_mprj_in_gates\[50\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xoutput690 output690/A vssd vssd vccd vccd la_data_in_core[41] sky130_fd_sc_hd__buf_2
Xuser_to_mprj_oen_buffers\[73\] _336_/Y mprj_logic_high_inst/HI[275] vssd vssd vccd
+ vccd output981/A sky130_fd_sc_hd__einvp_4
Xla_buf_enable\[95\] _358_/A la_buf_enable\[95\]/B vssd vssd vccd vccd la_buf\[95\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_47_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[21\] _453_/Y mprj_dat_buf\[21\]/TE vssd vssd vccd vccd output1090/A
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input339_A la_iena_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input241_A la_data_out_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input506_A la_oenb_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[37\]_A input318/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_dat_buf\[4\]_A _436_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput25 la_data_out_core[119] vssd vssd vccd vccd input25/X sky130_fd_sc_hd__buf_2
Xinput14 la_data_out_core[109] vssd vssd vccd vccd input14/X sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput36 la_data_out_core[13] vssd vssd vccd vccd input36/X sky130_fd_sc_hd__clkbuf_4
XFILLER_35_1095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput69 la_data_out_core[43] vssd vssd vccd vccd input69/X sky130_fd_sc_hd__clkbuf_4
Xinput58 la_data_out_core[33] vssd vssd vccd vccd input58/X sky130_fd_sc_hd__buf_4
Xinput47 la_data_out_core[23] vssd vssd vccd vccd input47/X sky130_fd_sc_hd__clkbuf_4
XFILLER_32_1972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[41\]_B user_to_mprj_in_gates\[41\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output725_A output725/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[28\]_A input308/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[114\]_A_N _377_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[1\] _593_/A la_buf_enable\[1\]/B vssd vssd vccd vccd la_buf\[1\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_31_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[93\]_A user_to_mprj_in_gates\[93\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[32\]_B user_to_mprj_in_gates\[32\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput407 la_oenb_mprj[117] vssd vssd vccd vccd _380_/A sky130_fd_sc_hd__clkbuf_4
Xinput418 la_oenb_mprj[127] vssd vssd vccd vccd _390_/A sky130_fd_sc_hd__buf_2
XFILLER_5_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput429 la_oenb_mprj[21] vssd vssd vccd vccd _613_/A sky130_fd_sc_hd__buf_2
XFILLER_9_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[19\]_A input298/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[32\] input313/X mprj_logic_high_inst/HI[362] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[32\]/B sky130_fd_sc_hd__and2_1
XFILLER_43_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[99\]_B user_to_mprj_in_gates\[99\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[10\] _602_/A la_buf_enable\[10\]/B vssd vssd vccd vccd la_buf\[10\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_22_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input191_A la_data_out_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input289_A la_iena_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[120\]_A _584_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[23\]_B user_to_mprj_in_gates\[23\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_input456_A la_oenb_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[84\]_A user_to_mprj_in_gates\[84\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input52_A la_data_out_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input623_A user_irq_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[110\]_TE la_buf\[110\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__597__A _597_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[25\]_TE mprj_adr_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output675_A output675/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_432 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[122\]_A user_to_mprj_in_gates\[122\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[111\]_A _575_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output842_A output842/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[14\]_B user_to_mprj_in_gates\[14\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[75\]_A user_to_mprj_in_gates\[75\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[113\]_A user_to_mprj_in_gates\[113\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[102\]_A _566_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[66\]_A user_to_mprj_in_gates\[66\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1037_A output1037/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput226 la_data_out_mprj[6] vssd vssd vccd vccd _470_/A sky130_fd_sc_hd__clkbuf_2
Xinput215 la_data_out_mprj[5] vssd vssd vccd vccd _469_/A sky130_fd_sc_hd__clkbuf_2
Xinput204 la_data_out_mprj[4] vssd vssd vccd vccd _468_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[106\] _369_/Y mprj_logic_high_inst/HI[308] vssd vssd vccd
+ vccd output890/A sky130_fd_sc_hd__einvp_4
Xinput259 la_data_out_mprj[9] vssd vssd vccd vccd _473_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput248 la_data_out_mprj[8] vssd vssd vccd vccd _472_/A sky130_fd_sc_hd__clkbuf_2
Xinput237 la_data_out_mprj[7] vssd vssd vccd vccd _471_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_1100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_650_ _650_/A vssd vssd vccd vccd _650_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_44_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_581_ _581_/A vssd vssd vccd vccd _581_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[58\] _650_/A la_buf_enable\[58\]/B vssd vssd vccd vccd la_buf\[58\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[36\] _628_/Y mprj_logic_high_inst/HI[238] vssd vssd vccd
+ vccd output940/A sky130_fd_sc_hd__einvp_4
XFILLER_22_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input204_A la_data_out_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_73 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input573_A mprj_dat_i_user[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[104\]_A user_to_mprj_in_gates\[104\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[57\]_A user_to_mprj_in_gates\[57\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[30\]_A _494_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[80\]_TE mprj_logic_high_inst/HI[282] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[19\]_TE la_buf\[19\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[97\]_A _561_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output792_A output792/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[120\]_B mprj_logic_high_inst/HI[450] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[48\]_A user_to_mprj_in_gates\[48\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[21\]_A _485_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[88\]_A _552_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[111\]_B mprj_logic_high_inst/HI[441] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1964 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[39\]_A user_to_mprj_in_gates\[39\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[12\]_A _476_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input154_A la_data_out_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[30\]_B la_buf_enable\[30\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input321_A la_iena_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input15_A la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_633_ _633_/A vssd vssd vccd vccd _633_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input419_A la_oenb_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[79\]_A _543_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[63\] _527_/Y la_buf\[63\]/TE vssd vssd vccd vccd output714/A sky130_fd_sc_hd__einvp_8
XFILLER_2_1895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_564_ _564_/A vssd vssd vccd vccd _564_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_38_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_495_ _495_/A vssd vssd vccd vccd _495_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_18_1815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[102\]_B mprj_logic_high_inst/HI[432] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_44_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[97\]_B la_buf_enable\[97\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[27\] _427_/Y mprj_adr_buf\[27\]/TE vssd vssd vccd vccd output1031/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output638_A output638/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_77 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_ack_gate input516/X repeater1125/A vssd vssd vccd vccd user_wb_ack_gate/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_49_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[21\]_B la_buf_enable\[21\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output805_A output805/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[72\]_A_N _335_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[52\] input79/X user_to_mprj_in_gates\[52\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[52\]/Y sky130_fd_sc_hd__nand2_1
Xinput590 mprj_dat_o_core[17] vssd vssd vccd vccd _449_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[87\]_A_N _350_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[88\]_B la_buf_enable\[88\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[10\]_A_N _602_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[90\]_A _353_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[25\]_A_N _617_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[29\]_A input571/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input7_A la_data_out_core[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[12\]_B la_buf_enable\[12\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[91\]_B mprj_logic_high_inst/HI[421] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_1715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[79\]_B la_buf_enable\[79\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[81\]_A _344_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input271_A la_iena_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input369_A la_iena_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input536_A mprj_adr_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[126\] _389_/A la_buf_enable\[126\]/B vssd vssd vccd vccd la_buf\[126\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_4_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[82\]_B mprj_logic_high_inst/HI[412] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_616_ _616_/A vssd vssd vccd vccd _616_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_17_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_547_ _547_/A vssd vssd vccd vccd _547_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_478_ _478_/A vssd vssd vccd vccd _478_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[72\]_A _335_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[22\] user_to_mprj_in_gates\[22\]/Y vssd vssd vccd vccd output797/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_9_564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output755_A output755/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output922_A output922/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[73\]_B mprj_logic_high_inst/HI[403] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[63\]_A _655_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput850 output850/A vssd vssd vccd vccd la_data_in_mprj[70] sky130_fd_sc_hd__buf_2
Xoutput861 output861/A vssd vssd vccd vccd la_data_in_mprj[80] sky130_fd_sc_hd__buf_2
Xoutput872 output872/A vssd vssd vccd vccd la_data_in_mprj[90] sky130_fd_sc_hd__buf_2
Xoutput894 output894/A vssd vssd vccd vccd la_oenb_core[10] sky130_fd_sc_hd__buf_2
Xoutput883 output883/A vssd vssd vccd vccd la_oenb_core[0] sky130_fd_sc_hd__buf_2
XFILLER_47_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1117_A output1117/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[62\] input346/X mprj_logic_high_inst/HI[392] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[62\]/B sky130_fd_sc_hd__and2_1
XFILLER_41_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[64\]_B mprj_logic_high_inst/HI[394] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_2268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input117_A la_data_out_core[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[40\] _632_/A la_buf_enable\[40\]/B vssd vssd vccd vccd la_buf\[40\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_1523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[0\] _592_/Y mprj_logic_high_inst/HI[202] vssd vssd vccd
+ vccd output883/A sky130_fd_sc_hd__einvp_4
XFILLER_27_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_401_ _401_/A vssd vssd vccd vccd _401_/Y sky130_fd_sc_hd__inv_12
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1932 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_332_ _332_/A vssd vssd vccd vccd _332_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_42_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input82_A la_data_out_core[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[115\]_TE mprj_logic_high_inst/HI[317] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[119\]_A _382_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[54\]_A _646_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input486_A la_oenb_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[26\] _490_/Y la_buf\[26\]/TE vssd vssd vccd vccd output673/A sky130_fd_sc_hd__einvp_8
XFILLER_13_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_438 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[55\]_B mprj_logic_high_inst/HI[385] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_52_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output872_A output872/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[28\] input570/X repeater1125/X vssd vssd vccd vccd user_wb_dat_gates\[28\]/Y
+ sky130_fd_sc_hd__nand2_8
XFILLER_33_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[15\] input38/X user_to_mprj_in_gates\[15\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[15\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_oen_buffers\[45\]_A _637_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[14\]_TE mprj_logic_high_inst/HI[216] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_buffers\[25\] user_wb_dat_gates\[25\]/Y vssd vssd vccd vccd output1062/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_29_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[126\] input33/X user_to_mprj_in_gates\[126\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[126\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[46\]_B mprj_logic_high_inst/HI[376] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[36\]_A _628_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1067_A output1067/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput680 output680/A vssd vssd vccd vccd la_data_in_core[32] sky130_fd_sc_hd__buf_2
Xoutput691 output691/A vssd vssd vccd vccd la_data_in_core[42] sky130_fd_sc_hd__buf_2
XFILLER_47_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[66\] _329_/Y mprj_logic_high_inst/HI[268] vssd vssd vccd
+ vccd output973/A sky130_fd_sc_hd__einvp_2
Xla_buf_enable\[88\] _351_/A la_buf_enable\[88\]/B vssd vssd vccd vccd la_buf\[88\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_8_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[14\] _446_/Y mprj_dat_buf\[14\]/TE vssd vssd vccd vccd output1082/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_19_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input234_A la_data_out_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[37\]_B mprj_logic_high_inst/HI[367] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_2043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[52\]_TE la_buf\[52\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input401_A la_oenb_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[37\]_TE mprj_logic_high_inst/HI[239] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_72 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput37 la_data_out_core[14] vssd vssd vccd vccd input37/X sky130_fd_sc_hd__buf_4
Xinput26 la_data_out_core[11] vssd vssd vccd vccd input26/X sky130_fd_sc_hd__clkbuf_4
Xinput15 la_data_out_core[10] vssd vssd vccd vccd input15/X sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_oen_buffers\[27\]_A _619_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput59 la_data_out_core[34] vssd vssd vccd vccd input59/X sky130_fd_sc_hd__buf_4
Xinput48 la_data_out_core[24] vssd vssd vccd vccd input48/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_2114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[123\] user_to_mprj_in_gates\[123\]/Y vssd vssd vccd vccd
+ output781/A sky130_fd_sc_hd__clkinv_4
XANTENNA_output718_A output718/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[23\]_A _423_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[28\]_B mprj_logic_high_inst/HI[358] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_37_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[0\]_A _592_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[18\]_A _610_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput419 la_oenb_mprj[12] vssd vssd vccd vccd _604_/A sky130_fd_sc_hd__clkbuf_2
Xinput408 la_oenb_mprj[118] vssd vssd vccd vccd _381_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[75\]_TE la_buf\[75\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[14\]_A _414_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[19\]_B mprj_logic_high_inst/HI[349] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_43_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[25\] input305/X mprj_logic_high_inst/HI[355] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[25\]/B sky130_fd_sc_hd__and2_1
XFILLER_52_750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input184_A la_data_out_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input449_A la_oenb_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input351_A la_iena_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input45_A la_data_out_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[93\] _557_/Y la_buf\[93\]/TE vssd vssd vccd vccd output747/A sky130_fd_sc_hd__einvp_4
XANTENNA_input616_A mprj_sel_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[24\]_TE mprj_dat_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[3\]_TE mprj_logic_high_inst/HI[205] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_1194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output668_A output668/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output835_A output835/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[98\]_TE la_buf\[98\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[82\] input112/X user_to_mprj_in_gates\[82\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[82\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput205 la_data_out_mprj[50] vssd vssd vccd vccd _514_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput216 la_data_out_mprj[60] vssd vssd vccd vccd _524_/A sky130_fd_sc_hd__clkbuf_2
Xinput227 la_data_out_mprj[70] vssd vssd vccd vccd _534_/A sky130_fd_sc_hd__buf_2
Xinput238 la_data_out_mprj[80] vssd vssd vccd vccd _544_/A sky130_fd_sc_hd__buf_4
Xinput249 la_data_out_mprj[90] vssd vssd vccd vccd _554_/A sky130_fd_sc_hd__clkbuf_2
X_580_ _580_/A vssd vssd vccd vccd _580_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[29\] _621_/Y mprj_logic_high_inst/HI[231] vssd vssd vccd
+ vccd output932/A sky130_fd_sc_hd__einvp_2
XFILLER_31_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_731 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input399_A la_oenb_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input566_A mprj_dat_i_user[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1066 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[4\] _468_/Y la_buf\[4\]/TE vssd vssd vccd vccd output699/A sky130_fd_sc_hd__einvp_8
XFILLER_49_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_654 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[113\]_A_N _376_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__401__A _401_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[1\] _401_/Y mprj_adr_buf\[1\]/TE vssd vssd vccd vccd output1023/A sky130_fd_sc_hd__einvp_4
XFILLER_23_1714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[27\]_A _459_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[52\] user_to_mprj_in_gates\[52\]/Y vssd vssd vccd vccd output830/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_1_1554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output785_A output785/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1832 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_gates\[10\] input551/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[10\]/Y
+ sky130_fd_sc_hd__nand2_2
XANTENNA_output952_A output952/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[18\]_A _450_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_buffers\[25\]_A user_wb_dat_gates\[25\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_39_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1954 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[100\]_TE la_buf\[100\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1998 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[15\]_TE mprj_adr_buf\[15\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[92\] input379/X mprj_logic_high_inst/HI[422] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[92\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input147_A la_data_out_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[70\] _333_/A la_buf_enable\[70\]/B vssd vssd vccd vccd la_buf\[70\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_28_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[16\]_A user_wb_dat_gates\[16\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
X_632_ _632_/A vssd vssd vccd vccd _632_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_1368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input314_A la_iena_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_563_ _563_/A vssd vssd vccd vccd _563_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_44_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[56\] _520_/Y la_buf\[56\]/TE vssd vssd vccd vccd output706/A sky130_fd_sc_hd__einvp_8
X_494_ _494_/A vssd vssd vccd vccd _494_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_wb_ena_buf input614/X user_to_mprj_wb_ena_buf/B vssd vssd vccd vccd
+ repeater1125/A sky130_fd_sc_hd__and2_4
XFILLER_9_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[112\] _576_/Y la_buf\[112\]/TE vssd vssd vccd vccd output641/A sky130_fd_sc_hd__einvp_4
XFILLER_49_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output700_A output700/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[3\]_TE mprj_dat_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput580 mprj_dat_i_user[8] vssd vssd vccd vccd input580/X sky130_fd_sc_hd__clkbuf_16
Xinput591 mprj_dat_o_core[18] vssd vssd vccd vccd _450_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_1649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[120\]_B la_buf_enable\[120\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[45\] input71/X user_to_mprj_in_gates\[45\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[45\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[123\]_TE la_buf\[123\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[7\] input109/X user_to_mprj_in_gates\[7\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[7\]/Y sky130_fd_sc_hd__nand2_2
XANTENNA_user_wb_dat_gates\[29\]_B repeater1125/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1097_A output1097/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[111\]_B la_buf_enable\[111\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[70\]_TE mprj_logic_high_inst/HI[272] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_buffers\[2\]_A user_wb_dat_gates\[2\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[96\] _359_/Y mprj_logic_high_inst/HI[298] vssd vssd vccd
+ vccd output1006/A sky130_fd_sc_hd__einvp_2
XFILLER_13_1779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[80\]_A input110/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input264_A la_iena_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input431_A la_oenb_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_476 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input529_A mprj_adr_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[9\] input387/X mprj_logic_high_inst/HI[339] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[9\]/B sky130_fd_sc_hd__and2_1
Xla_buf_enable\[119\] _382_/A la_buf_enable\[119\]/B vssd vssd vccd vccd la_buf\[119\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_24_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[5\]_A _469_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_615_ _615_/A vssd vssd vccd vccd _615_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[102\]_B la_buf_enable\[102\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_546_ _546_/A vssd vssd vccd vccd _546_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_477_ _477_/A vssd vssd vccd vccd _477_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[15\] user_to_mprj_in_gates\[15\]/Y vssd vssd vccd vccd output789/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output650_A output650/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output748_A output748/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[71\]_A input100/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output915_A output915/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[93\]_TE mprj_logic_high_inst/HI[295] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_19 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[62\]_A input90/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj2_pwrgood mprj2_pwrgood/A vssd vssd vccd vccd output1117/A sky130_fd_sc_hd__buf_12
Xoutput840 output840/A vssd vssd vccd vccd la_data_in_mprj[61] sky130_fd_sc_hd__buf_2
Xoutput851 output851/A vssd vssd vccd vccd la_data_in_mprj[71] sky130_fd_sc_hd__buf_2
Xoutput862 output862/A vssd vssd vccd vccd la_data_in_mprj[81] sky130_fd_sc_hd__buf_2
Xoutput873 output873/A vssd vssd vccd vccd la_data_in_mprj[91] sky130_fd_sc_hd__buf_2
Xoutput895 output895/A vssd vssd vccd vccd la_oenb_core[110] sky130_fd_sc_hd__buf_2
Xoutput884 output884/A vssd vssd vccd vccd la_oenb_core[100] sky130_fd_sc_hd__buf_2
XFILLER_43_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1012_A output1012/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[55\] input338/X mprj_logic_high_inst/HI[385] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[55\]/B sky130_fd_sc_hd__and2_1
XFILLER_41_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_400_ _400_/A vssd vssd vccd vccd _400_/Y sky130_fd_sc_hd__inv_2
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[11\] _603_/Y mprj_logic_high_inst/HI[213] vssd vssd vccd
+ vccd output905/A sky130_fd_sc_hd__einvp_4
XTAP_1557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_331_ _331_/A vssd vssd vccd vccd _331_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_19_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[33\] _625_/A la_buf_enable\[33\]/B vssd vssd vccd vccd la_buf\[33\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_in_buffers\[7\] user_to_mprj_in_gates\[7\]/Y vssd vssd vccd vccd output860/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_35_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input381_A la_iena_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[71\]_A_N _334_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input479_A la_oenb_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input75_A la_data_out_core[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[19\] _483_/Y la_buf\[19\]/TE vssd vssd vccd vccd output665/A sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[53\]_A input80/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[86\]_A_N _349_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_24 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_68 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output698_A output698/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[24\]_A_N _616_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[3\]_A user_to_mprj_in_gates\[3\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_529_ _529_/A vssd vssd vccd vccd _529_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output865_A output865/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[39\]_A_N _631_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[44\]_A input70/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[18\] user_wb_dat_gates\[18\]/Y vssd vssd vccd vccd output1054/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_29_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_vdd_pwrgood_A mprj_vdd_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[119\] input25/X user_to_mprj_in_gates\[119\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[119\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1298 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_932 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[35\]_A input60/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_6 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput681 output681/A vssd vssd vccd vccd la_data_in_core[33] sky130_fd_sc_hd__buf_2
Xoutput670 output670/A vssd vssd vccd vccd la_data_in_core[23] sky130_fd_sc_hd__buf_2
Xoutput692 output692/A vssd vssd vccd vccd la_data_in_core[43] sky130_fd_sc_hd__buf_2
XFILLER_47_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[59\] _651_/Y mprj_logic_high_inst/HI[261] vssd vssd vccd
+ vccd output965/A sky130_fd_sc_hd__einvp_2
XFILLER_8_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input227_A la_data_out_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input596_A mprj_dat_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[110\] input272/X mprj_logic_high_inst/HI[440] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[110\]/B sky130_fd_sc_hd__and2_1
Xinput27 la_data_out_core[120] vssd vssd vccd vccd input27/X sky130_fd_sc_hd__buf_2
Xinput16 la_data_out_core[110] vssd vssd vccd vccd input16/X sky130_fd_sc_hd__buf_4
XFILLER_11_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput49 la_data_out_core[25] vssd vssd vccd vccd input49/X sky130_fd_sc_hd__clkbuf_4
Xinput38 la_data_out_core[15] vssd vssd vccd vccd input38/X sky130_fd_sc_hd__buf_4
XANTENNA_user_to_mprj_in_gates\[26\]_A input50/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__404__A _404_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[110\]_A input16/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[116\] user_to_mprj_in_gates\[116\]/Y vssd vssd vccd vccd
+ output773/A sky130_fd_sc_hd__clkinv_4
XFILLER_2_582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[82\] user_to_mprj_in_gates\[82\]/Y vssd vssd vccd vccd output863/A
+ sky130_fd_sc_hd__inv_2
XFILLER_37_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output982_A output982/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_rstn_buf_A input3/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[17\]_A input40/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[101\]_A input6/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput409 la_oenb_mprj[119] vssd vssd vccd vccd _382_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[105\]_TE mprj_logic_high_inst/HI[307] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[18\] input297/X mprj_logic_high_inst/HI[348] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[18\]/B sky130_fd_sc_hd__and2_1
XFILLER_12_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input177_A la_data_out_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input344_A la_iena_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input38_A la_data_out_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input511_A la_oenb_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[86\] _550_/Y la_buf\[86\]/TE vssd vssd vccd vccd output739/A sky130_fd_sc_hd__einvp_2
XFILLER_19_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input609_A mprj_dat_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_718 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[101\] _364_/A la_buf_enable\[101\]/B vssd vssd vccd vccd la_buf\[101\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_1_1725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2016 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output730_A output730/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output828_A output828/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[75\] input104/X user_to_mprj_in_gates\[75\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[75\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[123\]_A input286/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[42\]_TE la_buf\[42\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[27\]_TE mprj_logic_high_inst/HI[229] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xinput206 la_data_out_mprj[51] vssd vssd vccd vccd _515_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput217 la_data_out_mprj[61] vssd vssd vccd vccd _525_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput228 la_data_out_mprj[71] vssd vssd vccd vccd _535_/A sky130_fd_sc_hd__buf_2
Xinput239 la_data_out_mprj[81] vssd vssd vccd vccd _545_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[114\]_A input276/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input294_A la_iena_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input559_A mprj_dat_i_user[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input461_A la_oenb_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_ena_buf\[1\] input625/X user_irq_ena_buf\[1\]/B vssd vssd vccd vccd user_irq_gates\[1\]/B
+ sky130_fd_sc_hd__and2_1
XFILLER_45_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[105\]_A input266/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output680_A output680/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[45\] user_to_mprj_in_gates\[45\]/Y vssd vssd vccd vccd output822/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_31_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output778_A output778/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[65\]_TE la_buf\[65\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output945_A output945/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[101\] input6/X user_to_mprj_in_gates\[101\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[101\]/Y sky130_fd_sc_hd__nand2_1
XTAP_1909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output1042_A output1042/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[14\]_TE mprj_dat_buf\[14\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__502__A _502_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[85\] input371/X mprj_logic_high_inst/HI[415] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[85\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[111\] _374_/Y mprj_logic_high_inst/HI[313] vssd vssd vccd
+ vccd output896/A sky130_fd_sc_hd__einvp_4
XFILLER_48_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[94\]_A input381/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[41\] _633_/Y mprj_logic_high_inst/HI[243] vssd vssd vccd
+ vccd output946/A sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[63\] _655_/A la_buf_enable\[63\]/B vssd vssd vccd vccd la_buf\[63\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_28_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_631_ _631_/A vssd vssd vccd vccd _631_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_562_ _562_/A vssd vssd vccd vccd _562_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_44_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input307_A la_iena_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_493_ _493_/A vssd vssd vccd vccd _493_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[88\]_TE la_buf\[88\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[49\] _513_/Y la_buf\[49\]/TE vssd vssd vccd vccd output698/A sky130_fd_sc_hd__einvp_4
XFILLER_34_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1432 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__412__A _412_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[105\] _569_/Y la_buf\[105\]/TE vssd vssd vccd vccd output633/A sky130_fd_sc_hd__einvp_4
XFILLER_45_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[85\]_A input371/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput570 mprj_dat_i_user[28] vssd vssd vccd vccd input570/X sky130_fd_sc_hd__clkbuf_2
Xinput581 mprj_dat_i_user[9] vssd vssd vccd vccd input581/X sky130_fd_sc_hd__clkbuf_16
XFILLER_36_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput592 mprj_dat_o_core[19] vssd vssd vccd vccd _451_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_output895_A output895/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[38\] input63/X user_to_mprj_in_gates\[38\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[38\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[76\]_A input361/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[112\]_A_N _375_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[127\]_A_N _390_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[80\]_B user_to_mprj_in_gates\[80\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[89\] _352_/Y mprj_logic_high_inst/HI[291] vssd vssd vccd
+ vccd output998/A sky130_fd_sc_hd__einvp_4
XFILLER_2_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input257_A la_data_out_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input20_A la_data_out_core[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input424_A la_oenb_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[67\]_A input351/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_614_ _614_/A vssd vssd vccd vccd _614_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_545_ _545_/A vssd vssd vccd vccd _545_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_476_ _476_/A vssd vssd vccd vccd _476_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_18_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__407__A _407_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[71\]_B user_to_mprj_in_gates\[71\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output643_A output643/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output810_A output810/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output908_A output908/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[58\]_A input341/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1026 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[62\]_B user_to_mprj_in_gates\[62\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xoutput830 output830/A vssd vssd vccd vccd la_data_in_mprj[52] sky130_fd_sc_hd__buf_2
Xoutput841 output841/A vssd vssd vccd vccd la_data_in_mprj[62] sky130_fd_sc_hd__buf_2
Xoutput852 output852/A vssd vssd vccd vccd la_data_in_mprj[72] sky130_fd_sc_hd__buf_2
Xoutput863 output863/A vssd vssd vccd vccd la_data_in_mprj[82] sky130_fd_sc_hd__buf_2
Xoutput896 output896/A vssd vssd vccd vccd la_oenb_core[111] sky130_fd_sc_hd__buf_2
Xoutput885 output885/A vssd vssd vccd vccd la_oenb_core[101] sky130_fd_sc_hd__buf_2
Xoutput874 output874/A vssd vssd vccd vccd la_data_in_mprj[92] sky130_fd_sc_hd__buf_2
XFILLER_43_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[49\]_A input331/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output1005_A output1005/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[48\] input330/X mprj_logic_high_inst/HI[378] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[48\]/B sky130_fd_sc_hd__and2_1
XTAP_2226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_330_ _330_/A vssd vssd vccd vccd _330_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_43 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[26\] _618_/A la_buf_enable\[26\]/B vssd vssd vccd vccd la_buf\[26\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_22_370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[53\]_B user_to_mprj_in_gates\[53\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input374_A la_iena_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input68_A la_data_out_core[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input541_A mprj_adr_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[113\]_TE la_buf\[113\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_764 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[28\]_TE mprj_adr_buf\[28\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_47 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_528_ _528_/A vssd vssd vccd vccd _528_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_mprj_dat_buf\[7\]_A _439_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_459_ _459_/A vssd vssd vccd vccd _459_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_20_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output858_A output858/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output760_A output760/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[44\]_B user_to_mprj_in_gates\[44\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__600__A _600_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[60\]_TE mprj_logic_high_inst/HI[262] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1290 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[35\]_B user_to_mprj_in_gates\[35\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[96\]_A user_to_mprj_in_gates\[96\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput671 output671/A vssd vssd vccd vccd la_data_in_core[24] sky130_fd_sc_hd__buf_2
Xoutput660 output660/A vssd vssd vccd vccd la_data_in_core[14] sky130_fd_sc_hd__buf_2
XANTENNA_output1122_A output1122/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput693 output693/A vssd vssd vccd vccd la_data_in_core[44] sky130_fd_sc_hd__buf_2
Xoutput682 output682/A vssd vssd vccd vccd la_data_in_core[34] sky130_fd_sc_hd__buf_2
XFILLER_47_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__510__A _510_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input122_A la_data_out_core[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1824 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[20\]_A user_to_mprj_in_gates\[20\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_2056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input491_A la_oenb_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2080 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input589_A mprj_dat_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput28 la_data_out_core[121] vssd vssd vccd vccd input28/X sky130_fd_sc_hd__clkbuf_4
Xinput17 la_data_out_core[111] vssd vssd vccd vccd input17/X sky130_fd_sc_hd__buf_4
XFILLER_52_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[123\]_A _587_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[31\] _495_/Y la_buf\[31\]/TE vssd vssd vccd vccd output679/A sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[103\] input264/X mprj_logic_high_inst/HI[433] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[103\]/B sky130_fd_sc_hd__and2_1
XFILLER_11_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_gates\[3\] input575/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[3\]/Y
+ sky130_fd_sc_hd__nand2_4
Xinput39 la_data_out_core[16] vssd vssd vccd vccd input39/X sky130_fd_sc_hd__buf_4
XANTENNA_user_to_mprj_in_gates\[26\]_B user_to_mprj_in_gates\[26\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[87\]_A user_to_mprj_in_gates\[87\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[110\]_B user_to_mprj_in_gates\[110\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[60\]_A _524_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[83\]_TE mprj_logic_high_inst/HI[285] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__420__A _420_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[109\] user_to_mprj_in_gates\[109\]/Y vssd vssd vccd vccd
+ output765/A sky130_fd_sc_hd__clkinv_4
XFILLER_4_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[75\] user_to_mprj_in_gates\[75\]/Y vssd vssd vccd vccd output855/A
+ sky130_fd_sc_hd__clkinv_2
XFILLER_4_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[11\]_A user_to_mprj_in_gates\[11\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_46_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output975_A output975/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[20\] input44/X user_to_mprj_in_gates\[20\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[20\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_1132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[125\]_A user_to_mprj_in_gates\[125\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[114\]_A _578_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[17\]_B user_to_mprj_in_gates\[17\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[30\] user_wb_dat_gates\[30\]/Y vssd vssd vccd vccd output1068/A
+ sky130_fd_sc_hd__inv_6
XFILLER_31_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[78\]_A user_to_mprj_in_gates\[78\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_B user_to_mprj_in_gates\[101\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[51\]_A _515_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__330__A _330_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[8\] _440_/Y mprj_dat_buf\[8\]/TE vssd vssd vccd vccd output1107/A sky130_fd_sc_hd__einvp_8
XFILLER_9_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[70\]_A_N _333_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[10\]_A input551/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[85\]_A_N _348_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[116\]_A user_to_mprj_in_gates\[116\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1072_A output1072/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[105\]_A _569_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__505__A _505_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[69\]_A user_to_mprj_in_gates\[69\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[42\]_A _506_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[71\] _334_/Y mprj_logic_high_inst/HI[273] vssd vssd vccd
+ vccd output979/A sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[60\]_B la_buf_enable\[60\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[23\]_A_N _615_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[93\] _356_/A la_buf_enable\[93\]/B vssd vssd vccd vccd la_buf\[93\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_47_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input337_A la_iena_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[38\]_A_N _630_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[79\] _543_/Y la_buf\[79\]/TE vssd vssd vccd vccd output731/A sky130_fd_sc_hd__einvp_2
XANTENNA_input504_A la_oenb_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[107\]_A user_to_mprj_in_gates\[107\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__415__A _415_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[33\]_A _497_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output723_A output723/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[51\]_B la_buf_enable\[51\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[68\] input96/X user_to_mprj_in_gates\[68\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[68\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[123\]_B mprj_logic_high_inst/HI[453] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[24\]_A _488_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[42\]_B la_buf_enable\[42\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput207 la_data_out_mprj[52] vssd vssd vccd vccd _516_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput218 la_data_out_mprj[62] vssd vssd vccd vccd _526_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput229 la_data_out_mprj[72] vssd vssd vccd vccd _536_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[114\]_B mprj_logic_high_inst/HI[444] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[30\] input311/X mprj_logic_high_inst/HI[360] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[30\]/B sky130_fd_sc_hd__and2_1
XFILLER_25_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input287_A la_iena_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[15\]_A _479_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input454_A la_oenb_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input50_A la_data_out_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[33\]_B la_buf_enable\[33\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input621_A user_irq_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[2\]_A input310/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[100\]_A _363_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[105\]_B mprj_logic_high_inst/HI[435] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_788 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[38\] user_to_mprj_in_gates\[38\]/Y vssd vssd vccd vccd output814/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output673_A output673/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output938_A output938/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output840_A output840/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[24\]_B la_buf_enable\[24\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[93\]_A _356_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output1035_A output1035/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[15\]_B la_buf_enable\[15\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[78\] input363/X mprj_logic_high_inst/HI[408] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[78\]/B sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[104\] _367_/Y mprj_logic_high_inst/HI[306] vssd vssd vccd
+ vccd output888/A sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[94\]_B mprj_logic_high_inst/HI[424] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_630_ _630_/A vssd vssd vccd vccd _630_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[56\] _648_/A la_buf_enable\[56\]/B vssd vssd vccd vccd la_buf\[56\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[34\] _626_/Y mprj_logic_high_inst/HI[236] vssd vssd vccd
+ vccd output938/A sky130_fd_sc_hd__einvp_4
X_561_ _561_/A vssd vssd vccd vccd _561_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_492_ _492_/A vssd vssd vccd vccd _492_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input202_A la_data_out_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2290 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[84\]_A _347_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[118\]_TE mprj_logic_high_inst/HI[320] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input98_A la_data_out_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input571_A mprj_dat_i_user[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_998 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput571 mprj_dat_i_user[29] vssd vssd vccd vccd input571/X sky130_fd_sc_hd__clkbuf_2
Xinput560 mprj_dat_i_user[19] vssd vssd vccd vccd input560/X sky130_fd_sc_hd__buf_12
XANTENNA_user_to_mprj_in_ena_buf\[85\]_B mprj_logic_high_inst/HI[415] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xinput582 mprj_dat_o_core[0] vssd vssd vccd vccd _432_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_2021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput593 mprj_dat_o_core[1] vssd vssd vccd vccd _433_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[32\]_TE la_buf\[32\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output790_A output790/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output888_A output888/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[75\]_A _338_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[17\]_TE mprj_logic_high_inst/HI[219] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__603__A _603_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[2\]_A input572/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[76\]_B mprj_logic_high_inst/HI[406] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[2\]_A input54/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[66\]_A _329_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1731 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[0\]_TE la_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__513__A _513_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input152_A la_data_out_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[67\]_B mprj_logic_high_inst/HI[397] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[55\]_TE la_buf\[55\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_613_ _613_/A vssd vssd vccd vccd _613_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input417_A la_oenb_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input13_A la_data_out_core[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[61\] _525_/Y la_buf\[61\]/TE vssd vssd vccd vccd output712/A sky130_fd_sc_hd__einvp_8
XFILLER_33_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_544_ _544_/A vssd vssd vccd vccd _544_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_475_ _475_/A vssd vssd vccd vccd _475_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[57\]_A _649_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[25\] _425_/Y mprj_adr_buf\[25\]/TE vssd vssd vccd vccd output1029/A
+ sky130_fd_sc_hd__einvp_8
XANTENNA__423__A _423_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output636_A output636/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output803_A output803/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[58\]_B mprj_logic_high_inst/HI[388] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput390 la_oenb_mprj[101] vssd vssd vccd vccd _364_/A sky130_fd_sc_hd__clkbuf_4
Xuser_to_mprj_in_gates\[50\] input77/X user_to_mprj_in_gates\[50\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[50\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[48\]_A _640_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__333__A _333_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput820 output820/A vssd vssd vccd vccd la_data_in_mprj[43] sky130_fd_sc_hd__buf_2
Xoutput831 output831/A vssd vssd vccd vccd la_data_in_mprj[53] sky130_fd_sc_hd__buf_2
Xoutput842 output842/A vssd vssd vccd vccd la_data_in_mprj[63] sky130_fd_sc_hd__buf_2
Xoutput853 output853/A vssd vssd vccd vccd la_data_in_mprj[73] sky130_fd_sc_hd__buf_2
Xoutput864 output864/A vssd vssd vccd vccd la_data_in_mprj[83] sky130_fd_sc_hd__buf_2
Xoutput886 output886/A vssd vssd vccd vccd la_oenb_core[102] sky130_fd_sc_hd__buf_2
Xoutput897 output897/A vssd vssd vccd vccd la_oenb_core[112] sky130_fd_sc_hd__buf_2
XANTENNA_la_buf\[78\]_TE la_buf\[78\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput875 output875/A vssd vssd vccd vccd la_data_in_mprj[93] sky130_fd_sc_hd__buf_2
XANTENNA_input5_A la_data_out_core[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[49\]_B mprj_logic_high_inst/HI[379] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__508__A _508_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[39\]_A _631_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[19\] _611_/A la_buf_enable\[19\]/B vssd vssd vccd vccd la_buf\[19\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_52_1572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input367_A la_iena_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_irq_gates\[2\] input623/X user_irq_gates\[2\]/B vssd vssd vccd vccd user_irq_gates\[2\]/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_29_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input534_A mprj_adr_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[124\] _387_/A la_buf_enable\[124\]/B vssd vssd vccd vccd la_buf\[124\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[27\]_TE mprj_dat_buf\[27\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_527_ _527_/A vssd vssd vccd vccd _527_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__418__A _418_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[6\]_TE mprj_logic_high_inst/HI[208] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_458_ _458_/A vssd vssd vccd vccd _458_/Y sky130_fd_sc_hd__inv_6
XFILLER_32_157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_389_ _389_/A vssd vssd vccd vccd _389_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[20\] user_to_mprj_in_gates\[20\]/Y vssd vssd vccd vccd output795/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_9_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output753_A output753/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output920_A output920/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[98\] input129/X user_to_mprj_in_gates\[98\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[98\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[26\]_A _426_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[111\]_A_N _374_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[126\]_A_N _389_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[3\]_A _595_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput650 output650/A vssd vssd vccd vccd la_data_in_core[120] sky130_fd_sc_hd__buf_2
Xoutput672 output672/A vssd vssd vccd vccd la_data_in_core[25] sky130_fd_sc_hd__buf_2
Xoutput661 output661/A vssd vssd vccd vccd la_data_in_core[15] sky130_fd_sc_hd__buf_2
Xoutput694 output694/A vssd vssd vccd vccd la_data_in_core[45] sky130_fd_sc_hd__buf_2
Xoutput683 output683/A vssd vssd vccd vccd la_data_in_core[35] sky130_fd_sc_hd__buf_2
XFILLER_43_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output1115_A output1115/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[17\]_A _417_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[60\] input344/X mprj_logic_high_inst/HI[390] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[60\]/B sky130_fd_sc_hd__and2_1
XFILLER_25_1950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_sel_buf\[1\]_TE mprj_sel_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_964 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input115_A la_data_out_core[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_64 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput18 la_data_out_core[112] vssd vssd vccd vccd input18/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_input80_A la_data_out_core[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input484_A la_oenb_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput29 la_data_out_core[122] vssd vssd vccd vccd input29/X sky130_fd_sc_hd__buf_4
Xla_buf\[24\] _488_/Y la_buf\[24\]/TE vssd vssd vccd vccd output671/A sky130_fd_sc_hd__einvp_8
XFILLER_32_1976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_irq_buffers\[0\]_A user_irq_gates\[0\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[68\] user_to_mprj_in_gates\[68\]/Y vssd vssd vccd vccd output847/A
+ sky130_fd_sc_hd__inv_2
XFILLER_45_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output870_A output870/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output968_A output968/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[26\] input568/X repeater1125/X vssd vssd vccd vccd user_wb_dat_gates\[26\]/Y
+ sky130_fd_sc_hd__nand2_8
XTAP_1890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[13\] input36/X user_to_mprj_in_gates\[13\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[13\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_buffers\[23\] user_wb_dat_gates\[23\]/Y vssd vssd vccd vccd output1060/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_31_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__611__A _611_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[124\] input31/X user_to_mprj_in_gates\[124\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[124\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[10\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_764 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[103\]_TE la_buf\[103\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[18\]_TE mprj_adr_buf\[18\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1065_A output1065/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__521__A _521_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[2\]_TE mprj_adr_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[64\] _656_/Y mprj_logic_high_inst/HI[266] vssd vssd vccd
+ vccd output971/A sky130_fd_sc_hd__einvp_4
Xla_buf_enable\[86\] _349_/A la_buf_enable\[86\]/B vssd vssd vccd vccd la_buf\[86\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_43_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[12\] _444_/Y mprj_dat_buf\[12\]/TE vssd vssd vccd vccd output1080/A
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input232_A la_data_out_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_cyc_buf_A _393_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[50\]_TE mprj_logic_high_inst/HI[252] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__431__A _431_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[121\] user_to_mprj_in_gates\[121\]/Y vssd vssd vccd vccd
+ output779/A sky130_fd_sc_hd__clkinv_4
XFILLER_3_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[6\]_TE mprj_dat_buf\[6\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output716_A output716/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[126\]_TE la_buf\[126\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__606__A _606_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[2\]_A _402_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__341__A _341_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput208 la_data_out_mprj[53] vssd vssd vccd vccd _517_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_wb_dat_buffers\[28\]_A user_wb_dat_gates\[28\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_29_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput219 la_data_out_mprj[63] vssd vssd vccd vccd _527_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[73\]_TE mprj_logic_high_inst/HI[275] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[23\] input303/X mprj_logic_high_inst/HI[353] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[23\]/B sky130_fd_sc_hd__and2_1
XFILLER_12_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__516__A _516_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_296 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_77 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input182_A la_data_out_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input447_A la_oenb_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input43_A la_data_out_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_buffers\[19\]_A user_wb_dat_gates\[19\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_43_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[2\]_B mprj_logic_high_inst/HI[332] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf\[91\] _555_/Y la_buf\[91\]/TE vssd vssd vccd vccd output745/A sky130_fd_sc_hd__einvp_8
XANTENNA_input614_A mprj_iena_wb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__426__A _426_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output666_A output666/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output833_A output833/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[80\] input110/X user_to_mprj_in_gates\[80\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[80\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[84\]_A_N _347_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[123\]_B la_buf_enable\[123\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[96\]_TE mprj_logic_high_inst/HI[298] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[99\]_A_N _362_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[22\]_A_N _614_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__336__A _336_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[92\]_A input123/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[37\]_A_N _629_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output1028_A output1028/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_66 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[114\]_B la_buf_enable\[114\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_560_ _560_/A vssd vssd vccd vccd _560_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[49\] _641_/A la_buf_enable\[49\]/B vssd vssd vccd vccd la_buf\[49\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[27\] _619_/Y mprj_logic_high_inst/HI[229] vssd vssd vccd
+ vccd output930/A sky130_fd_sc_hd__einvp_2
Xuser_to_mprj_oen_buffers\[9\] _601_/Y mprj_logic_high_inst/HI[211] vssd vssd vccd
+ vccd output1010/A sky130_fd_sc_hd__einvp_4
X_491_ _491_/A vssd vssd vccd vccd _491_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_25_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_buffers\[5\]_A user_wb_dat_gates\[5\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input397_A la_oenb_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[83\]_A input113/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input564_A mprj_dat_i_user[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[2\] _466_/Y la_buf\[2\]/TE vssd vssd vccd vccd output677/A sky130_fd_sc_hd__einvp_8
XFILLER_5_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput572 mprj_dat_i_user[2] vssd vssd vccd vccd input572/X sky130_fd_sc_hd__buf_8
Xinput550 mprj_dat_i_user[0] vssd vssd vccd vccd input550/X sky130_fd_sc_hd__buf_12
Xinput561 mprj_dat_i_user[1] vssd vssd vccd vccd input561/X sky130_fd_sc_hd__clkbuf_16
XANTENNA_la_buf\[8\]_A _472_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[105\]_B la_buf_enable\[105\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput583 mprj_dat_o_core[10] vssd vssd vccd vccd _442_/A sky130_fd_sc_hd__clkbuf_2
Xinput594 mprj_dat_o_core[20] vssd vssd vccd vccd _452_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[50\] user_to_mprj_in_gates\[50\]/Y vssd vssd vccd vccd output828/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_44_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output783_A output783/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output950_A output950/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[74\]_A input103/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[2\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[2\]_B user_to_mprj_in_gates\[2\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_41_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[65\]_A input93/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[90\] input377/X mprj_logic_high_inst/HI[420] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[90\]/B sky130_fd_sc_hd__and2_1
XFILLER_11_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input145_A la_data_out_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_612_ _612_/A vssd vssd vccd vccd _612_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input312_A la_iena_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_543_ _543_/A vssd vssd vccd vccd _543_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1674 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_474_ _474_/A vssd vssd vccd vccd _474_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[54\] _518_/Y la_buf\[54\]/TE vssd vssd vccd vccd output704/A sky130_fd_sc_hd__einvp_8
XFILLER_25_380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[126\] input289/X mprj_logic_high_inst/HI[456] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[126\]/B sky130_fd_sc_hd__and2_1
XFILLER_13_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[56\]_A input83/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[110\] _574_/Y la_buf\[110\]/TE vssd vssd vccd vccd output639/A sky130_fd_sc_hd__einvp_2
Xmprj_adr_buf\[18\] _418_/Y mprj_adr_buf\[18\]/TE vssd vssd vccd vccd output1021/A
+ sky130_fd_sc_hd__einvp_4
XFILLER_5_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output629_A output629/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[98\] user_to_mprj_in_gates\[98\]/Y vssd vssd vccd vccd output880/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_7_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput380 la_iena_mprj[93] vssd vssd vccd vccd input380/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[6\]_A user_to_mprj_in_gates\[6\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xinput391 la_oenb_mprj[102] vssd vssd vccd vccd _365_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_output998_A output998/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[43\] input69/X user_to_mprj_in_gates\[43\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[43\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_buffers\[8\] user_wb_dat_gates\[8\]/Y vssd vssd vccd vccd output1075/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_36_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[47\]_A input73/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__614__A _614_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput821 output821/A vssd vssd vccd vccd la_data_in_mprj[44] sky130_fd_sc_hd__buf_2
Xoutput810 output810/A vssd vssd vccd vccd la_data_in_mprj[34] sky130_fd_sc_hd__buf_2
Xoutput832 output832/A vssd vssd vccd vccd la_data_in_mprj[54] sky130_fd_sc_hd__buf_2
Xoutput843 output843/A vssd vssd vccd vccd la_data_in_mprj[64] sky130_fd_sc_hd__buf_2
Xoutput854 output854/A vssd vssd vccd vccd la_data_in_mprj[74] sky130_fd_sc_hd__buf_2
Xoutput887 output887/A vssd vssd vccd vccd la_oenb_core[103] sky130_fd_sc_hd__buf_2
XFILLER_28_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[5\] input87/X user_to_mprj_in_gates\[5\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[5\]/Y sky130_fd_sc_hd__nand2_2
Xoutput865 output865/A vssd vssd vccd vccd la_data_in_mprj[84] sky130_fd_sc_hd__buf_2
Xoutput876 output876/A vssd vssd vccd vccd la_data_in_mprj[94] sky130_fd_sc_hd__buf_2
Xoutput898 output898/A vssd vssd vccd vccd la_oenb_core[113] sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_oen_buffers\[108\]_TE mprj_logic_high_inst/HI[310] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XTAP_350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1095_A output1095/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_45 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[38\]_A input63/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__524__A _524_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[122\]_A input29/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[94\] _357_/Y mprj_logic_high_inst/HI[296] vssd vssd vccd
+ vccd output1004/A sky130_fd_sc_hd__einvp_4
XFILLER_46_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input262_A la_iena_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[22\]_TE la_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input527_A mprj_adr_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[7\] input365/X mprj_logic_high_inst/HI[337] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[7\]/B sky130_fd_sc_hd__and2_1
Xla_buf_enable\[117\] _380_/A la_buf_enable\[117\]/B vssd vssd vccd vccd la_buf\[117\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_8_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_526_ _526_/A vssd vssd vccd vccd _526_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_33_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_457_ _457_/A vssd vssd vccd vccd _457_/Y sky130_fd_sc_hd__inv_4
XFILLER_20_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_388_ _388_/A vssd vssd vccd vccd _388_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[29\]_A input53/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__434__A _434_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_A input19/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[13\] user_to_mprj_in_gates\[13\]/Y vssd vssd vccd vccd output787/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_9_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output746_A output746/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output913_A output913/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__609__A _609_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__344__A _344_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[104\]_A input9/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[45\]_TE la_buf\[45\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput651 output651/A vssd vssd vccd vccd la_data_in_core[121] sky130_fd_sc_hd__buf_2
Xoutput640 output640/A vssd vssd vccd vccd la_data_in_core[111] sky130_fd_sc_hd__buf_2
Xoutput662 output662/A vssd vssd vccd vccd la_data_in_core[16] sky130_fd_sc_hd__buf_2
Xoutput695 output695/A vssd vssd vccd vccd la_data_in_core[46] sky130_fd_sc_hd__buf_2
Xoutput684 output684/A vssd vssd vccd vccd la_data_in_core[36] sky130_fd_sc_hd__buf_2
Xoutput673 output673/A vssd vssd vccd vccd la_data_in_core[26] sky130_fd_sc_hd__buf_2
XFILLER_28_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1010_A output1010/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output1108_A output1108/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[53\] input336/X mprj_logic_high_inst/HI[383] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[53\]/B sky130_fd_sc_hd__and2_1
XTAP_180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__519__A _519_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input108_A la_data_out_core[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_618 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[31\] _623_/A la_buf_enable\[31\]/B vssd vssd vccd vccd la_buf\[31\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_in_buffers\[5\] user_to_mprj_in_gates\[5\]/Y vssd vssd vccd vccd output838/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_52_2060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput19 la_data_out_core[113] vssd vssd vccd vccd input19/X sky130_fd_sc_hd__clkbuf_4
XFILLER_32_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input477_A la_oenb_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input73_A la_data_out_core[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[17\] _481_/Y la_buf\[17\]/TE vssd vssd vccd vccd output663/A sky130_fd_sc_hd__einvp_8
XFILLER_6_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__429__A _429_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output696_A output696/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_509_ _509_/A vssd vssd vccd vccd _509_/Y sky130_fd_sc_hd__inv_2
XTAP_1891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[68\]_TE la_buf\[68\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output863_A output863/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[19\] input560/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[19\]/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_31_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_buffers\[16\] user_wb_dat_gates\[16\]/Y vssd vssd vccd vccd output1052/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_29_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[2\]_B la_buf_enable\[2\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[126\]_A input289/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[117\] input23/X user_to_mprj_in_gates\[117\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[117\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA__339__A _339_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output1058_A output1058/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[17\]_TE mprj_dat_buf\[17\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[127\] _390_/Y mprj_logic_high_inst/HI[329] vssd vssd vccd
+ vccd output913/A sky130_fd_sc_hd__einvp_4
XFILLER_43_2059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[57\] _649_/Y mprj_logic_high_inst/HI[259] vssd vssd vccd
+ vccd output963/A sky130_fd_sc_hd__einvp_2
XFILLER_47_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[79\] _342_/A la_buf_enable\[79\]/B vssd vssd vccd vccd la_buf\[79\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_43_1369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_54 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[117\]_A input279/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input225_A la_data_out_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input594_A mprj_dat_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[110\]_A_N _373_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[125\]_A_N _388_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[114\] user_to_mprj_in_gates\[114\]/Y vssd vssd vccd vccd
+ output771/A sky130_fd_sc_hd__clkinv_4
XANTENNA_output709_A output709/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[80\] user_to_mprj_in_gates\[80\]/Y vssd vssd vccd vccd output861/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_4_2053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[108\]_A input269/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output980_A output980/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__622__A _622_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput1120 output1120/A vssd vssd vccd vccd user_clock2 sky130_fd_sc_hd__buf_2
Xinput209 la_data_out_mprj[54] vssd vssd vccd vccd _518_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[16\] input295/X mprj_logic_high_inst/HI[346] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[16\]/B sky130_fd_sc_hd__and2_1
XFILLER_12_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[30\]_A input311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__532__A _532_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input175_A la_data_out_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input342_A la_iena_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[97\]_A input384/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input36_A la_data_out_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[84\] _548_/Y la_buf\[84\]/TE vssd vssd vccd vccd output737/A sky130_fd_sc_hd__einvp_4
XFILLER_1_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input607_A mprj_dat_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[21\]_A input301/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output659_A output659/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__442__A _442_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output826_A output826/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[88\]_A input374/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[73\] input102/X user_to_mprj_in_gates\[73\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[73\]/Y sky130_fd_sc_hd__nand2_1
XTAP_735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__617__A _617_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_234 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[12\]_A input291/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[92\]_B user_to_mprj_in_gates\[92\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__352__A _352_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[79\]_A input364/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[40\]_TE mprj_logic_high_inst/HI[242] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__527__A _527_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_490_ _490_/A vssd vssd vccd vccd _490_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input292_A la_iena_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[83\]_B user_to_mprj_in_gates\[83\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_input557_A mprj_dat_i_user[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[116\]_TE la_buf\[116\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput573 mprj_dat_i_user[30] vssd vssd vccd vccd input573/X sky130_fd_sc_hd__clkbuf_2
Xinput562 mprj_dat_i_user[20] vssd vssd vccd vccd input562/X sky130_fd_sc_hd__clkbuf_16
Xinput551 mprj_dat_i_user[10] vssd vssd vccd vccd input551/X sky130_fd_sc_hd__buf_12
XFILLER_48_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput540 mprj_adr_o_core[30] vssd vssd vccd vccd _430_/A sky130_fd_sc_hd__buf_2
XFILLER_35_304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput584 mprj_dat_o_core[11] vssd vssd vccd vccd _443_/A sky130_fd_sc_hd__buf_2
Xinput595 mprj_dat_o_core[21] vssd vssd vccd vccd _453_/A sky130_fd_sc_hd__buf_2
XFILLER_1_1333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__437__A _437_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[43\] user_to_mprj_in_gates\[43\]/Y vssd vssd vccd vccd output820/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_16_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output776_A output776/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[74\]_B user_to_mprj_in_gates\[74\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output943_A output943/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[63\]_TE mprj_logic_high_inst/HI[265] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XTAP_510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__347__A _347_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[65\]_B user_to_mprj_in_gates\[65\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output1040_A output1040/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[83\] input369/X mprj_logic_high_inst/HI[413] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[83\]/B sky130_fd_sc_hd__and2_1
XFILLER_11_1496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[61\] _653_/A la_buf_enable\[61\]/B vssd vssd vccd vccd la_buf\[61\]/TE
+ sky130_fd_sc_hd__and2b_1
X_611_ _611_/A vssd vssd vccd vccd _611_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input138_A la_data_out_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[50\]_A user_to_mprj_in_gates\[50\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_542_ _542_/A vssd vssd vccd vccd _542_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input305_A la_iena_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_473_ _473_/A vssd vssd vccd vccd _473_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[47\] _511_/Y la_buf\[47\]/TE vssd vssd vccd vccd output696/A sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[83\]_A_N _346_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[56\]_B user_to_mprj_in_gates\[56\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[119\] input281/X mprj_logic_high_inst/HI[449] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[119\]/B sky130_fd_sc_hd__and2_1
XFILLER_13_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[90\]_A _554_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1298 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[86\]_TE mprj_logic_high_inst/HI[288] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[98\]_A_N _361_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[103\] _567_/Y la_buf\[103\]/TE vssd vssd vccd vccd output631/A sky130_fd_sc_hd__einvp_2
XANTENNA_la_buf_enable\[21\]_A_N _613_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[41\]_A user_to_mprj_in_gates\[41\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xinput370 la_iena_mprj[84] vssd vssd vccd vccd input370/X sky130_fd_sc_hd__clkbuf_1
Xinput381 la_iena_mprj[94] vssd vssd vccd vccd input381/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput392 la_oenb_mprj[103] vssd vssd vccd vccd _366_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_output893_A output893/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[36\]_A_N _628_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[36\] input61/X user_to_mprj_in_gates\[36\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[36\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_1163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[47\]_B user_to_mprj_in_gates\[47\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[81\]_A _545_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput800 output800/A vssd vssd vccd vccd la_data_in_mprj[25] sky130_fd_sc_hd__buf_2
Xoutput811 output811/A vssd vssd vccd vccd la_data_in_mprj[35] sky130_fd_sc_hd__buf_2
Xoutput833 output833/A vssd vssd vccd vccd la_data_in_mprj[55] sky130_fd_sc_hd__buf_2
Xoutput822 output822/A vssd vssd vccd vccd la_data_in_mprj[45] sky130_fd_sc_hd__buf_2
Xoutput844 output844/A vssd vssd vccd vccd la_data_in_mprj[65] sky130_fd_sc_hd__buf_2
Xoutput855 output855/A vssd vssd vccd vccd la_data_in_mprj[75] sky130_fd_sc_hd__buf_2
XFILLER_8_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__630__A _630_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput888 output888/A vssd vssd vccd vccd la_oenb_core[104] sky130_fd_sc_hd__buf_2
XFILLER_28_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput866 output866/A vssd vssd vccd vccd la_data_in_mprj[85] sky130_fd_sc_hd__buf_2
Xoutput877 output877/A vssd vssd vccd vccd la_data_in_mprj[95] sky130_fd_sc_hd__buf_2
Xoutput899 output899/A vssd vssd vccd vccd la_oenb_core[114] sky130_fd_sc_hd__buf_2
XTAP_351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[32\]_A user_to_mprj_in_gates\[32\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output1088_A output1088/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[38\]_B user_to_mprj_in_gates\[38\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[99\]_A user_to_mprj_in_gates\[99\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[122\]_B user_to_mprj_in_gates\[122\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[72\]_A _536_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[90\]_B la_buf_enable\[90\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[87\] _350_/Y mprj_logic_high_inst/HI[289] vssd vssd vccd
+ vccd output996/A sky130_fd_sc_hd__einvp_2
XANTENNA__540__A _540_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input255_A la_data_out_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[23\]_A user_to_mprj_in_gates\[23\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_input422_A la_oenb_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[31\]_A input574/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_525_ _525_/A vssd vssd vccd vccd _525_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[126\]_A _590_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_456_ _456_/A vssd vssd vccd vccd _456_/Y sky130_fd_sc_hd__inv_6
XFILLER_41_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_387_ _387_/A vssd vssd vccd vccd _387_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1040 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[29\]_B user_to_mprj_in_gates\[29\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_B user_to_mprj_in_gates\[113\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[63\]_A _527_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[30\] _430_/Y mprj_adr_buf\[30\]/TE vssd vssd vccd vccd output1035/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output641_A output641/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[81\]_B la_buf_enable\[81\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__450__A _450_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output739_A output739/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output906_A output906/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[14\]_A user_to_mprj_in_gates\[14\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[22\]_A input564/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[117\]_A _581_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__625__A _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[104\]_B user_to_mprj_in_gates\[104\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[54\]_A _518_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[72\]_B la_buf_enable\[72\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput652 output652/A vssd vssd vccd vccd la_data_in_core[122] sky130_fd_sc_hd__buf_2
Xoutput641 output641/A vssd vssd vccd vccd la_data_in_core[112] sky130_fd_sc_hd__buf_2
Xoutput630 output630/A vssd vssd vccd vccd la_data_in_core[102] sky130_fd_sc_hd__buf_2
Xoutput663 output663/A vssd vssd vccd vccd la_data_in_core[17] sky130_fd_sc_hd__buf_2
XANTENNA__360__A _360_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_wb_ena_buf_A input614/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput696 output696/A vssd vssd vccd vccd la_data_in_core[47] sky130_fd_sc_hd__buf_2
Xoutput674 output674/A vssd vssd vccd vccd la_data_in_core[27] sky130_fd_sc_hd__buf_2
Xoutput685 output685/A vssd vssd vccd vccd la_data_in_core[37] sky130_fd_sc_hd__buf_2
XANTENNA_mprj_stb_buf_A _394_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output1003_A output1003/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[46\] input328/X mprj_logic_high_inst/HI[376] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[46\]/B sky130_fd_sc_hd__and2_1
XTAP_2015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[13\]_A input554/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[119\]_A user_to_mprj_in_gates\[119\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_33 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[108\]_A _572_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__535__A _535_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[24\] _616_/A la_buf_enable\[24\]/B vssd vssd vccd vccd la_buf\[24\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_22_170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[45\]_A _509_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input372_A la_iena_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input66_A la_data_out_core[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[63\]_B la_buf_enable\[63\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_708 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_508_ _508_/A vssd vssd vccd vccd _508_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output689_A output689/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_439_ _439_/A vssd vssd vccd vccd _439_/Y sky130_fd_sc_hd__inv_4
XANTENNA__445__A _445_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output856_A output856/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[36\]_A _500_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[54\]_B la_buf_enable\[54\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[121\]_A _384_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[126\]_B mprj_logic_high_inst/HI[456] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1044 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_788 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[12\]_TE la_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__355__A _355_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[27\]_A _491_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[45\]_B la_buf_enable\[45\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1120_A output1120/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_7 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[112\]_A _375_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[117\]_B mprj_logic_high_inst/HI[447] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input120_A la_data_out_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input218_A la_data_out_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input587_A mprj_dat_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[18\]_A _482_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[1\] input561/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[1\]/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_7_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[101\] input262/X mprj_logic_high_inst/HI[431] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[101\]/B sky130_fd_sc_hd__and2_1
XANTENNA_la_buf_enable\[36\]_B la_buf_enable\[36\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[5\]_A input343/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[103\]_A _366_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[107\] user_to_mprj_in_gates\[107\]/Y vssd vssd vccd vccd
+ output763/A sky130_fd_sc_hd__clkinv_4
XFILLER_26_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[108\]_B mprj_logic_high_inst/HI[438] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_38_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[73\] user_to_mprj_in_gates\[73\]/Y vssd vssd vccd vccd output853/A
+ sky130_fd_sc_hd__inv_2
XFILLER_4_1331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[35\]_TE la_buf\[35\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output973_A output973/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[31\] input574/X repeater1125/X vssd vssd vccd vccd user_wb_dat_gates\[31\]/Y
+ sky130_fd_sc_hd__nand2_8
XFILLER_33_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[27\]_B la_buf_enable\[27\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput1110 output1110/A vssd vssd vccd vccd mprj_sel_o_user[1] sky130_fd_sc_hd__buf_2
XFILLER_44_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput1121 output1121/A vssd vssd vccd vccd user_irq[0] sky130_fd_sc_hd__buf_2
XFILLER_0_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[6\] _438_/Y mprj_dat_buf\[6\]/TE vssd vssd vccd vccd output1105/A sky130_fd_sc_hd__einvp_8
XFILLER_9_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1242 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[96\]_A _359_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_736 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[30\]_B mprj_logic_high_inst/HI[360] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[3\]_TE la_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1070_A output1070/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[18\]_B la_buf_enable\[18\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input168_A la_data_out_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[20\]_A _612_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[91\] _354_/A la_buf_enable\[91\]/B vssd vssd vccd vccd la_buf\[91\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_47_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[97\]_B mprj_logic_high_inst/HI[427] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[58\]_TE la_buf\[58\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input335_A la_iena_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input29_A la_data_out_core[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[77\] _541_/Y la_buf\[77\]/TE vssd vssd vccd vccd output729/A sky130_fd_sc_hd__einvp_4
XANTENNA_input502_A la_oenb_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[87\]_A _350_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[21\]_B mprj_logic_high_inst/HI[351] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output721_A output721/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[11\]_A _603_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output819_A output819/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[88\]_B mprj_logic_high_inst/HI[418] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[66\] input94/X user_to_mprj_in_gates\[66\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[66\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[78\]_A _341_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[12\]_B mprj_logic_high_inst/HI[342] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__633__A _633_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[5\]_A input577/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[79\]_B mprj_logic_high_inst/HI[409] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[5\]_A input87/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[69\]_A _332_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[124\]_A_N _387_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_382 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__543__A _543_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input285_A la_iena_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input452_A la_oenb_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput530 mprj_adr_o_core[21] vssd vssd vccd vccd _421_/A sky130_fd_sc_hd__buf_2
Xinput563 mprj_dat_i_user[21] vssd vssd vccd vccd input563/X sky130_fd_sc_hd__buf_8
Xinput552 mprj_dat_i_user[11] vssd vssd vccd vccd input552/X sky130_fd_sc_hd__buf_12
Xinput541 mprj_adr_o_core[31] vssd vssd vccd vccd _431_/A sky130_fd_sc_hd__buf_2
Xinput574 mprj_dat_i_user[31] vssd vssd vccd vccd input574/X sky130_fd_sc_hd__clkbuf_2
Xinput585 mprj_dat_o_core[12] vssd vssd vccd vccd _444_/A sky130_fd_sc_hd__buf_2
Xinput596 mprj_dat_o_core[22] vssd vssd vccd vccd _454_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[9\]_TE mprj_logic_high_inst/HI[211] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[36\] user_to_mprj_in_gates\[36\]/Y vssd vssd vccd vccd output812/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output671_A output671/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__453__A _453_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output769_A output769/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output936_A output936/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__628__A _628_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__363__A _363_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1033_A output1033/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[76\] input361/X mprj_logic_high_inst/HI[406] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[76\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[102\] _365_/Y mprj_logic_high_inst/HI[304] vssd vssd vccd
+ vccd output886/A sky130_fd_sc_hd__einvp_2
XFILLER_44_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_610_ _610_/A vssd vssd vccd vccd _610_/Y sky130_fd_sc_hd__inv_2
X_541_ _541_/A vssd vssd vccd vccd _541_/Y sky130_fd_sc_hd__inv_2
XANTENNA__538__A _538_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[32\] _624_/Y mprj_logic_high_inst/HI[234] vssd vssd vccd
+ vccd output936/A sky130_fd_sc_hd__einvp_8
XFILLER_17_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[54\] _646_/A la_buf_enable\[54\]/B vssd vssd vccd vccd la_buf\[54\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_38_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_472_ _472_/A vssd vssd vccd vccd _472_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input200_A la_data_out_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[20\]_A _452_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input96_A la_data_out_core[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xrepeater1125 repeater1125/A vssd vssd vccd vccd repeater1125/X sky130_fd_sc_hd__buf_12
XFILLER_5_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput360 la_iena_mprj[75] vssd vssd vccd vccd input360/X sky130_fd_sc_hd__clkbuf_1
Xinput371 la_iena_mprj[85] vssd vssd vccd vccd input371/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__448__A _448_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput382 la_iena_mprj[95] vssd vssd vccd vccd input382/X sky130_fd_sc_hd__clkbuf_1
Xinput393 la_oenb_mprj[104] vssd vssd vccd vccd _367_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output886_A output886/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[11\]_A _443_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[29\] input53/X user_to_mprj_in_gates\[29\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[29\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_16_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[30\]_TE mprj_logic_high_inst/HI[232] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xoutput801 output801/A vssd vssd vccd vccd la_data_in_mprj[26] sky130_fd_sc_hd__buf_2
Xoutput812 output812/A vssd vssd vccd vccd la_data_in_mprj[36] sky130_fd_sc_hd__buf_2
XANTENNA_mprj_adr_buf\[29\]_A _429_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput834 output834/A vssd vssd vccd vccd la_data_in_mprj[56] sky130_fd_sc_hd__buf_2
XFILLER_6_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput823 output823/A vssd vssd vccd vccd la_data_in_mprj[46] sky130_fd_sc_hd__buf_2
Xoutput845 output845/A vssd vssd vccd vccd la_data_in_mprj[66] sky130_fd_sc_hd__buf_2
XFILLER_47_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput856 output856/A vssd vssd vccd vccd la_data_in_mprj[76] sky130_fd_sc_hd__buf_2
Xoutput867 output867/A vssd vssd vccd vccd la_data_in_mprj[86] sky130_fd_sc_hd__buf_2
Xoutput878 output878/A vssd vssd vccd vccd la_data_in_mprj[96] sky130_fd_sc_hd__buf_2
Xoutput889 output889/A vssd vssd vccd vccd la_oenb_core[105] sky130_fd_sc_hd__buf_2
XFILLER_28_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__358__A _358_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[6\]_A _598_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[106\]_TE la_buf\[106\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[5\]_TE mprj_adr_buf\[5\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[28\] _460_/Y mprj_dat_buf\[28\]/TE vssd vssd vccd vccd output1097/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_2_768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input150_A la_data_out_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input248_A la_data_out_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1716 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input415_A la_oenb_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input11_A la_data_out_core[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[31\]_B repeater1125/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_524_ _524_/A vssd vssd vccd vccd _524_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_455_ _455_/A vssd vssd vccd vccd _455_/Y sky130_fd_sc_hd__inv_4
XFILLER_26_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[53\]_TE mprj_logic_high_inst/HI[255] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_386_ _386_/A vssd vssd vccd vccd _386_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[23\] _423_/Y mprj_adr_buf\[23\]/TE vssd vssd vccd vccd output1027/A
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[9\]_TE mprj_dat_buf\[9\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output634_A output634/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output801_A output801/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput190 la_data_out_mprj[37] vssd vssd vccd vccd _501_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[22\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[8\] _600_/A la_buf_enable\[8\]/B vssd vssd vccd vccd la_buf\[8\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_18_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__641__A _641_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput653 output653/A vssd vssd vccd vccd la_data_in_core[123] sky130_fd_sc_hd__buf_2
Xoutput642 output642/A vssd vssd vccd vccd la_data_in_core[113] sky130_fd_sc_hd__buf_2
Xoutput631 output631/A vssd vssd vccd vccd la_data_in_core[103] sky130_fd_sc_hd__buf_2
XFILLER_47_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_wb_ena_buf_B user_to_mprj_wb_ena_buf/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput697 output697/A vssd vssd vccd vccd la_data_in_core[48] sky130_fd_sc_hd__buf_2
Xoutput686 output686/A vssd vssd vccd vccd la_data_in_core[38] sky130_fd_sc_hd__buf_2
Xoutput675 output675/A vssd vssd vccd vccd la_data_in_core[28] sky130_fd_sc_hd__buf_2
Xoutput664 output664/A vssd vssd vccd vccd la_data_in_core[18] sky130_fd_sc_hd__buf_2
XFILLER_28_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input3_A caravel_rstn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[82\]_A_N _345_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[91\]_TE la_buf\[91\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1828 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[13\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[76\]_TE mprj_logic_high_inst/HI[278] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[39\] input320/X mprj_logic_high_inst/HI[369] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[39\]/B sky130_fd_sc_hd__and2_1
XTAP_1348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[97\]_A_N _360_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_23 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[20\]_A_N _612_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[17\] _609_/A la_buf_enable\[17\]/B vssd vssd vccd vccd la_buf\[17\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_10_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input198_A la_data_out_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_878 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__551__A _551_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[35\]_A_N _627_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input365_A la_iena_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input59_A la_data_out_core[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_irq_gates\[0\] input621/X user_irq_gates\[0\]/B vssd vssd vccd vccd user_irq_gates\[0\]/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_2_510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input532_A mprj_adr_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[122\] _385_/A la_buf_enable\[122\]/B vssd vssd vccd vccd la_buf\[122\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_4_2225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_507_ _507_/A vssd vssd vccd vccd _507_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_438_ _438_/A vssd vssd vccd vccd _438_/Y sky130_fd_sc_hd__inv_4
X_369_ _369_/A vssd vssd vccd vccd _369_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output751_A output751/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__461__A _461_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output849_A output849/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[96\] input127/X user_to_mprj_in_gates\[96\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[96\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_1964 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[99\]_TE mprj_logic_high_inst/HI[301] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1056 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__636__A _636_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[5\]_A _405_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__371__A _371_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1113_A output1113/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input113_A la_data_out_core[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__546__A _546_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input482_A la_oenb_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[22\] _486_/Y la_buf\[22\]/TE vssd vssd vccd vccd output669/A sky130_fd_sc_hd__einvp_8
XFILLER_32_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[5\]_B mprj_logic_high_inst/HI[335] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_stb_buf_TE mprj_stb_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[66\] user_to_mprj_in_gates\[66\]/Y vssd vssd vccd vccd output845/A
+ sky130_fd_sc_hd__inv_2
XFILLER_37_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__456__A _456_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output799_A output799/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output966_A output966/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[24\] input566/X repeater1125/X vssd vssd vccd vccd user_wb_dat_gates\[24\]/Y
+ sky130_fd_sc_hd__nand2_8
XTAP_1690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[11\] input26/X user_to_mprj_in_gates\[11\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[11\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_buffers\[21\] user_wb_dat_gates\[21\]/Y vssd vssd vccd vccd output1058/A
+ sky130_fd_sc_hd__clkinv_8
Xoutput1100 output1100/A vssd vssd vccd vccd mprj_dat_o_user[30] sky130_fd_sc_hd__buf_2
Xoutput1111 output1111/A vssd vssd vccd vccd mprj_sel_o_user[2] sky130_fd_sc_hd__buf_2
Xoutput1122 output1122/A vssd vssd vccd vccd user_irq[1] sky130_fd_sc_hd__buf_2
XFILLER_44_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[126\]_B la_buf_enable\[126\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[122\] input29/X user_to_mprj_in_gates\[122\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[122\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__366__A _366_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[95\]_A input126/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output1063_A output1063/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[31\]_TE mprj_adr_buf\[31\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[62\] _654_/Y mprj_logic_high_inst/HI[264] vssd vssd vccd
+ vccd output969/A sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[84\] _347_/A la_buf_enable\[84\]/B vssd vssd vccd vccd la_buf\[84\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_27_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[117\]_B la_buf_enable\[117\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[10\] _442_/Y mprj_dat_buf\[10\]/TE vssd vssd vccd vccd output1078/A
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input230_A la_data_out_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input328_A la_iena_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_buffers\[8\]_A user_wb_dat_gates\[8\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[86\]_A input116/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[126\] _590_/Y la_buf\[126\]/TE vssd vssd vccd vccd output656/A sky130_fd_sc_hd__einvp_2
XFILLER_32_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output714_A output714/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[108\]_B la_buf_enable\[108\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[10\]_A input15/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[59\] input86/X user_to_mprj_in_gates\[59\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[59\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_A input106/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[5\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[5\]_B user_to_mprj_in_gates\[5\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[21\] input301/X mprj_logic_high_inst/HI[351] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[21\]/B sky130_fd_sc_hd__and2_1
XFILLER_52_372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[68\]_A input96/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[25\]_TE la_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input180_A la_data_out_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input278_A la_iena_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input41_A la_data_out_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input445_A la_oenb_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput520 mprj_adr_o_core[12] vssd vssd vccd vccd _412_/A sky130_fd_sc_hd__clkbuf_2
Xinput564 mprj_dat_i_user[22] vssd vssd vccd vccd input564/X sky130_fd_sc_hd__buf_8
Xinput553 mprj_dat_i_user[12] vssd vssd vccd vccd input553/X sky130_fd_sc_hd__buf_12
XFILLER_48_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput542 mprj_adr_o_core[3] vssd vssd vccd vccd _403_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input612_A mprj_dat_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput531 mprj_adr_o_core[22] vssd vssd vccd vccd _422_/A sky130_fd_sc_hd__clkbuf_2
Xinput575 mprj_dat_i_user[3] vssd vssd vccd vccd input575/X sky130_fd_sc_hd__buf_8
XFILLER_1_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput586 mprj_dat_o_core[13] vssd vssd vccd vccd _445_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput597 mprj_dat_o_core[23] vssd vssd vccd vccd _455_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[59\]_A input86/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[29\] user_to_mprj_in_gates\[29\]/Y vssd vssd vccd vccd output804/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output664_A output664/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output831_A output831/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output929_A output929/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_634 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[9\]_A user_to_mprj_in_gates\[9\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__644__A _644_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1746 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[48\]_TE la_buf\[48\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output1026_A output1026/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[69\] input353/X mprj_logic_high_inst/HI[399] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[69\]/B sky130_fd_sc_hd__and2_1
XFILLER_40_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_540_ _540_/A vssd vssd vccd vccd _540_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[25\] _617_/Y mprj_logic_high_inst/HI[227] vssd vssd vccd
+ vccd output928/A sky130_fd_sc_hd__einvp_2
Xla_buf_enable\[47\] _639_/A la_buf_enable\[47\]/B vssd vssd vccd vccd la_buf\[47\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_32_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[7\] _599_/Y mprj_logic_high_inst/HI[209] vssd vssd vccd
+ vccd output988/A sky130_fd_sc_hd__einvp_2
XFILLER_25_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_471_ _471_/A vssd vssd vccd vccd _471_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[125\]_A input32/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__554__A _554_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input395_A la_oenb_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input89_A la_data_out_core[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input562_A mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[0\] _464_/Y la_buf\[0\]/TE vssd vssd vccd vccd output627/A sky130_fd_sc_hd__einvp_8
XFILLER_4_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput350 la_iena_mprj[66] vssd vssd vccd vccd input350/X sky130_fd_sc_hd__clkbuf_1
Xinput361 la_iena_mprj[76] vssd vssd vccd vccd input361/X sky130_fd_sc_hd__clkbuf_1
Xinput372 la_iena_mprj[86] vssd vssd vccd vccd input372/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput383 la_iena_mprj[96] vssd vssd vccd vccd input383/X sky130_fd_sc_hd__clkbuf_1
Xinput394 la_oenb_mprj[105] vssd vssd vccd vccd _368_/A sky130_fd_sc_hd__buf_2
XFILLER_35_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__464__A _464_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_A input22/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output879_A output879/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output781_A output781/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput802 output802/A vssd vssd vccd vccd la_data_in_mprj[27] sky130_fd_sc_hd__buf_2
Xoutput835 output835/A vssd vssd vccd vccd la_data_in_mprj[57] sky130_fd_sc_hd__buf_2
Xoutput824 output824/A vssd vssd vccd vccd la_data_in_mprj[47] sky130_fd_sc_hd__buf_2
Xoutput813 output813/A vssd vssd vccd vccd la_data_in_mprj[37] sky130_fd_sc_hd__buf_2
Xoutput846 output846/A vssd vssd vccd vccd la_data_in_mprj[67] sky130_fd_sc_hd__buf_2
XANTENNA_la_buf_enable\[123\]_A_N _386_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput857 output857/A vssd vssd vccd vccd la_data_in_mprj[77] sky130_fd_sc_hd__buf_2
Xoutput868 output868/A vssd vssd vccd vccd la_data_in_mprj[87] sky130_fd_sc_hd__buf_2
Xoutput879 output879/A vssd vssd vccd vccd la_data_in_mprj[97] sky130_fd_sc_hd__buf_2
XTAP_320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__639__A _639_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__374__A _374_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[107\]_A input12/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input143_A la_data_out_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__549__A _549_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input310_A la_iena_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input408_A la_oenb_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_523_ _523_/A vssd vssd vccd vccd _523_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_454_ _454_/A vssd vssd vccd vccd _454_/Y sky130_fd_sc_hd__inv_4
Xla_buf\[52\] _516_/Y la_buf\[52\]/TE vssd vssd vccd vccd output702/A sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[124\] input287/X mprj_logic_high_inst/HI[454] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[124\]/B sky130_fd_sc_hd__and2_1
XFILLER_13_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_385_ _385_/A vssd vssd vccd vccd _385_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[16\] _416_/Y mprj_adr_buf\[16\]/TE vssd vssd vccd vccd output1019/A
+ sky130_fd_sc_hd__einvp_4
XFILLER_5_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output627_A output627/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[96\] user_to_mprj_in_gates\[96\]/Y vssd vssd vccd vccd output878/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_42_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__459__A _459_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_rstn_buf input3/X mprj_rstn_buf/TE vssd vssd vccd vccd output1124/A sky130_fd_sc_hd__einvp_2
Xinput180 la_data_out_mprj[28] vssd vssd vccd vccd _492_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput191 la_data_out_mprj[38] vssd vssd vccd vccd _502_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_output996_A output996/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[41\] input67/X user_to_mprj_in_gates\[41\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[41\]/Y sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_buffers\[6\] user_wb_dat_gates\[6\]/Y vssd vssd vccd vccd output1073/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_36_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[5\]_B la_buf_enable\[5\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput654 output654/A vssd vssd vccd vccd la_data_in_core[124] sky130_fd_sc_hd__buf_2
Xoutput643 output643/A vssd vssd vccd vccd la_data_in_core[114] sky130_fd_sc_hd__buf_2
Xoutput632 output632/A vssd vssd vccd vccd la_data_in_core[104] sky130_fd_sc_hd__buf_2
XFILLER_47_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput687 output687/A vssd vssd vccd vccd la_data_in_core[39] sky130_fd_sc_hd__buf_2
Xoutput676 output676/A vssd vssd vccd vccd la_data_in_core[29] sky130_fd_sc_hd__buf_2
Xoutput665 output665/A vssd vssd vccd vccd la_data_in_core[19] sky130_fd_sc_hd__buf_2
XFILLER_28_1033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[3\] input65/X user_to_mprj_in_gates\[3\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[3\]/Y sky130_fd_sc_hd__nand2_1
Xoutput698 output698/A vssd vssd vccd vccd la_data_in_core[49] sky130_fd_sc_hd__buf_2
XFILLER_28_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1954 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__369__A _369_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[121\]_TE mprj_logic_high_inst/HI[323] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1093_A output1093/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[60\]_A input344/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[92\] _355_/Y mprj_logic_high_inst/HI[294] vssd vssd vccd
+ vccd output1002/A sky130_fd_sc_hd__einvp_4
XANTENNA_input260_A la_iena_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input358_A la_iena_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[5\] input343/X mprj_logic_high_inst/HI[335] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[5\]/B sky130_fd_sc_hd__and2_1
XANTENNA_input525_A mprj_adr_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[115\] _378_/A la_buf_enable\[115\]/B vssd vssd vccd vccd la_buf\[115\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_oen_buffers\[20\]_TE mprj_logic_high_inst/HI[222] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_506_ _506_/A vssd vssd vccd vccd _506_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_33_415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[51\]_A input334/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_437_ _437_/A vssd vssd vccd vccd _437_/Y sky130_fd_sc_hd__inv_4
XFILLER_20_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_368_ _368_/A vssd vssd vccd vccd _368_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[11\] user_to_mprj_in_gates\[11\]/Y vssd vssd vccd vccd output777/A
+ sky130_fd_sc_hd__inv_6
XANTENNA_output744_A output744/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output911_A output911/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[89\] input119/X user_to_mprj_in_gates\[89\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[89\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[42\]_A input324/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__652__A _652_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[43\]_TE mprj_logic_high_inst/HI[245] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1106_A output1106/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[51\] input334/X mprj_logic_high_inst/HI[381] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[51\]/B sky130_fd_sc_hd__and2_1
XFILLER_5_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_cyc_buf _393_/Y mprj_cyc_buf/TE vssd vssd vccd vccd output1044/A sky130_fd_sc_hd__einvp_8
XTAP_1113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input106_A la_data_out_core[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[33\]_A input314/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[3\] user_to_mprj_in_gates\[3\]/Y vssd vssd vccd vccd output816/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_42_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__562__A _562_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input475_A la_oenb_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input71_A la_data_out_core[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[119\]_TE la_buf\[119\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[15\] _479_/Y la_buf\[15\]/TE vssd vssd vccd vccd output661/A sky130_fd_sc_hd__einvp_8
XFILLER_32_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[0\]_A _432_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[8\] _408_/Y mprj_adr_buf\[8\]/TE vssd vssd vccd vccd output1042/A sky130_fd_sc_hd__einvp_4
XFILLER_4_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[24\]_A input304/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[59\] user_to_mprj_in_gates\[59\]/Y vssd vssd vccd vccd output837/A
+ sky130_fd_sc_hd__inv_2
XANTENNA_output694_A output694/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output959_A output959/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__472__A _472_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output861_A output861/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[17\] input558/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[17\]/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_50_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[81\]_A_N _344_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[81\]_TE la_buf\[81\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput1101 output1101/A vssd vssd vccd vccd mprj_dat_o_user[31] sky130_fd_sc_hd__buf_2
Xoutput1112 output1112/A vssd vssd vccd vccd mprj_sel_o_user[3] sky130_fd_sc_hd__buf_2
XFILLER_44_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_buffers\[14\] user_wb_dat_gates\[14\]/Y vssd vssd vccd vccd output1050/A
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_user_to_mprj_oen_buffers\[66\]_TE mprj_logic_high_inst/HI[268] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xoutput1123 output1123/A vssd vssd vccd vccd user_irq[2] sky130_fd_sc_hd__buf_2
XANTENNA_la_buf_enable\[96\]_A_N _359_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[115\] input21/X user_to_mprj_in_gates\[115\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[115\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA__647__A _647_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_540 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[34\]_A_N _626_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[15\]_A input294/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[95\]_B user_to_mprj_in_gates\[95\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[49\]_A_N _641_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__382__A _382_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output1056_A output1056/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_clk2_buf_TE mprj_clk2_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[99\] input386/X mprj_logic_high_inst/HI[429] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[99\]/B sky130_fd_sc_hd__and2_1
XFILLER_3_105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[125\] _388_/Y mprj_logic_high_inst/HI[327] vssd vssd vccd
+ vccd output911/A sky130_fd_sc_hd__einvp_4
XANTENNA_mprj_dat_buf\[30\]_TE mprj_dat_buf\[30\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[55\] _647_/Y mprj_logic_high_inst/HI[257] vssd vssd vccd
+ vccd output961/A sky130_fd_sc_hd__einvp_4
XFILLER_27_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[80\]_A user_to_mprj_in_gates\[80\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_48_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[77\] _340_/A la_buf_enable\[77\]/B vssd vssd vccd vccd la_buf\[77\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_input223_A la_data_out_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_ena_buf\[2\]_A input626/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__557__A _557_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[86\]_B user_to_mprj_in_gates\[86\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_input592_A mprj_dat_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[89\]_TE mprj_logic_high_inst/HI[291] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[119\] _583_/Y la_buf\[119\]/TE vssd vssd vccd vccd output648/A sky130_fd_sc_hd__einvp_2
XFILLER_10_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[112\] user_to_mprj_in_gates\[112\]/Y vssd vssd vccd vccd
+ output769/A sky130_fd_sc_hd__clkinv_4
XTAP_749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[10\]_B user_to_mprj_in_gates\[10\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[71\]_A user_to_mprj_in_gates\[71\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output707_A output707/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__467__A _467_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_B user_to_mprj_in_gates\[77\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[62\]_A user_to_mprj_in_gates\[62\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__377__A _377_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[14\] input293/X mprj_logic_high_inst/HI[344] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[14\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[68\]_B user_to_mprj_in_gates\[68\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input173_A la_data_out_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[100\]_A user_to_mprj_in_gates\[100\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input340_A la_iena_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input438_A la_oenb_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput510 la_oenb_mprj[95] vssd vssd vccd vccd _358_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_buffers\[53\]_A user_to_mprj_in_gates\[53\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xinput521 mprj_adr_o_core[13] vssd vssd vccd vccd _413_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input34_A la_data_out_core[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput554 mprj_dat_i_user[13] vssd vssd vccd vccd input554/X sky130_fd_sc_hd__buf_12
XFILLER_48_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput543 mprj_adr_o_core[4] vssd vssd vccd vccd _404_/A sky130_fd_sc_hd__buf_12
Xinput532 mprj_adr_o_core[23] vssd vssd vccd vccd _423_/A sky130_fd_sc_hd__clkbuf_2
Xinput565 mprj_dat_i_user[23] vssd vssd vccd vccd input565/X sky130_fd_sc_hd__buf_6
Xinput576 mprj_dat_i_user[4] vssd vssd vccd vccd input576/X sky130_fd_sc_hd__clkbuf_16
XFILLER_48_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[82\] _546_/Y la_buf\[82\]/TE vssd vssd vccd vccd output735/A sky130_fd_sc_hd__einvp_4
Xinput587 mprj_dat_o_core[14] vssd vssd vccd vccd _446_/A sky130_fd_sc_hd__clkbuf_2
Xinput598 mprj_dat_o_core[24] vssd vssd vccd vccd _456_/A sky130_fd_sc_hd__buf_2
XANTENNA_input605_A mprj_dat_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_B user_to_mprj_in_gates\[59\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[93\]_A _557_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output657_A output657/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output824_A output824/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[44\]_A user_to_mprj_in_gates\[44\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[71\] input100/X user_to_mprj_in_gates\[71\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[71\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[21\]_TE mprj_adr_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[84\]_A _548_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1878 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[35\]_A user_to_mprj_in_gates\[35\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1019_A output1019/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_470_ _470_/A vssd vssd vccd vccd _470_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[18\] _610_/Y mprj_logic_high_inst/HI[220] vssd vssd vccd
+ vccd output920/A sky130_fd_sc_hd__einvp_2
XFILLER_41_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[125\]_B user_to_mprj_in_gates\[125\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[75\]_A _539_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_590 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input388_A la_oenb_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input290_A la_iena_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[93\]_B la_buf_enable\[93\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input555_A mprj_dat_i_user[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__570__A _570_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1716 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_82 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[26\]_A user_to_mprj_in_gates\[26\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput340 la_iena_mprj[57] vssd vssd vccd vccd input340/X sky130_fd_sc_hd__clkbuf_1
Xinput351 la_iena_mprj[67] vssd vssd vccd vccd input351/X sky130_fd_sc_hd__clkbuf_1
Xinput362 la_iena_mprj[77] vssd vssd vccd vccd input362/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput373 la_iena_mprj[87] vssd vssd vccd vccd input373/X sky130_fd_sc_hd__clkbuf_1
Xinput384 la_iena_mprj[97] vssd vssd vccd vccd input384/X sky130_fd_sc_hd__clkbuf_1
Xinput395 la_oenb_mprj[106] vssd vssd vccd vccd _369_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_599_ _599_/A vssd vssd vccd vccd _599_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[41\] user_to_mprj_in_gates\[41\]/Y vssd vssd vccd vccd output818/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_in_gates\[116\]_B user_to_mprj_in_gates\[116\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[66\]_A _530_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output774_A output774/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output941_A output941/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[84\]_B la_buf_enable\[84\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__480__A _480_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput803 output803/A vssd vssd vccd vccd la_data_in_mprj[28] sky130_fd_sc_hd__buf_2
XFILLER_47_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput825 output825/A vssd vssd vccd vccd la_data_in_mprj[48] sky130_fd_sc_hd__buf_2
Xoutput814 output814/A vssd vssd vccd vccd la_data_in_mprj[38] sky130_fd_sc_hd__buf_2
Xoutput836 output836/A vssd vssd vccd vccd la_data_in_mprj[58] sky130_fd_sc_hd__buf_2
XFILLER_47_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput847 output847/A vssd vssd vccd vccd la_data_in_mprj[68] sky130_fd_sc_hd__buf_2
Xoutput858 output858/A vssd vssd vccd vccd la_data_in_mprj[78] sky130_fd_sc_hd__buf_2
Xoutput869 output869/A vssd vssd vccd vccd la_data_in_mprj[88] sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_buffers\[17\]_A user_to_mprj_in_gates\[17\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[25\]_A input567/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[15\]_TE la_buf\[15\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__655__A _655_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[107\]_B user_to_mprj_in_gates\[107\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[57\]_A _521_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[75\]_B la_buf_enable\[75\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__390__A _390_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[81\] input367/X mprj_logic_high_inst/HI[411] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[81\]/B sky130_fd_sc_hd__and2_1
XFILLER_24_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[16\]_A input557/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input136_A la_data_out_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_522_ _522_/A vssd vssd vccd vccd _522_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input303_A la_iena_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_453_ _453_/A vssd vssd vccd vccd _453_/Y sky130_fd_sc_hd__inv_6
XFILLER_32_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__565__A _565_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_384_ _384_/A vssd vssd vccd vccd _384_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[45\] _509_/Y la_buf\[45\]/TE vssd vssd vccd vccd output694/A sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[48\]_A _512_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[117\] input279/X mprj_logic_high_inst/HI[447] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[117\]/B sky130_fd_sc_hd__and2_1
XFILLER_13_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[66\]_B la_buf_enable\[66\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[101\] _565_/Y la_buf\[101\]/TE vssd vssd vccd vccd output629/A sky130_fd_sc_hd__einvp_4
XFILLER_9_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput170 la_data_out_mprj[19] vssd vssd vccd vccd _483_/A sky130_fd_sc_hd__clkbuf_2
Xinput181 la_data_out_mprj[29] vssd vssd vccd vccd _493_/A sky130_fd_sc_hd__clkbuf_2
Xuser_to_mprj_in_buffers\[89\] user_to_mprj_in_gates\[89\]/Y vssd vssd vccd vccd output870/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_7_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[38\]_TE la_buf\[38\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput192 la_data_out_mprj[39] vssd vssd vccd vccd _503_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_output989_A output989/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output891_A output891/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__475__A _475_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[34\] input59/X user_to_mprj_in_gates\[34\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[34\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[39\]_A _503_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[57\]_B la_buf_enable\[57\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput644 output644/A vssd vssd vccd vccd la_data_in_core[115] sky130_fd_sc_hd__buf_2
Xoutput633 output633/A vssd vssd vccd vccd la_data_in_core[105] sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_oen_buffers\[124\]_A _387_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput655 output655/A vssd vssd vccd vccd la_data_in_core[125] sky130_fd_sc_hd__buf_2
Xoutput688 output688/A vssd vssd vccd vccd la_data_in_core[3] sky130_fd_sc_hd__buf_2
Xoutput677 output677/A vssd vssd vccd vccd la_data_in_core[2] sky130_fd_sc_hd__buf_2
Xoutput666 output666/A vssd vssd vccd vccd la_data_in_core[1] sky130_fd_sc_hd__buf_2
Xoutput699 output699/A vssd vssd vccd vccd la_data_in_core[4] sky130_fd_sc_hd__buf_2
XFILLER_47_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__385__A _385_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_14 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[60\]_B mprj_logic_high_inst/HI[390] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output1086_A output1086/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[6\]_TE la_buf\[6\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[48\]_B la_buf_enable\[48\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[115\]_A _378_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[85\] _348_/Y mprj_logic_high_inst/HI[287] vssd vssd vccd
+ vccd output994/A sky130_fd_sc_hd__einvp_2
XANTENNA_user_to_mprj_oen_buffers\[50\]_A _642_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input253_A la_data_out_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_578 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input420_A la_oenb_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input518_A mprj_adr_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[108\] _371_/A la_buf_enable\[108\]/B vssd vssd vccd vccd la_buf\[108\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_46_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_505_ _505_/A vssd vssd vccd vccd _505_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[51\]_B mprj_logic_high_inst/HI[381] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_436_ _436_/A vssd vssd vccd vccd _436_/Y sky130_fd_sc_hd__inv_4
XANTENNA_la_buf_enable\[122\]_A_N _385_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_367_ _367_/A vssd vssd vccd vccd _367_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[39\]_B la_buf_enable\[39\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[8\]_A input376/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[41\]_A _633_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[106\]_A _369_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output737_A output737/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output904_A output904/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[42\]_B mprj_logic_high_inst/HI[372] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_51_257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[32\]_A _624_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1001_A output1001/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[99\]_A _362_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[44\] input326/X mprj_logic_high_inst/HI[374] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[44\]/B sky130_fd_sc_hd__and2_1
XFILLER_5_1879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[33\]_B mprj_logic_high_inst/HI[363] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_1169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[22\] _614_/A la_buf_enable\[22\]/B vssd vssd vccd vccd la_buf\[22\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_23_482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input468_A la_oenb_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input370_A la_iena_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input64_A la_data_out_core[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[23\]_A _615_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[24\]_B mprj_logic_high_inst/HI[354] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output687_A output687/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_419_ _419_/A vssd vssd vccd vccd _419_/Y sky130_fd_sc_hd__inv_8
XFILLER_14_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output854_A output854/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[111\]_TE mprj_logic_high_inst/HI[313] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[14\]_A _606_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput1102 output1102/A vssd vssd vccd vccd mprj_dat_o_user[3] sky130_fd_sc_hd__buf_2
Xoutput1113 output1113/A vssd vssd vccd vccd mprj_stb_o_user sky130_fd_sc_hd__buf_2
Xoutput1124 output1124/A vssd vssd vccd vccd user_reset sky130_fd_sc_hd__buf_2
XFILLER_44_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[108\] input13/X user_to_mprj_in_gates\[108\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[108\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[10\]_A _410_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[15\]_B mprj_logic_high_inst/HI[345] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_52_566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[8\]_A input580/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[10\]_TE mprj_logic_high_inst/HI[212] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output1049_A output1049/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[118\] _381_/Y mprj_logic_high_inst/HI[320] vssd vssd vccd
+ vccd output903/A sky130_fd_sc_hd__einvp_2
XFILLER_5_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[8\]_A input120/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[48\] _640_/Y mprj_logic_high_inst/HI[250] vssd vssd vccd
+ vccd output953/A sky130_fd_sc_hd__einvp_2
XFILLER_28_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[2\]_B user_irq_ena_buf\[2\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input216_A la_data_out_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__573__A _573_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input585_A mprj_dat_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[105\] user_to_mprj_in_gates\[105\]/Y vssd vssd vccd vccd
+ output761/A sky130_fd_sc_hd__clkinv_4
XFILLER_43_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[71\] user_to_mprj_in_gates\[71\]/Y vssd vssd vccd vccd output851/A
+ sky130_fd_sc_hd__inv_2
XFILLER_47_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output971_A output971/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__483__A _483_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[33\]_TE mprj_logic_high_inst/HI[235] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[4\] _436_/Y mprj_dat_buf\[4\]/TE vssd vssd vccd vccd output1103/A sky130_fd_sc_hd__einvp_8
XFILLER_29_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[109\]_TE la_buf\[109\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__393__A _393_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[8\]_TE mprj_adr_buf\[8\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input166_A la_data_out_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput500 la_oenb_mprj[86] vssd vssd vccd vccd _349_/A sky130_fd_sc_hd__clkbuf_4
Xinput511 la_oenb_mprj[96] vssd vssd vccd vccd _359_/A sky130_fd_sc_hd__clkbuf_4
Xinput555 mprj_dat_i_user[14] vssd vssd vccd vccd input555/X sky130_fd_sc_hd__buf_12
XFILLER_48_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2080 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__568__A _568_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input333_A la_iena_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput544 mprj_adr_o_core[5] vssd vssd vccd vccd _405_/A sky130_fd_sc_hd__clkbuf_4
Xinput522 mprj_adr_o_core[14] vssd vssd vccd vccd _414_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput533 mprj_adr_o_core[24] vssd vssd vccd vccd _424_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input27_A la_data_out_core[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput566 mprj_dat_i_user[24] vssd vssd vccd vccd input566/X sky130_fd_sc_hd__buf_2
Xinput577 mprj_dat_i_user[5] vssd vssd vccd vccd input577/X sky130_fd_sc_hd__buf_12
XFILLER_48_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[80\]_A_N _343_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput588 mprj_dat_o_core[15] vssd vssd vccd vccd _447_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[71\]_TE la_buf\[71\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input500_A la_oenb_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput599 mprj_dat_o_core[25] vssd vssd vccd vccd _457_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[75\] _539_/Y la_buf\[75\]/TE vssd vssd vccd vccd output727/A sky130_fd_sc_hd__einvp_4
XANTENNA_mprj_dat_buf\[23\]_A _455_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[56\]_TE mprj_logic_high_inst/HI[258] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[30\]_A user_wb_dat_gates\[30\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_43_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[95\]_A_N _358_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[33\]_A_N _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output817_A output817/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[48\]_A_N _640_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__478__A _478_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[64\] input92/X user_to_mprj_in_gates\[64\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[64\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA_mprj_dat_buf\[14\]_A _446_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_buffers\[21\]_A user_wb_dat_gates\[21\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_35_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[20\]_TE mprj_dat_buf\[20\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[94\]_TE la_buf\[94\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__388__A _388_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[79\]_TE mprj_logic_high_inst/HI[281] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[9\]_A _601_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_buffers\[12\]_A user_wb_dat_gates\[12\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_40_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input283_A la_iena_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input450_A la_oenb_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input548_A mprj_adr_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput330 la_iena_mprj[48] vssd vssd vccd vccd input330/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput341 la_iena_mprj[58] vssd vssd vccd vccd input341/X sky130_fd_sc_hd__clkbuf_1
Xinput352 la_iena_mprj[68] vssd vssd vccd vccd input352/X sky130_fd_sc_hd__clkbuf_1
Xinput363 la_iena_mprj[78] vssd vssd vccd vccd input363/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput374 la_iena_mprj[88] vssd vssd vccd vccd input374/X sky130_fd_sc_hd__clkbuf_1
Xinput385 la_iena_mprj[98] vssd vssd vccd vccd input385/X sky130_fd_sc_hd__clkbuf_1
Xinput396 la_oenb_mprj[107] vssd vssd vccd vccd _370_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_598_ _598_/A vssd vssd vccd vccd _598_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[34\] user_to_mprj_in_gates\[34\]/Y vssd vssd vccd vccd output810/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output767_A output767/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output934_A output934/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput826 output826/A vssd vssd vccd vccd la_data_in_mprj[49] sky130_fd_sc_hd__buf_2
Xoutput804 output804/A vssd vssd vccd vccd la_data_in_mprj[29] sky130_fd_sc_hd__buf_2
Xoutput815 output815/A vssd vssd vccd vccd la_data_in_mprj[39] sky130_fd_sc_hd__buf_2
Xoutput837 output837/A vssd vssd vccd vccd la_data_in_mprj[59] sky130_fd_sc_hd__buf_2
XFILLER_47_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput848 output848/A vssd vssd vccd vccd la_data_in_mprj[69] sky130_fd_sc_hd__buf_2
Xoutput859 output859/A vssd vssd vccd vccd la_data_in_mprj[79] sky130_fd_sc_hd__buf_2
XFILLER_45_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[25\]_B repeater1125/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output1031_A output1031/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[74\] input359/X mprj_logic_high_inst/HI[404] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[74\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[100\] _363_/Y mprj_logic_high_inst/HI[302] vssd vssd vccd
+ vccd output884/A sky130_fd_sc_hd__einvp_2
XFILLER_24_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[16\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input129_A la_data_out_core[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[30\] _622_/Y mprj_logic_high_inst/HI[232] vssd vssd vccd
+ vccd output934/A sky130_fd_sc_hd__einvp_4
XFILLER_2_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_521_ _521_/A vssd vssd vccd vccd _521_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[52\] _644_/A la_buf_enable\[52\]/B vssd vssd vccd vccd la_buf\[52\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_1465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_452_ _452_/A vssd vssd vccd vccd _452_/Y sky130_fd_sc_hd__inv_4
XFILLER_32_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[1\]_A _465_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_383_ _383_/A vssd vssd vccd vccd _383_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input498_A la_oenb_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input94_A la_data_out_core[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__581__A _581_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[38\] _502_/Y la_buf\[38\]/TE vssd vssd vccd vccd output686/A sky130_fd_sc_hd__einvp_8
XFILLER_13_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[11\]_TE mprj_adr_buf\[11\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_irq_gates\[1\]_A input622/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2150 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput171 la_data_out_mprj[1] vssd vssd vccd vccd _465_/A sky130_fd_sc_hd__clkbuf_2
Xinput160 la_data_out_mprj[125] vssd vssd vccd vccd _589_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput182 la_data_out_mprj[2] vssd vssd vccd vccd _466_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput193 la_data_out_mprj[3] vssd vssd vccd vccd _467_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output884_A output884/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[27\] input51/X user_to_mprj_in_gates\[27\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[27\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_31_152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__491__A _491_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput645 output645/A vssd vssd vccd vccd la_data_in_core[116] sky130_fd_sc_hd__buf_2
Xoutput634 output634/A vssd vssd vccd vccd la_data_in_core[106] sky130_fd_sc_hd__buf_2
Xoutput656 output656/A vssd vssd vccd vccd la_data_in_core[126] sky130_fd_sc_hd__buf_2
Xoutput678 output678/A vssd vssd vccd vccd la_data_in_core[30] sky130_fd_sc_hd__buf_2
Xoutput667 output667/A vssd vssd vccd vccd la_data_in_core[20] sky130_fd_sc_hd__buf_2
XFILLER_47_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput689 output689/A vssd vssd vccd vccd la_data_in_core[40] sky130_fd_sc_hd__buf_2
XTAP_141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_adr_buf\[8\]_A _408_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2076 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1079_A output1079/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[78\] _341_/Y mprj_logic_high_inst/HI[280] vssd vssd vccd
+ vccd output986/A sky130_fd_sc_hd__einvp_4
Xmprj_dat_buf\[26\] _458_/Y mprj_dat_buf\[26\]/TE vssd vssd vccd vccd output1095/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_28_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input246_A la_data_out_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input413_A la_oenb_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__576__A _576_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_504_ _504_/A vssd vssd vccd vccd _504_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_82 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_435_ _435_/A vssd vssd vccd vccd _435_/Y sky130_fd_sc_hd__inv_4
XFILLER_14_675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_366_ _366_/A vssd vssd vccd vccd _366_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[8\]_B mprj_logic_high_inst/HI[338] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[21\] _421_/Y mprj_adr_buf\[21\]/TE vssd vssd vccd vccd output1025/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output632_A output632/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[40\]_A input66/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_64 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__486__A _486_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[6\] _598_/A la_buf_enable\[6\]/B vssd vssd vccd vccd la_buf\[6\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[31\]_A input56/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input1_A caravel_clk vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__396__A _396_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[37\] input318/X mprj_logic_high_inst/HI[367] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[37\]/B sky130_fd_sc_hd__and2_1
XFILLER_15_417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[98\]_A input129/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[15\] _607_/A la_buf_enable\[15\]/B vssd vssd vccd vccd la_buf\[15\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_23_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[28\]_TE la_buf\[28\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input196_A la_data_out_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input363_A la_iena_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input57_A la_data_out_core[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[22\]_A input46/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input530_A mprj_adr_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[120\] _383_/A la_buf_enable\[120\]/B vssd vssd vccd vccd la_buf\[120\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_4_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[89\]_A input119/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_418_ _418_/A vssd vssd vccd vccd _418_/Y sky130_fd_sc_hd__inv_12
XFILLER_14_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_349_ _349_/A vssd vssd vccd vccd _349_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output847_A output847/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput1103 output1103/A vssd vssd vccd vccd mprj_dat_o_user[4] sky130_fd_sc_hd__buf_2
Xoutput1114 output1114/A vssd vssd vccd vccd mprj_we_o_user sky130_fd_sc_hd__buf_2
XFILLER_6_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[94\] input125/X user_to_mprj_in_gates\[94\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[94\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[13\]_A input36/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[8\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1111_A output1111/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[121\]_A_N _384_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[8\]_B user_to_mprj_in_gates\[8\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_47_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input111_A la_data_out_core[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input209_A la_data_out_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input578_A mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input480_A la_oenb_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[20\] _484_/Y la_buf\[20\]/TE vssd vssd vccd vccd output667/A sky130_fd_sc_hd__einvp_8
XFILLER_32_1587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_542 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[64\] user_to_mprj_in_gates\[64\]/Y vssd vssd vccd vccd output843/A
+ sky130_fd_sc_hd__clkinv_4
XTAP_2180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output797_A output797/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_wb_dat_gates\[22\] input564/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[22\]/Y
+ sky130_fd_sc_hd__nand2_2
XANTENNA_output964_A output964/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[120\] input27/X user_to_mprj_in_gates\[120\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[120\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_29_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[110\]_A input272/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output1061_A output1061/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[60\] _652_/Y mprj_logic_high_inst/HI[262] vssd vssd vccd
+ vccd output967/A sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[82\] _345_/A la_buf_enable\[82\]/B vssd vssd vccd vccd la_buf\[82\]/TE
+ sky130_fd_sc_hd__and2b_1
Xinput501 la_oenb_mprj[87] vssd vssd vccd vccd _350_/A sky130_fd_sc_hd__clkbuf_4
Xinput512 la_oenb_mprj[97] vssd vssd vccd vccd _360_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input159_A la_data_out_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput545 mprj_adr_o_core[6] vssd vssd vccd vccd _406_/A sky130_fd_sc_hd__clkbuf_2
Xinput523 mprj_adr_o_core[15] vssd vssd vccd vccd _415_/A sky130_fd_sc_hd__buf_2
XFILLER_5_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput534 mprj_adr_o_core[25] vssd vssd vccd vccd _425_/A sky130_fd_sc_hd__buf_2
Xinput567 mprj_dat_i_user[25] vssd vssd vccd vccd input567/X sky130_fd_sc_hd__clkbuf_2
Xinput578 mprj_dat_i_user[6] vssd vssd vccd vccd input578/X sky130_fd_sc_hd__buf_12
Xinput556 mprj_dat_i_user[15] vssd vssd vccd vccd input556/X sky130_fd_sc_hd__buf_12
XFILLER_44_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input326_A la_iena_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput589 mprj_dat_o_core[16] vssd vssd vccd vccd _448_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[101\]_TE mprj_logic_high_inst/HI[303] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__584__A _584_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[68\] _532_/Y la_buf\[68\]/TE vssd vssd vccd vccd output719/A sky130_fd_sc_hd__einvp_8
XFILLER_16_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[101\]_A input262/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[124\] _588_/Y la_buf\[124\]/TE vssd vssd vccd vccd output654/A sky130_fd_sc_hd__einvp_4
XFILLER_32_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output712_A output712/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[57\] input84/X user_to_mprj_in_gates\[57\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[57\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[119\]_A input25/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__494__A _494_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1560 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[124\]_TE mprj_logic_high_inst/HI[326] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[90\]_A input377/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input276_A la_iena_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_758 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__579__A _579_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input443_A la_oenb_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput320 la_iena_mprj[39] vssd vssd vccd vccd input320/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[23\]_TE mprj_logic_high_inst/HI[225] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xinput331 la_iena_mprj[49] vssd vssd vccd vccd input331/X sky130_fd_sc_hd__clkbuf_1
Xinput342 la_iena_mprj[59] vssd vssd vccd vccd input342/X sky130_fd_sc_hd__clkbuf_1
Xinput353 la_iena_mprj[69] vssd vssd vccd vccd input353/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input610_A mprj_dat_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput364 la_iena_mprj[79] vssd vssd vccd vccd input364/X sky130_fd_sc_hd__clkbuf_1
Xinput375 la_iena_mprj[89] vssd vssd vccd vccd input375/X sky130_fd_sc_hd__clkbuf_1
Xinput386 la_iena_mprj[99] vssd vssd vccd vccd input386/X sky130_fd_sc_hd__clkbuf_1
Xinput397 la_oenb_mprj[108] vssd vssd vccd vccd _371_/A sky130_fd_sc_hd__buf_2
XFILLER_40_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[81\]_A input367/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_597_ _597_/A vssd vssd vccd vccd _597_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[27\] user_to_mprj_in_gates\[27\]/Y vssd vssd vccd vccd output802/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_51_1760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output662_A output662/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput827 output827/A vssd vssd vccd vccd la_data_in_mprj[4] sky130_fd_sc_hd__buf_2
Xoutput816 output816/A vssd vssd vccd vccd la_data_in_mprj[3] sky130_fd_sc_hd__buf_2
Xoutput805 output805/A vssd vssd vccd vccd la_data_in_mprj[2] sky130_fd_sc_hd__buf_2
XANTENNA_output927_A output927/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_97 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput849 output849/A vssd vssd vccd vccd la_data_in_mprj[6] sky130_fd_sc_hd__buf_2
Xoutput838 output838/A vssd vssd vccd vccd la_data_in_mprj[5] sky130_fd_sc_hd__buf_2
XFILLER_45_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__489__A _489_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[72\]_A input357/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[8\]_B la_buf_enable\[8\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[61\]_TE la_buf\[61\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[46\]_TE mprj_logic_high_inst/HI[248] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[94\]_A_N _357_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__399__A _399_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1024_A output1024/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[67\] input351/X mprj_logic_high_inst/HI[397] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[67\]/B sky130_fd_sc_hd__and2_1
XFILLER_2_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_520_ _520_/A vssd vssd vccd vccd _520_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_ena_buf\[63\]_A input347/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[23\] _615_/Y mprj_logic_high_inst/HI[225] vssd vssd vccd
+ vccd output926/A sky130_fd_sc_hd__einvp_4
Xuser_to_mprj_oen_buffers\[5\] _597_/Y mprj_logic_high_inst/HI[207] vssd vssd vccd
+ vccd output966/A sky130_fd_sc_hd__einvp_4
Xla_buf_enable\[45\] _637_/A la_buf_enable\[45\]/B vssd vssd vccd vccd la_buf\[45\]/TE
+ sky130_fd_sc_hd__and2b_1
X_451_ _451_/A vssd vssd vccd vccd _451_/Y sky130_fd_sc_hd__inv_6
X_382_ _382_/A vssd vssd vccd vccd _382_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf_enable\[32\]_A_N _624_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input393_A la_oenb_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input87_A la_data_out_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[47\]_A_N _639_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input560_A mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[10\]_TE mprj_dat_buf\[10\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_irq_gates\[1\]_B user_irq_gates\[1\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput172 la_data_out_mprj[20] vssd vssd vccd vccd _484_/A sky130_fd_sc_hd__clkbuf_2
Xinput150 la_data_out_mprj[116] vssd vssd vccd vccd _580_/A sky130_fd_sc_hd__clkbuf_2
Xinput161 la_data_out_mprj[126] vssd vssd vccd vccd _590_/A sky130_fd_sc_hd__clkbuf_4
Xinput194 la_data_out_mprj[40] vssd vssd vccd vccd _504_/A sky130_fd_sc_hd__clkbuf_2
Xinput183 la_data_out_mprj[30] vssd vssd vccd vccd _494_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[54\]_A input337/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_649_ _649_/A vssd vssd vccd vccd _649_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_17_662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output877_A output877/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[84\]_TE la_buf\[84\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[69\]_TE mprj_logic_high_inst/HI[271] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xoutput635 output635/A vssd vssd vccd vccd la_data_in_core[107] sky130_fd_sc_hd__buf_2
Xoutput657 output657/A vssd vssd vccd vccd la_data_in_core[127] sky130_fd_sc_hd__buf_2
Xoutput646 output646/A vssd vssd vccd vccd la_data_in_core[117] sky130_fd_sc_hd__buf_2
Xoutput679 output679/A vssd vssd vccd vccd la_data_in_core[31] sky130_fd_sc_hd__buf_2
Xoutput668 output668/A vssd vssd vccd vccd la_data_in_core[21] sky130_fd_sc_hd__buf_2
XFILLER_47_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_sel_buf\[2\]_A _398_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[45\]_A input327/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1354 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_514 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_dat_buf\[19\] _451_/Y mprj_dat_buf\[19\]/TE vssd vssd vccd vccd output1087/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input239_A la_data_out_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input141_A la_data_out_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[36\]_A input317/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input406_A la_oenb_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_503_ _503_/A vssd vssd vccd vccd _503_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_434_ _434_/A vssd vssd vccd vccd _434_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_26_492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1296 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__592__A _592_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[50\] _514_/Y la_buf\[50\]/TE vssd vssd vccd vccd output700/A sky130_fd_sc_hd__einvp_8
XTAP_1886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_365_ _365_/A vssd vssd vccd vccd _365_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[122\] input285/X mprj_logic_high_inst/HI[452] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[122\]/B sky130_fd_sc_hd__and2_1
XFILLER_14_687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[3\]_A _435_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2024 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_6 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[14\] _414_/Y mprj_adr_buf\[14\]/TE vssd vssd vccd vccd output1017/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_48_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[40\]_B user_to_mprj_in_gates\[40\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[94\] user_to_mprj_in_gates\[94\]/Y vssd vssd vccd vccd output876/A
+ sky130_fd_sc_hd__inv_2
XFILLER_49_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[27\]_A input307/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output994_A output994/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_buffers\[4\] user_wb_dat_gates\[4\]/Y vssd vssd vccd vccd output1071/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_51_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[31\]_B user_to_mprj_in_gates\[31\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[1\] input43/X user_to_mprj_in_gates\[1\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[1\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_buffers\[92\]_A user_to_mprj_in_gates\[92\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[18\]_A input297/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[98\]_B user_to_mprj_in_gates\[98\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output1091_A output1091/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input189_A la_data_out_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[90\] _353_/Y mprj_logic_high_inst/HI[292] vssd vssd vccd
+ vccd output1000/A sky130_fd_sc_hd__einvp_8
XFILLER_30_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[22\]_B user_to_mprj_in_gates\[22\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_input356_A la_iena_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[83\]_A user_to_mprj_in_gates\[83\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[98\] _562_/Y la_buf\[98\]/TE vssd vssd vccd vccd output752/A sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[3\] input321/X mprj_logic_high_inst/HI[333] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[3\]/B sky130_fd_sc_hd__and2_1
XANTENNA_input523_A mprj_adr_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__587__A _587_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[113\] _376_/A la_buf_enable\[113\]/B vssd vssd vccd vccd la_buf\[113\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_19_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_2304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[89\]_B user_to_mprj_in_gates\[89\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_417_ _417_/A vssd vssd vccd vccd _417_/Y sky130_fd_sc_hd__inv_6
XFILLER_42_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_348_ _348_/A vssd vssd vccd vccd _348_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[121\]_A user_to_mprj_in_gates\[121\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output742_A output742/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput1104 output1104/A vssd vssd vccd vccd mprj_dat_o_user[5] sky130_fd_sc_hd__buf_2
XANTENNA_la_buf\[110\]_A _574_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput1115 output1115/A vssd vssd vccd vccd user1_vcc_powergood sky130_fd_sc_hd__buf_2
XFILLER_45_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[13\]_B user_to_mprj_in_gates\[13\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[74\]_A user_to_mprj_in_gates\[74\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[87\] input117/X user_to_mprj_in_gates\[87\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[87\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__497__A _497_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_532 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[24\]_TE mprj_adr_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[112\]_A user_to_mprj_in_gates\[112\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[101\]_A _565_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[65\]_A user_to_mprj_in_gates\[65\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output1104_A output1104/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input104_A la_data_out_core[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[1\] user_to_mprj_in_gates\[1\]/Y vssd vssd vccd vccd output794/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_38_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input473_A la_oenb_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[103\]_A user_to_mprj_in_gates\[103\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[13\] _477_/Y la_buf\[13\]/TE vssd vssd vccd vccd output659/A sky130_fd_sc_hd__einvp_8
Xla_buf\[9\] _473_/Y la_buf\[9\]/TE vssd vssd vccd vccd output754/A sky130_fd_sc_hd__einvp_8
XFILLER_48_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[56\]_A user_to_mprj_in_gates\[56\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[6\] _406_/Y mprj_adr_buf\[6\]/TE vssd vssd vccd vccd output1040/A sky130_fd_sc_hd__einvp_8
XFILLER_43_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[57\] user_to_mprj_in_gates\[57\]/Y vssd vssd vccd vccd output835/A
+ sky130_fd_sc_hd__clkinv_4
XTAP_2181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output692_A output692/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[96\]_A _560_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output957_A output957/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[15\] input556/X repeater1125/A vssd vssd vccd vccd user_wb_dat_gates\[15\]/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_50_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[47\]_A user_to_mprj_in_gates\[47\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[12\] user_wb_dat_gates\[12\]/Y vssd vssd vccd vccd output1048/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[20\]_A _484_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[113\] input19/X user_to_mprj_in_gates\[113\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[113\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[18\]_TE la_buf\[18\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[87\]_A _551_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[110\]_B mprj_logic_high_inst/HI[440] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1054_A output1054/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[97\] input384/X mprj_logic_high_inst/HI[427] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[97\]/B sky130_fd_sc_hd__and2_1
XFILLER_49_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[38\]_A user_to_mprj_in_gates\[38\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[123\] _386_/Y mprj_logic_high_inst/HI[325] vssd vssd vccd
+ vccd output909/A sky130_fd_sc_hd__einvp_4
XANTENNA_la_buf\[11\]_A _475_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput502 la_oenb_mprj[88] vssd vssd vccd vccd _351_/A sky130_fd_sc_hd__clkbuf_4
Xuser_to_mprj_oen_buffers\[53\] _645_/Y mprj_logic_high_inst/HI[255] vssd vssd vccd
+ vccd output959/A sky130_fd_sc_hd__einvp_8
Xinput513 la_oenb_mprj[98] vssd vssd vccd vccd _361_/A sky130_fd_sc_hd__clkbuf_2
Xinput546 mprj_adr_o_core[7] vssd vssd vccd vccd _407_/A sky130_fd_sc_hd__buf_2
Xinput524 mprj_adr_o_core[16] vssd vssd vccd vccd _416_/A sky130_fd_sc_hd__buf_2
XFILLER_5_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput535 mprj_adr_o_core[26] vssd vssd vccd vccd _426_/A sky130_fd_sc_hd__buf_2
Xinput568 mprj_dat_i_user[26] vssd vssd vccd vccd input568/X sky130_fd_sc_hd__clkbuf_2
Xinput557 mprj_dat_i_user[16] vssd vssd vccd vccd input557/X sky130_fd_sc_hd__buf_12
Xinput579 mprj_dat_i_user[7] vssd vssd vccd vccd input579/X sky130_fd_sc_hd__buf_8
XFILLER_47_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[75\] _338_/A la_buf_enable\[75\]/B vssd vssd vccd vccd la_buf\[75\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_29_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_830 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input319_A la_iena_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input221_A la_data_out_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[78\]_A _542_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[101\]_B mprj_logic_high_inst/HI[431] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_34_72 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input590_A mprj_dat_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[96\]_B la_buf_enable\[96\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[117\] _581_/Y la_buf\[117\]/TE vssd vssd vccd vccd output646/A sky130_fd_sc_hd__einvp_4
XANTENNA_user_to_mprj_in_buffers\[29\]_A user_to_mprj_in_gates\[29\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[110\] user_to_mprj_in_gates\[110\]/Y vssd vssd vccd vccd
+ output767/A sky130_fd_sc_hd__clkinv_4
XTAP_538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[20\]_B la_buf_enable\[20\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output705_A output705/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[119\]_B user_to_mprj_in_gates\[119\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[69\]_A _533_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[87\]_B la_buf_enable\[87\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[120\]_A_N _383_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[28\]_A input570/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[11\]_B la_buf_enable\[11\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[9\]_TE la_buf\[9\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[90\]_B mprj_logic_high_inst/HI[420] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[12\] input291/X mprj_logic_high_inst/HI[342] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[12\]/B sky130_fd_sc_hd__and2_1
XANTENNA_la_buf_enable\[78\]_B la_buf_enable\[78\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[80\]_A _343_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input171_A la_data_out_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input269_A la_iena_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[19\]_A input560/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input436_A la_oenb_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput321 la_iena_mprj[3] vssd vssd vccd vccd input321/X sky130_fd_sc_hd__clkbuf_1
Xinput310 la_iena_mprj[2] vssd vssd vccd vccd input310/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input32_A la_data_out_core[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput354 la_iena_mprj[6] vssd vssd vccd vccd input354/X sky130_fd_sc_hd__clkbuf_1
Xinput343 la_iena_mprj[5] vssd vssd vccd vccd input343/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput332 la_iena_mprj[4] vssd vssd vccd vccd input332/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[80\] _544_/Y la_buf\[80\]/TE vssd vssd vccd vccd output733/A sky130_fd_sc_hd__einvp_4
Xinput387 la_iena_mprj[9] vssd vssd vccd vccd input387/X sky130_fd_sc_hd__clkbuf_2
Xinput365 la_iena_mprj[7] vssd vssd vccd vccd input365/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput376 la_iena_mprj[8] vssd vssd vccd vccd input376/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input603_A mprj_dat_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__595__A _595_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput398 la_oenb_mprj[109] vssd vssd vccd vccd _372_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[81\]_B mprj_logic_high_inst/HI[411] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_32_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_596_ _596_/A vssd vssd vccd vccd _596_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[69\]_B la_buf_enable\[69\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output655_A output655/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[71\]_A _334_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput828 output828/A vssd vssd vccd vccd la_data_in_mprj[50] sky130_fd_sc_hd__buf_2
XFILLER_6_65 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput817 output817/A vssd vssd vccd vccd la_data_in_mprj[40] sky130_fd_sc_hd__buf_2
Xoutput806 output806/A vssd vssd vccd vccd la_data_in_mprj[30] sky130_fd_sc_hd__buf_2
Xoutput839 output839/A vssd vssd vccd vccd la_data_in_mprj[60] sky130_fd_sc_hd__buf_2
XFILLER_45_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output822_A output822/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[72\]_B mprj_logic_high_inst/HI[402] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[62\]_A _654_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[127\]_A _390_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output1017_A output1017/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[63\]_B mprj_logic_high_inst/HI[393] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_450_ _450_/A vssd vssd vccd vccd _450_/Y sky130_fd_sc_hd__inv_6
XFILLER_26_663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[16\] _608_/Y mprj_logic_high_inst/HI[218] vssd vssd vccd
+ vccd output918/A sky130_fd_sc_hd__einvp_4
X_381_ _381_/A vssd vssd vccd vccd _381_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[38\] _630_/A la_buf_enable\[38\]/B vssd vssd vccd vccd la_buf\[38\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_40_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input386_A la_iena_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[53\]_A _645_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[118\]_A _381_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input553_A mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput140 la_data_out_mprj[107] vssd vssd vccd vccd _571_/A sky130_fd_sc_hd__clkbuf_4
Xinput151 la_data_out_mprj[117] vssd vssd vccd vccd _581_/A sky130_fd_sc_hd__clkbuf_4
Xinput162 la_data_out_mprj[127] vssd vssd vccd vccd _591_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput195 la_data_out_mprj[41] vssd vssd vccd vccd _505_/A sky130_fd_sc_hd__clkbuf_2
Xinput173 la_data_out_mprj[21] vssd vssd vccd vccd _485_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput184 la_data_out_mprj[31] vssd vssd vccd vccd _495_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[54\]_B mprj_logic_high_inst/HI[384] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_648_ _648_/A vssd vssd vccd vccd _648_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_17_674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_579_ _579_/A vssd vssd vccd vccd _579_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output772_A output772/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[114\]_TE mprj_logic_high_inst/HI[316] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[44\]_A _636_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[109\]_A _372_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput636 output636/A vssd vssd vccd vccd la_data_in_core[108] sky130_fd_sc_hd__buf_2
XFILLER_47_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput647 output647/A vssd vssd vccd vccd la_data_in_core[118] sky130_fd_sc_hd__buf_2
Xoutput669 output669/A vssd vssd vccd vccd la_data_in_core[22] sky130_fd_sc_hd__buf_2
Xoutput658 output658/A vssd vssd vccd vccd la_data_in_core[12] sky130_fd_sc_hd__buf_2
XFILLER_47_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[45\]_B mprj_logic_high_inst/HI[375] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_42_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2056 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[13\]_TE mprj_logic_high_inst/HI[215] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[35\]_A _627_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_6 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[31\]_A _431_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input134_A la_data_out_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[36\]_B mprj_logic_high_inst/HI[366] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_502_ _502_/A vssd vssd vccd vccd _502_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input301_A la_iena_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_433_ _433_/A vssd vssd vccd vccd _433_/Y sky130_fd_sc_hd__inv_4
XTAP_1876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[43\] _507_/Y la_buf\[43\]/TE vssd vssd vccd vccd output692/A sky130_fd_sc_hd__einvp_8
X_364_ _364_/A vssd vssd vccd vccd _364_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[115\] input277/X mprj_logic_high_inst/HI[445] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[115\]/B sky130_fd_sc_hd__and2_1
XFILLER_42_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[26\]_A _618_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_850 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_11 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[87\] user_to_mprj_in_gates\[87\]/Y vssd vssd vccd vccd output868/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_3_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[22\]_A _422_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[51\]_TE la_buf\[51\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[27\]_B mprj_logic_high_inst/HI[357] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_output987_A output987/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[32\] input57/X user_to_mprj_in_gates\[32\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[32\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[36\]_TE mprj_logic_high_inst/HI[238] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[93\]_A_N _356_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[17\]_A _609_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[31\]_A_N _623_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[13\]_A _413_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[46\]_A_N _638_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[18\]_B mprj_logic_high_inst/HI[348] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output1084_A output1084/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[83\] _346_/Y mprj_logic_high_inst/HI[285] vssd vssd vccd
+ vccd output992/A sky130_fd_sc_hd__einvp_4
XFILLER_30_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[31\] _463_/Y mprj_dat_buf\[31\]/TE vssd vssd vccd vccd output1101/A
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input349_A la_iena_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input251_A la_data_out_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input516_A mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[74\]_TE la_buf\[74\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[106\] _369_/A la_buf_enable\[106\]/B vssd vssd vccd vccd la_buf\[106\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_19_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[59\]_TE mprj_logic_high_inst/HI[261] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_416_ _416_/A vssd vssd vccd vccd _416_/Y sky130_fd_sc_hd__inv_12
XFILLER_53_82 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_347_ _347_/A vssd vssd vccd vccd _347_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput1105 output1105/A vssd vssd vccd vccd mprj_dat_o_user[6] sky130_fd_sc_hd__buf_2
XFILLER_48_1722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput1116 output1116/A vssd vssd vccd vccd user1_vdd_powergood sky130_fd_sc_hd__buf_2
XANTENNA_output735_A output735/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output902_A output902/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[23\]_TE mprj_dat_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[2\]_TE mprj_logic_high_inst/HI[204] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[97\]_TE la_buf\[97\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[42\] input324/X mprj_logic_high_inst/HI[372] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[42\]/B sky130_fd_sc_hd__and2_1
XFILLER_5_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[20\] _612_/A la_buf_enable\[20\]/B vssd vssd vccd vccd la_buf\[20\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_32_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input299_A la_iena_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input62_A la_data_out_core[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input466_A la_oenb_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__598__A _598_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[26\]_A _458_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output685_A output685/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1710 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_786 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output852_A output852/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[17\]_A _449_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1758 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_buffers\[24\]_A user_wb_dat_gates\[24\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[106\] input11/X user_to_mprj_in_gates\[106\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[106\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output1047_A output1047/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[116\] _379_/Y mprj_logic_high_inst/HI[318] vssd vssd vccd
+ vccd output901/A sky130_fd_sc_hd__einvp_4
Xinput503 la_oenb_mprj[89] vssd vssd vccd vccd _352_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput514 la_oenb_mprj[99] vssd vssd vccd vccd _362_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput525 mprj_adr_o_core[17] vssd vssd vccd vccd _417_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput536 mprj_adr_o_core[27] vssd vssd vccd vccd _427_/A sky130_fd_sc_hd__buf_2
Xinput569 mprj_dat_i_user[27] vssd vssd vccd vccd input569/X sky130_fd_sc_hd__clkbuf_2
Xinput558 mprj_dat_i_user[17] vssd vssd vccd vccd input558/X sky130_fd_sc_hd__buf_12
XFILLER_47_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput547 mprj_adr_o_core[8] vssd vssd vccd vccd _408_/A sky130_fd_sc_hd__buf_2
XFILLER_5_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[46\] _638_/Y mprj_logic_high_inst/HI[248] vssd vssd vccd
+ vccd output951/A sky130_fd_sc_hd__einvp_2
Xla_buf_enable\[68\] _331_/A la_buf_enable\[68\]/B vssd vssd vccd vccd la_buf\[68\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_28_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_buffers\[15\]_A user_wb_dat_gates\[15\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_40_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input214_A la_data_out_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input583_A mprj_dat_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1998 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[14\]_TE mprj_adr_buf\[14\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[103\] user_to_mprj_in_gates\[103\]/Y vssd vssd vccd vccd
+ output759/A sky130_fd_sc_hd__clkinv_4
XFILLER_43_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1830 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[28\]_B repeater1125/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[2\] _434_/Y mprj_dat_buf\[2\]/TE vssd vssd vccd vccd output1099/A sky130_fd_sc_hd__einvp_8
XFILLER_44_1268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_dat_buf\[2\]_TE mprj_dat_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[110\]_B la_buf_enable\[110\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[122\]_TE la_buf\[122\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_buffers\[1\]_A user_wb_dat_gates\[1\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input164_A la_data_out_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[19\]_B repeater1125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput300 la_iena_mprj[20] vssd vssd vccd vccd input300/X sky130_fd_sc_hd__clkbuf_1
Xinput311 la_iena_mprj[30] vssd vssd vccd vccd input311/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_988 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input331_A la_iena_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput333 la_iena_mprj[50] vssd vssd vccd vccd input333/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input429_A la_oenb_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput322 la_iena_mprj[40] vssd vssd vccd vccd input322/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput344 la_iena_mprj[60] vssd vssd vccd vccd input344/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input25_A la_data_out_core[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_95 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput388 la_oenb_mprj[0] vssd vssd vccd vccd _592_/A sky130_fd_sc_hd__clkbuf_2
Xinput355 la_iena_mprj[70] vssd vssd vccd vccd input355/X sky130_fd_sc_hd__clkbuf_1
Xinput366 la_iena_mprj[80] vssd vssd vccd vccd input366/X sky130_fd_sc_hd__clkbuf_1
Xinput377 la_iena_mprj[90] vssd vssd vccd vccd input377/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput399 la_oenb_mprj[10] vssd vssd vccd vccd _602_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[73\] _537_/Y la_buf\[73\]/TE vssd vssd vccd vccd output725/A sky130_fd_sc_hd__einvp_4
XANTENNA_la_buf\[4\]_A _468_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[101\]_B la_buf_enable\[101\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_595_ _595_/A vssd vssd vccd vccd _595_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1702 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput818 output818/A vssd vssd vccd vccd la_data_in_mprj[41] sky130_fd_sc_hd__buf_2
Xoutput807 output807/A vssd vssd vccd vccd la_data_in_mprj[31] sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_gates\[70\]_A input99/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output648_A output648/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput829 output829/A vssd vssd vccd vccd la_data_in_mprj[51] sky130_fd_sc_hd__buf_2
XFILLER_45_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output815_A output815/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[62\] input90/X user_to_mprj_in_gates\[62\]/B vssd vssd vccd
+ vccd user_to_mprj_in_gates\[62\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[61\]_A input89/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_380_ _380_/A vssd vssd vccd vccd _380_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[92\]_TE mprj_logic_high_inst/HI[294] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input281_A la_iena_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_63 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input379_A la_iena_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[52\]_A input79/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input546_A mprj_adr_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput130 la_data_out_core[99] vssd vssd vccd vccd input130/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput163 la_data_out_mprj[12] vssd vssd vccd vccd _476_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput141 la_data_out_mprj[108] vssd vssd vccd vccd _572_/A sky130_fd_sc_hd__clkbuf_2
Xinput152 la_data_out_mprj[118] vssd vssd vccd vccd _582_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput196 la_data_out_mprj[42] vssd vssd vccd vccd _506_/A sky130_fd_sc_hd__clkbuf_2
Xinput174 la_data_out_mprj[22] vssd vssd vccd vccd _486_/A sky130_fd_sc_hd__clkbuf_2
Xinput185 la_data_out_mprj[32] vssd vssd vccd vccd _496_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_647_ _647_/A vssd vssd vccd vccd _647_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_38_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_578_ _578_/A vssd vssd vccd vccd _578_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[2\]_A user_to_mprj_in_gates\[2\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[32\] user_to_mprj_in_gates\[32\]/Y vssd vssd vccd vccd output808/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output765_A output765/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output932_A output932/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[43\]_A input69/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput648 output648/A vssd vssd vccd vccd la_data_in_core[119] sky130_fd_sc_hd__buf_2
Xoutput637 output637/A vssd vssd vccd vccd la_data_in_core[109] sky130_fd_sc_hd__buf_2
Xoutput659 output659/A vssd vssd vccd vccd la_data_in_core[13] sky130_fd_sc_hd__buf_2
XFILLER_47_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

