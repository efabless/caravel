magic
tech sky130A
magscale 1 2
timestamp 1638030917
<< locali >>
rect 5089 13311 5123 13481
rect 6193 11543 6227 11713
rect 10333 10455 10367 10557
rect 10149 9911 10183 10081
rect 6193 9367 6227 9469
rect 7481 7939 7515 8041
rect 10425 7191 10459 7293
rect 10701 6647 10735 6817
rect 10609 5083 10643 5185
rect 5549 3043 5583 3145
<< viali >>
rect 5089 13481 5123 13515
rect 10241 13481 10275 13515
rect 2421 13345 2455 13379
rect 3525 13345 3559 13379
rect 4905 13345 4939 13379
rect 7665 13413 7699 13447
rect 11529 13413 11563 13447
rect 5917 13345 5951 13379
rect 7021 13345 7055 13379
rect 7205 13345 7239 13379
rect 8953 13345 8987 13379
rect 10793 13345 10827 13379
rect 11989 13345 12023 13379
rect 12173 13345 12207 13379
rect 1869 13277 1903 13311
rect 2513 13277 2547 13311
rect 3341 13277 3375 13311
rect 4353 13277 4387 13311
rect 5089 13277 5123 13311
rect 5181 13277 5215 13311
rect 5641 13277 5675 13311
rect 5825 13277 5859 13311
rect 9597 13277 9631 13311
rect 12357 13277 12391 13311
rect 2329 13209 2363 13243
rect 2973 13209 3007 13243
rect 3065 13209 3099 13243
rect 3433 13209 3467 13243
rect 4813 13209 4847 13243
rect 5733 13209 5767 13243
rect 9413 13209 9447 13243
rect 9505 13209 9539 13243
rect 10057 13209 10091 13243
rect 10149 13209 10183 13243
rect 10701 13209 10735 13243
rect 12817 13209 12851 13243
rect 12909 13209 12943 13243
rect 3157 13141 3191 13175
rect 7297 13141 7331 13175
rect 10609 13141 10643 13175
rect 11897 13141 11931 13175
rect 6377 12937 6411 12971
rect 7389 12937 7423 12971
rect 2973 12869 3007 12903
rect 3249 12869 3283 12903
rect 5825 12869 5859 12903
rect 6929 12869 6963 12903
rect 7941 12869 7975 12903
rect 10333 12869 10367 12903
rect 1409 12801 1443 12835
rect 2881 12801 2915 12835
rect 3525 12801 3559 12835
rect 4445 12801 4479 12835
rect 5181 12801 5215 12835
rect 6101 12801 6135 12835
rect 6561 12801 6595 12835
rect 7021 12801 7055 12835
rect 7757 12801 7791 12835
rect 8033 12801 8067 12835
rect 8953 12801 8987 12835
rect 9689 12801 9723 12835
rect 10609 12801 10643 12835
rect 11621 12801 11655 12835
rect 11897 12801 11931 12835
rect 12817 12801 12851 12835
rect 3433 12733 3467 12767
rect 6837 12733 6871 12767
rect 9597 12733 9631 12767
rect 10793 12733 10827 12767
rect 11345 12733 11379 12767
rect 11805 12733 11839 12767
rect 4813 12665 4847 12699
rect 11253 12665 11287 12699
rect 13185 12665 13219 12699
rect 3341 12393 3375 12427
rect 3801 12393 3835 12427
rect 9873 12393 9907 12427
rect 10149 12393 10183 12427
rect 12541 12393 12575 12427
rect 12909 12393 12943 12427
rect 6193 12325 6227 12359
rect 7757 12325 7791 12359
rect 8401 12325 8435 12359
rect 4261 12257 4295 12291
rect 4353 12257 4387 12291
rect 5549 12257 5583 12291
rect 5733 12257 5767 12291
rect 7941 12257 7975 12291
rect 9229 12257 9263 12291
rect 9413 12257 9447 12291
rect 10885 12257 10919 12291
rect 10977 12257 11011 12291
rect 2145 12189 2179 12223
rect 2881 12189 2915 12223
rect 3065 12189 3099 12223
rect 4997 12189 5031 12223
rect 6285 12189 6319 12223
rect 7481 12189 7515 12223
rect 9965 12189 9999 12223
rect 11529 12189 11563 12223
rect 12173 12189 12207 12223
rect 12449 12189 12483 12223
rect 12725 12189 12759 12223
rect 13185 12189 13219 12223
rect 3249 12121 3283 12155
rect 4169 12121 4203 12155
rect 8493 12121 8527 12155
rect 8677 12121 8711 12155
rect 12817 12121 12851 12155
rect 5089 12053 5123 12087
rect 5825 12053 5859 12087
rect 8585 12053 8619 12087
rect 9505 12053 9539 12087
rect 10425 12053 10459 12087
rect 10793 12053 10827 12087
rect 13277 12053 13311 12087
rect 1409 11849 1443 11883
rect 1777 11849 1811 11883
rect 4077 11849 4111 11883
rect 5917 11849 5951 11883
rect 9229 11849 9263 11883
rect 9689 11849 9723 11883
rect 10241 11849 10275 11883
rect 2697 11781 2731 11815
rect 7757 11781 7791 11815
rect 8585 11781 8619 11815
rect 12449 11781 12483 11815
rect 13461 11781 13495 11815
rect 2881 11713 2915 11747
rect 4169 11713 4203 11747
rect 6101 11713 6135 11747
rect 6193 11713 6227 11747
rect 6377 11713 6411 11747
rect 6653 11713 6687 11747
rect 7113 11713 7147 11747
rect 7297 11713 7331 11747
rect 7481 11713 7515 11747
rect 8401 11713 8435 11747
rect 9045 11713 9079 11747
rect 9597 11713 9631 11747
rect 10701 11713 10735 11747
rect 10793 11713 10827 11747
rect 11529 11713 11563 11747
rect 11713 11713 11747 11747
rect 12541 11713 12575 11747
rect 13277 11713 13311 11747
rect 1869 11645 1903 11679
rect 1961 11645 1995 11679
rect 2237 11645 2271 11679
rect 2789 11645 2823 11679
rect 3433 11645 3467 11679
rect 3893 11645 3927 11679
rect 4629 11645 4663 11679
rect 5181 11645 5215 11679
rect 5273 11645 5307 11679
rect 5825 11645 5859 11679
rect 3341 11577 3375 11611
rect 5089 11577 5123 11611
rect 5365 11577 5399 11611
rect 8493 11645 8527 11679
rect 9781 11645 9815 11679
rect 10517 11645 10551 11679
rect 6469 11577 6503 11611
rect 10149 11577 10183 11611
rect 11621 11577 11655 11611
rect 4537 11509 4571 11543
rect 6193 11509 6227 11543
rect 6837 11509 6871 11543
rect 11161 11509 11195 11543
rect 12357 11509 12391 11543
rect 3341 11305 3375 11339
rect 5825 11305 5859 11339
rect 8309 11305 8343 11339
rect 8953 11305 8987 11339
rect 10149 11305 10183 11339
rect 11253 11305 11287 11339
rect 3065 11237 3099 11271
rect 5273 11237 5307 11271
rect 6193 11237 6227 11271
rect 7205 11237 7239 11271
rect 12817 11237 12851 11271
rect 6561 11169 6595 11203
rect 9413 11169 9447 11203
rect 9505 11169 9539 11203
rect 10425 11169 10459 11203
rect 10885 11169 10919 11203
rect 1593 11101 1627 11135
rect 3065 11101 3099 11135
rect 3249 11101 3283 11135
rect 3985 11101 4019 11135
rect 4905 11101 4939 11135
rect 6009 11101 6043 11135
rect 6101 11101 6135 11135
rect 6285 11101 6319 11135
rect 8125 11101 8159 11135
rect 8401 11101 8435 11135
rect 8585 11101 8619 11135
rect 10333 11101 10367 11135
rect 10517 11101 10551 11135
rect 10609 11101 10643 11135
rect 10793 11101 10827 11135
rect 11069 11101 11103 11135
rect 11529 11101 11563 11135
rect 13001 11101 13035 11135
rect 13185 11101 13219 11135
rect 6745 11033 6779 11067
rect 6837 11033 6871 11067
rect 8769 11033 8803 11067
rect 9321 11033 9355 11067
rect 13369 10965 13403 10999
rect 2145 10761 2179 10795
rect 3617 10761 3651 10795
rect 4353 10761 4387 10795
rect 11069 10761 11103 10795
rect 11529 10761 11563 10795
rect 11989 10761 12023 10795
rect 3341 10693 3375 10727
rect 4445 10693 4479 10727
rect 4813 10693 4847 10727
rect 6377 10693 6411 10727
rect 6561 10693 6595 10727
rect 6745 10693 6779 10727
rect 7941 10693 7975 10727
rect 8769 10693 8803 10727
rect 11897 10693 11931 10727
rect 12909 10693 12943 10727
rect 13553 10693 13587 10727
rect 1685 10625 1719 10659
rect 1777 10625 1811 10659
rect 2605 10625 2639 10659
rect 3525 10625 3559 10659
rect 3801 10625 3835 10659
rect 4537 10625 4571 10659
rect 5457 10625 5491 10659
rect 5825 10625 5859 10659
rect 5917 10625 5951 10659
rect 6101 10625 6135 10659
rect 7113 10625 7147 10659
rect 7205 10625 7239 10659
rect 7389 10625 7423 10659
rect 7849 10625 7883 10659
rect 8401 10625 8435 10659
rect 8585 10625 8619 10659
rect 9781 10625 9815 10659
rect 10149 10625 10183 10659
rect 10425 10625 10459 10659
rect 10609 10625 10643 10659
rect 10701 10625 10735 10659
rect 10885 10625 10919 10659
rect 12357 10625 12391 10659
rect 12817 10625 12851 10659
rect 13001 10625 13035 10659
rect 13461 10625 13495 10659
rect 1501 10557 1535 10591
rect 7665 10557 7699 10591
rect 9873 10557 9907 10591
rect 10333 10557 10367 10591
rect 10793 10557 10827 10591
rect 12173 10557 12207 10591
rect 6009 10489 6043 10523
rect 6929 10489 6963 10523
rect 7297 10489 7331 10523
rect 8309 10489 8343 10523
rect 5641 10421 5675 10455
rect 9505 10421 9539 10455
rect 9965 10421 9999 10455
rect 10057 10421 10091 10455
rect 10333 10421 10367 10455
rect 3065 10217 3099 10251
rect 5733 10217 5767 10251
rect 6929 10217 6963 10251
rect 7297 10217 7331 10251
rect 10333 10217 10367 10251
rect 10885 10217 10919 10251
rect 11161 10217 11195 10251
rect 11529 10217 11563 10251
rect 12725 10217 12759 10251
rect 9321 10149 9355 10183
rect 10701 10149 10735 10183
rect 5273 10081 5307 10115
rect 5457 10081 5491 10115
rect 6101 10081 6135 10115
rect 7481 10081 7515 10115
rect 8585 10081 8619 10115
rect 9413 10081 9447 10115
rect 10149 10081 10183 10115
rect 13277 10081 13311 10115
rect 3801 10013 3835 10047
rect 5181 10013 5215 10047
rect 6009 10013 6043 10047
rect 6193 10013 6227 10047
rect 6285 10013 6319 10047
rect 6469 10013 6503 10047
rect 7205 10013 7239 10047
rect 7389 10013 7423 10047
rect 7573 10013 7607 10047
rect 8401 10013 8435 10047
rect 8953 10013 8987 10047
rect 9229 10013 9263 10047
rect 9505 10013 9539 10047
rect 9689 10013 9723 10047
rect 2973 9945 3007 9979
rect 8493 9945 8527 9979
rect 10609 10013 10643 10047
rect 10793 10013 10827 10047
rect 10977 10013 11011 10047
rect 11161 10013 11195 10047
rect 11345 10013 11379 10047
rect 12449 10013 12483 10047
rect 13093 9945 13127 9979
rect 3893 9877 3927 9911
rect 4813 9877 4847 9911
rect 8033 9877 8067 9911
rect 10149 9877 10183 9911
rect 12541 9877 12575 9911
rect 13185 9877 13219 9911
rect 8769 9673 8803 9707
rect 3433 9605 3467 9639
rect 5089 9605 5123 9639
rect 7849 9605 7883 9639
rect 8033 9605 8067 9639
rect 8309 9605 8343 9639
rect 9045 9605 9079 9639
rect 10609 9605 10643 9639
rect 10793 9605 10827 9639
rect 10977 9605 11011 9639
rect 1685 9537 1719 9571
rect 3157 9537 3191 9571
rect 3709 9537 3743 9571
rect 4353 9537 4387 9571
rect 4629 9537 4663 9571
rect 5181 9537 5215 9571
rect 6469 9537 6503 9571
rect 6745 9537 6779 9571
rect 6837 9537 6871 9571
rect 7205 9537 7239 9571
rect 8493 9537 8527 9571
rect 8601 9537 8635 9571
rect 9229 9537 9263 9571
rect 9321 9537 9355 9571
rect 9505 9537 9539 9571
rect 10425 9537 10459 9571
rect 10885 9537 10919 9571
rect 11529 9537 11563 9571
rect 12541 9537 12575 9571
rect 13369 9537 13403 9571
rect 4997 9469 5031 9503
rect 6193 9469 6227 9503
rect 2973 9401 3007 9435
rect 9413 9401 9447 9435
rect 12817 9401 12851 9435
rect 4445 9333 4479 9367
rect 5549 9333 5583 9367
rect 6193 9333 6227 9367
rect 6929 9333 6963 9367
rect 7021 9333 7055 9367
rect 7757 9333 7791 9367
rect 8309 9333 8343 9367
rect 13277 9333 13311 9367
rect 2237 9129 2271 9163
rect 6285 9129 6319 9163
rect 8033 9129 8067 9163
rect 9137 9129 9171 9163
rect 9505 9129 9539 9163
rect 10701 9129 10735 9163
rect 11253 9129 11287 9163
rect 2881 9061 2915 9095
rect 3341 9061 3375 9095
rect 3893 9061 3927 9095
rect 6653 9061 6687 9095
rect 7297 9061 7331 9095
rect 12449 9061 12483 9095
rect 1593 8993 1627 9027
rect 1777 8993 1811 9027
rect 2421 8993 2455 9027
rect 3801 8993 3835 9027
rect 4353 8993 4387 9027
rect 9229 8993 9263 9027
rect 12541 8993 12575 9027
rect 1869 8925 1903 8959
rect 2973 8925 3007 8959
rect 3617 8925 3651 8959
rect 4445 8925 4479 8959
rect 6469 8925 6503 8959
rect 6561 8925 6595 8959
rect 6745 8925 6779 8959
rect 7481 8925 7515 8959
rect 9137 8925 9171 8959
rect 10149 8925 10183 8959
rect 11161 8925 11195 8959
rect 11713 8925 11747 8959
rect 11989 8925 12023 8959
rect 12633 8925 12667 8959
rect 13369 8925 13403 8959
rect 3157 8857 3191 8891
rect 4629 8857 4663 8891
rect 7849 8857 7883 8891
rect 8125 8857 8159 8891
rect 8309 8857 8343 8891
rect 9689 8857 9723 8891
rect 9873 8857 9907 8891
rect 10057 8857 10091 8891
rect 10701 8857 10735 8891
rect 10885 8857 10919 8891
rect 10977 8857 11011 8891
rect 13553 8857 13587 8891
rect 3433 8789 3467 8823
rect 4813 8789 4847 8823
rect 7573 8789 7607 8823
rect 7665 8789 7699 8823
rect 10241 8789 10275 8823
rect 10517 8789 10551 8823
rect 11805 8789 11839 8823
rect 6837 8585 6871 8619
rect 7297 8585 7331 8619
rect 7941 8585 7975 8619
rect 8033 8585 8067 8619
rect 8861 8585 8895 8619
rect 3157 8517 3191 8551
rect 3249 8517 3283 8551
rect 8217 8517 8251 8551
rect 8493 8517 8527 8551
rect 8677 8517 8711 8551
rect 10425 8517 10459 8551
rect 1593 8449 1627 8483
rect 3065 8449 3099 8483
rect 3433 8449 3467 8483
rect 4169 8449 4203 8483
rect 4445 8449 4479 8483
rect 5917 8449 5951 8483
rect 6561 8449 6595 8483
rect 7205 8449 7239 8483
rect 7665 8449 7699 8483
rect 7849 8449 7883 8483
rect 8309 8449 8343 8483
rect 8769 8449 8803 8483
rect 9505 8449 9539 8483
rect 9689 8449 9723 8483
rect 9781 8449 9815 8483
rect 9965 8449 9999 8483
rect 10241 8449 10275 8483
rect 10701 8449 10735 8483
rect 11345 8449 11379 8483
rect 11529 8449 11563 8483
rect 12449 8449 12483 8483
rect 13185 8449 13219 8483
rect 7481 8381 7515 8415
rect 9597 8381 9631 8415
rect 10609 8381 10643 8415
rect 10793 8381 10827 8415
rect 5733 8313 5767 8347
rect 10885 8313 10919 8347
rect 12817 8313 12851 8347
rect 6469 8245 6503 8279
rect 9321 8245 9355 8279
rect 10149 8245 10183 8279
rect 13369 8245 13403 8279
rect 2145 8041 2179 8075
rect 4353 8041 4387 8075
rect 7481 8041 7515 8075
rect 10977 8041 11011 8075
rect 3065 7973 3099 8007
rect 4169 7973 4203 8007
rect 5365 7973 5399 8007
rect 8953 7973 8987 8007
rect 13277 7973 13311 8007
rect 1501 7905 1535 7939
rect 1685 7905 1719 7939
rect 2237 7905 2271 7939
rect 2973 7905 3007 7939
rect 3525 7905 3559 7939
rect 4905 7905 4939 7939
rect 5457 7905 5491 7939
rect 6837 7905 6871 7939
rect 7297 7905 7331 7939
rect 7481 7905 7515 7939
rect 7573 7905 7607 7939
rect 8677 7905 8711 7939
rect 9505 7905 9539 7939
rect 11253 7905 11287 7939
rect 12817 7905 12851 7939
rect 13369 7905 13403 7939
rect 2697 7837 2731 7871
rect 3801 7837 3835 7871
rect 4445 7837 4479 7871
rect 4629 7837 4663 7871
rect 5733 7837 5767 7871
rect 6009 7837 6043 7871
rect 6653 7837 6687 7871
rect 7757 7837 7791 7871
rect 8217 7837 8251 7871
rect 8769 7837 8803 7871
rect 9321 7837 9355 7871
rect 9873 7837 9907 7871
rect 10057 7837 10091 7871
rect 10517 7837 10551 7871
rect 11069 7837 11103 7871
rect 11713 7837 11747 7871
rect 11989 7837 12023 7871
rect 12725 7837 12759 7871
rect 1777 7769 1811 7803
rect 2789 7769 2823 7803
rect 6745 7769 6779 7803
rect 8033 7769 8067 7803
rect 8125 7769 8159 7803
rect 9413 7769 9447 7803
rect 11161 7769 11195 7803
rect 11805 7769 11839 7803
rect 4169 7701 4203 7735
rect 8309 7701 8343 7735
rect 9873 7701 9907 7735
rect 10609 7701 10643 7735
rect 3065 7497 3099 7531
rect 3157 7497 3191 7531
rect 6653 7497 6687 7531
rect 7941 7497 7975 7531
rect 8033 7497 8067 7531
rect 10885 7497 10919 7531
rect 11989 7497 12023 7531
rect 12265 7497 12299 7531
rect 8677 7429 8711 7463
rect 9505 7429 9539 7463
rect 12633 7429 12667 7463
rect 2421 7361 2455 7395
rect 2605 7361 2639 7395
rect 2881 7361 2915 7395
rect 3617 7361 3651 7395
rect 3893 7361 3927 7395
rect 4445 7361 4479 7395
rect 6469 7361 6503 7395
rect 6929 7361 6963 7395
rect 7297 7361 7331 7395
rect 7573 7361 7607 7395
rect 8401 7361 8435 7395
rect 8585 7361 8619 7395
rect 8821 7361 8855 7395
rect 9137 7361 9171 7395
rect 9321 7361 9355 7395
rect 9689 7361 9723 7395
rect 9873 7361 9907 7395
rect 10149 7361 10183 7395
rect 10333 7361 10367 7395
rect 11529 7361 11563 7395
rect 12173 7361 12207 7395
rect 12725 7361 12759 7395
rect 13369 7361 13403 7395
rect 7113 7293 7147 7327
rect 7832 7293 7866 7327
rect 8125 7293 8159 7327
rect 9965 7293 9999 7327
rect 10057 7293 10091 7327
rect 10425 7293 10459 7327
rect 10977 7293 11011 7327
rect 11069 7293 11103 7327
rect 12817 7293 12851 7327
rect 2421 7225 2455 7259
rect 3893 7225 3927 7259
rect 7021 7225 7055 7259
rect 4445 7157 4479 7191
rect 7389 7157 7423 7191
rect 8953 7157 8987 7191
rect 10425 7157 10459 7191
rect 10517 7157 10551 7191
rect 11621 7157 11655 7191
rect 13185 7157 13219 7191
rect 3893 6953 3927 6987
rect 5076 6953 5110 6987
rect 6561 6953 6595 6987
rect 7389 6953 7423 6987
rect 12817 6953 12851 6987
rect 10057 6885 10091 6919
rect 11805 6885 11839 6919
rect 6837 6817 6871 6851
rect 8677 6817 8711 6851
rect 8769 6817 8803 6851
rect 9413 6817 9447 6851
rect 9505 6817 9539 6851
rect 10701 6817 10735 6851
rect 11437 6817 11471 6851
rect 13369 6817 13403 6851
rect 2605 6749 2639 6783
rect 3341 6749 3375 6783
rect 3801 6749 3835 6783
rect 3985 6749 4019 6783
rect 4813 6749 4847 6783
rect 6929 6749 6963 6783
rect 7205 6749 7239 6783
rect 7568 6749 7602 6783
rect 7885 6749 7919 6783
rect 8033 6749 8067 6783
rect 8401 6749 8435 6783
rect 8493 6749 8527 6783
rect 9229 6749 9263 6783
rect 9321 6749 9355 6783
rect 9689 6749 9723 6783
rect 10189 6749 10223 6783
rect 10333 6749 10367 6783
rect 10609 6749 10643 6783
rect 7113 6681 7147 6715
rect 7665 6681 7699 6715
rect 7757 6681 7791 6715
rect 8217 6681 8251 6715
rect 10425 6681 10459 6715
rect 10793 6749 10827 6783
rect 10977 6749 11011 6783
rect 11069 6749 11103 6783
rect 11195 6749 11229 6783
rect 11713 6749 11747 6783
rect 12235 6749 12269 6783
rect 12541 6749 12575 6783
rect 13185 6749 13219 6783
rect 2789 6613 2823 6647
rect 3249 6613 3283 6647
rect 9045 6613 9079 6647
rect 10701 6613 10735 6647
rect 12173 6613 12207 6647
rect 12357 6613 12391 6647
rect 12725 6613 12759 6647
rect 13277 6613 13311 6647
rect 5825 6409 5859 6443
rect 6193 6409 6227 6443
rect 8125 6409 8159 6443
rect 10425 6409 10459 6443
rect 13461 6409 13495 6443
rect 10517 6341 10551 6375
rect 11069 6341 11103 6375
rect 11989 6341 12023 6375
rect 3893 6273 3927 6307
rect 4629 6273 4663 6307
rect 5365 6273 5399 6307
rect 5641 6273 5675 6307
rect 6009 6273 6043 6307
rect 8401 6273 8435 6307
rect 8861 6273 8895 6307
rect 9045 6273 9079 6307
rect 9597 6273 9631 6307
rect 9781 6273 9815 6307
rect 10057 6273 10091 6307
rect 10313 6273 10347 6307
rect 10701 6273 10735 6307
rect 10885 6273 10919 6307
rect 11345 6273 11379 6307
rect 1685 6205 1719 6239
rect 1961 6205 1995 6239
rect 6377 6205 6411 6239
rect 6653 6205 6687 6239
rect 10609 6205 10643 6239
rect 11713 6205 11747 6239
rect 3801 6137 3835 6171
rect 8953 6137 8987 6171
rect 3433 6069 3467 6103
rect 4077 6069 4111 6103
rect 5181 6069 5215 6103
rect 8493 6069 8527 6103
rect 9689 6069 9723 6103
rect 10057 6069 10091 6103
rect 11161 6069 11195 6103
rect 7665 5865 7699 5899
rect 8677 5865 8711 5899
rect 11529 5865 11563 5899
rect 13461 5865 13495 5899
rect 2789 5797 2823 5831
rect 7941 5797 7975 5831
rect 2237 5729 2271 5763
rect 3157 5729 3191 5763
rect 8125 5729 8159 5763
rect 8217 5729 8251 5763
rect 10057 5729 10091 5763
rect 1685 5661 1719 5695
rect 1961 5661 1995 5695
rect 2053 5661 2087 5695
rect 2513 5661 2547 5695
rect 2881 5661 2915 5695
rect 3065 5661 3099 5695
rect 3893 5661 3927 5695
rect 7573 5661 7607 5695
rect 8033 5661 8067 5695
rect 8401 5661 8435 5695
rect 8493 5661 8527 5695
rect 8953 5661 8987 5695
rect 9046 5661 9080 5695
rect 9229 5661 9263 5695
rect 9321 5661 9355 5695
rect 9418 5661 9452 5695
rect 9781 5661 9815 5695
rect 11713 5661 11747 5695
rect 1593 5593 1627 5627
rect 3341 5593 3375 5627
rect 3525 5593 3559 5627
rect 4169 5593 4203 5627
rect 11989 5593 12023 5627
rect 5641 5525 5675 5559
rect 9597 5525 9631 5559
rect 1961 5321 1995 5355
rect 4169 5321 4203 5355
rect 6469 5321 6503 5355
rect 12725 5321 12759 5355
rect 2973 5253 3007 5287
rect 9229 5253 9263 5287
rect 9321 5253 9355 5287
rect 10793 5253 10827 5287
rect 1409 5185 1443 5219
rect 1593 5185 1627 5219
rect 2054 5185 2088 5219
rect 2876 5185 2910 5219
rect 3065 5185 3099 5219
rect 3249 5185 3283 5219
rect 3612 5185 3646 5219
rect 3709 5185 3743 5219
rect 3801 5185 3835 5219
rect 3985 5185 4019 5219
rect 4445 5185 4479 5219
rect 4997 5185 5031 5219
rect 5180 5185 5214 5219
rect 5549 5185 5583 5219
rect 5825 5185 5859 5219
rect 6009 5185 6043 5219
rect 8309 5185 8343 5219
rect 8769 5185 8803 5219
rect 8953 5185 8987 5219
rect 10517 5185 10551 5219
rect 10609 5185 10643 5219
rect 10977 5185 11011 5219
rect 11069 5185 11103 5219
rect 11713 5185 11747 5219
rect 12541 5185 12575 5219
rect 2421 5117 2455 5151
rect 2513 5117 2547 5151
rect 4077 5117 4111 5151
rect 4629 5117 4663 5151
rect 5273 5117 5307 5151
rect 5365 5117 5399 5151
rect 5733 5117 5767 5151
rect 7941 5117 7975 5151
rect 8217 5117 8251 5151
rect 10425 5117 10459 5151
rect 11345 5117 11379 5151
rect 2697 5049 2731 5083
rect 5917 5049 5951 5083
rect 10609 5049 10643 5083
rect 11621 5049 11655 5083
rect 1685 4981 1719 5015
rect 3433 4981 3467 5015
rect 8401 4981 8435 5015
rect 10149 4981 10183 5015
rect 10333 4981 10367 5015
rect 11253 4981 11287 5015
rect 4445 4777 4479 4811
rect 6745 4777 6779 4811
rect 9689 4777 9723 4811
rect 2881 4709 2915 4743
rect 3893 4709 3927 4743
rect 7573 4709 7607 4743
rect 10057 4709 10091 4743
rect 12173 4709 12207 4743
rect 2329 4641 2363 4675
rect 3045 4641 3079 4675
rect 3525 4641 3559 4675
rect 6377 4641 6411 4675
rect 11069 4641 11103 4675
rect 1501 4573 1535 4607
rect 1777 4573 1811 4607
rect 2053 4573 2087 4607
rect 2237 4573 2271 4607
rect 2421 4573 2455 4607
rect 3157 4573 3191 4607
rect 3433 4573 3467 4607
rect 3801 4573 3835 4607
rect 4263 4573 4297 4607
rect 5181 4573 5215 4607
rect 5457 4573 5491 4607
rect 5641 4573 5675 4607
rect 5917 4573 5951 4607
rect 6469 4573 6503 4607
rect 6561 4573 6595 4607
rect 7205 4573 7239 4607
rect 9137 4573 9171 4607
rect 9505 4573 9539 4607
rect 9873 4573 9907 4607
rect 9965 4573 9999 4607
rect 10149 4573 10183 4607
rect 10701 4573 10735 4607
rect 10885 4573 10919 4607
rect 11161 4573 11195 4607
rect 11345 4573 11379 4607
rect 11621 4573 11655 4607
rect 11897 4573 11931 4607
rect 12009 4573 12043 4607
rect 5273 4505 5307 4539
rect 5365 4505 5399 4539
rect 7389 4505 7423 4539
rect 11529 4505 11563 4539
rect 2513 4437 2547 4471
rect 4261 4437 4295 4471
rect 4997 4437 5031 4471
rect 5733 4437 5767 4471
rect 8953 4437 8987 4471
rect 9413 4437 9447 4471
rect 3893 4233 3927 4267
rect 9597 4233 9631 4267
rect 9873 4233 9907 4267
rect 3525 4165 3559 4199
rect 3985 4165 4019 4199
rect 4629 4165 4663 4199
rect 6745 4165 6779 4199
rect 10885 4165 10919 4199
rect 11805 4165 11839 4199
rect 1777 4097 1811 4131
rect 1960 4097 1994 4131
rect 2145 4097 2179 4131
rect 2329 4097 2363 4131
rect 2605 4097 2639 4131
rect 3065 4097 3099 4131
rect 3249 4097 3283 4131
rect 3341 4097 3375 4131
rect 3709 4097 3743 4131
rect 6469 4097 6503 4131
rect 6653 4097 6687 4131
rect 6842 4097 6876 4131
rect 7389 4097 7423 4131
rect 7573 4097 7607 4131
rect 9965 4097 9999 4131
rect 10334 4097 10368 4131
rect 10529 4097 10563 4131
rect 10701 4097 10735 4131
rect 10977 4097 11011 4131
rect 11074 4097 11108 4131
rect 11529 4097 11563 4131
rect 2053 4029 2087 4063
rect 4353 4029 4387 4063
rect 7849 4029 7883 4063
rect 8125 4029 8159 4063
rect 10149 4029 10183 4063
rect 10241 4029 10275 4063
rect 13277 4029 13311 4063
rect 2513 3961 2547 3995
rect 7297 3961 7331 3995
rect 2697 3893 2731 3927
rect 6101 3893 6135 3927
rect 7021 3893 7055 3927
rect 7757 3893 7791 3927
rect 11253 3893 11287 3927
rect 3893 3689 3927 3723
rect 9045 3689 9079 3723
rect 9689 3689 9723 3723
rect 10057 3689 10091 3723
rect 12633 3689 12667 3723
rect 2421 3621 2455 3655
rect 3525 3621 3559 3655
rect 5733 3621 5767 3655
rect 2559 3553 2593 3587
rect 5365 3553 5399 3587
rect 5641 3553 5675 3587
rect 6653 3553 6687 3587
rect 6929 3553 6963 3587
rect 8401 3553 8435 3587
rect 9505 3553 9539 3587
rect 9597 3553 9631 3587
rect 9781 3553 9815 3587
rect 1868 3485 1902 3519
rect 1961 3485 1995 3519
rect 2053 3485 2087 3519
rect 2237 3485 2271 3519
rect 2329 3485 2363 3519
rect 2697 3485 2731 3519
rect 2973 3485 3007 3519
rect 3157 3485 3191 3519
rect 3249 3485 3283 3519
rect 3393 3485 3427 3519
rect 6009 3485 6043 3519
rect 9229 3485 9263 3519
rect 9321 3485 9355 3519
rect 9689 3485 9723 3519
rect 10241 3485 10275 3519
rect 12449 3485 12483 3519
rect 12725 3485 12759 3519
rect 1593 3417 1627 3451
rect 6101 3417 6135 3451
rect 10517 3417 10551 3451
rect 5917 3349 5951 3383
rect 6285 3349 6319 3383
rect 11989 3349 12023 3383
rect 12909 3349 12943 3383
rect 4721 3145 4755 3179
rect 5273 3145 5307 3179
rect 5549 3145 5583 3179
rect 10701 3145 10735 3179
rect 10977 3145 11011 3179
rect 3157 3077 3191 3111
rect 5191 3077 5225 3111
rect 5457 3077 5491 3111
rect 7297 3077 7331 3111
rect 10057 3077 10091 3111
rect 1593 3009 1627 3043
rect 1869 3009 1903 3043
rect 1961 3009 1995 3043
rect 2237 3009 2271 3043
rect 2421 3009 2455 3043
rect 2605 3009 2639 3043
rect 2881 3009 2915 3043
rect 3065 3009 3099 3043
rect 3893 3009 3927 3043
rect 4813 3009 4847 3043
rect 5089 3009 5123 3043
rect 5549 3009 5583 3043
rect 5641 3009 5675 3043
rect 5825 3009 5859 3043
rect 6469 3009 6503 3043
rect 6745 3009 6779 3043
rect 7200 3009 7234 3043
rect 7389 3009 7423 3043
rect 7573 3009 7607 3043
rect 9689 3009 9723 3043
rect 9873 3009 9907 3043
rect 10149 3009 10183 3043
rect 10293 3009 10327 3043
rect 10885 3009 10919 3043
rect 11069 3009 11103 3043
rect 11713 3009 11747 3043
rect 6101 2941 6135 2975
rect 6193 2941 6227 2975
rect 6837 2941 6871 2975
rect 9413 2941 9447 2975
rect 11253 2941 11287 2975
rect 11989 2941 12023 2975
rect 4905 2873 4939 2907
rect 7021 2873 7055 2907
rect 7941 2873 7975 2907
rect 10425 2873 10459 2907
rect 1777 2805 1811 2839
rect 2053 2805 2087 2839
rect 3985 2805 4019 2839
rect 13461 2805 13495 2839
rect 2973 2601 3007 2635
rect 3893 2601 3927 2635
rect 4445 2601 4479 2635
rect 7573 2601 7607 2635
rect 8585 2601 8619 2635
rect 9045 2601 9079 2635
rect 11897 2601 11931 2635
rect 2421 2533 2455 2567
rect 5089 2533 5123 2567
rect 8125 2533 8159 2567
rect 12725 2533 12759 2567
rect 1961 2465 1995 2499
rect 2605 2465 2639 2499
rect 3617 2465 3651 2499
rect 5457 2465 5491 2499
rect 5825 2465 5859 2499
rect 5917 2465 5951 2499
rect 6653 2465 6687 2499
rect 7113 2465 7147 2499
rect 9781 2465 9815 2499
rect 13277 2465 13311 2499
rect 1685 2397 1719 2431
rect 1868 2397 1902 2431
rect 2053 2397 2087 2431
rect 2237 2397 2271 2431
rect 2697 2397 2731 2431
rect 3137 2397 3171 2431
rect 3249 2397 3283 2431
rect 3801 2397 3835 2431
rect 4323 2397 4357 2431
rect 4629 2397 4663 2431
rect 5273 2397 5307 2431
rect 5549 2397 5583 2431
rect 5732 2397 5766 2431
rect 6101 2397 6135 2431
rect 6285 2397 6319 2431
rect 6561 2397 6595 2431
rect 7205 2397 7239 2431
rect 7695 2397 7729 2431
rect 8217 2397 8251 2431
rect 8769 2397 8803 2431
rect 9224 2397 9258 2431
rect 9320 2397 9354 2431
rect 9597 2397 9631 2431
rect 9689 2397 9723 2431
rect 9965 2397 9999 2431
rect 12081 2397 12115 2431
rect 12357 2397 12391 2431
rect 12889 2397 12923 2431
rect 13001 2397 13035 2431
rect 3525 2329 3559 2363
rect 4721 2329 4755 2363
rect 4905 2329 4939 2363
rect 6837 2329 6871 2363
rect 9413 2329 9447 2363
rect 10241 2329 10275 2363
rect 13369 2329 13403 2363
rect 4261 2261 4295 2295
rect 7757 2261 7791 2295
rect 11713 2261 11747 2295
rect 12541 2261 12575 2295
rect 3617 2057 3651 2091
rect 8125 2057 8159 2091
rect 10408 2057 10442 2091
rect 11069 2057 11103 2091
rect 5733 1989 5767 2023
rect 10701 1989 10735 2023
rect 3525 1921 3559 1955
rect 3893 1921 3927 1955
rect 4077 1921 4111 1955
rect 8401 1921 8435 1955
rect 10557 1921 10591 1955
rect 10793 1921 10827 1955
rect 10977 1921 11011 1955
rect 11253 1921 11287 1955
rect 1593 1853 1627 1887
rect 1869 1853 1903 1887
rect 6009 1853 6043 1887
rect 6377 1853 6411 1887
rect 6653 1853 6687 1887
rect 8677 1853 8711 1887
rect 10149 1853 10183 1887
rect 11529 1853 11563 1887
rect 11805 1853 11839 1887
rect 3341 1717 3375 1751
rect 4261 1717 4295 1751
rect 13277 1717 13311 1751
rect 2789 1513 2823 1547
rect 3893 1513 3927 1547
rect 5181 1513 5215 1547
rect 5365 1513 5399 1547
rect 6101 1513 6135 1547
rect 6653 1513 6687 1547
rect 7481 1513 7515 1547
rect 9597 1513 9631 1547
rect 11345 1513 11379 1547
rect 13461 1513 13495 1547
rect 8953 1445 8987 1479
rect 11713 1377 11747 1411
rect 11989 1377 12023 1411
rect 1777 1309 1811 1343
rect 2605 1309 2639 1343
rect 3433 1309 3467 1343
rect 3525 1309 3559 1343
rect 4025 1309 4059 1343
rect 4169 1309 4203 1343
rect 4445 1309 4479 1343
rect 5457 1309 5491 1343
rect 5549 1309 5583 1343
rect 5825 1309 5859 1343
rect 6193 1309 6227 1343
rect 6377 1309 6411 1343
rect 6561 1309 6595 1343
rect 7297 1309 7331 1343
rect 9413 1309 9447 1343
rect 11161 1309 11195 1343
rect 4261 1241 4295 1275
rect 9137 1241 9171 1275
rect 9321 1241 9355 1275
rect 1593 1173 1627 1207
rect 3525 1173 3559 1207
rect 5641 1173 5675 1207
<< metal1 >>
rect 3970 13744 3976 13796
rect 4028 13784 4034 13796
rect 7558 13784 7564 13796
rect 4028 13756 7564 13784
rect 4028 13744 4034 13756
rect 7558 13744 7564 13756
rect 7616 13744 7622 13796
rect 566 13676 572 13728
rect 624 13716 630 13728
rect 7190 13716 7196 13728
rect 624 13688 7196 13716
rect 624 13676 630 13688
rect 7190 13676 7196 13688
rect 7248 13676 7254 13728
rect 1104 13626 13892 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 12214 13626
rect 12266 13574 12278 13626
rect 12330 13574 12342 13626
rect 12394 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 13892 13626
rect 1104 13552 13892 13574
rect 5077 13515 5135 13521
rect 5077 13481 5089 13515
rect 5123 13512 5135 13515
rect 10229 13515 10287 13521
rect 10229 13512 10241 13515
rect 5123 13484 10241 13512
rect 5123 13481 5135 13484
rect 5077 13475 5135 13481
rect 10229 13481 10241 13484
rect 10275 13481 10287 13515
rect 10229 13475 10287 13481
rect 7653 13447 7711 13453
rect 2332 13416 6040 13444
rect 1394 13268 1400 13320
rect 1452 13308 1458 13320
rect 1857 13311 1915 13317
rect 1857 13308 1869 13311
rect 1452 13280 1869 13308
rect 1452 13268 1458 13280
rect 1857 13277 1869 13280
rect 1903 13277 1915 13311
rect 1857 13271 1915 13277
rect 2130 13268 2136 13320
rect 2188 13308 2194 13320
rect 2332 13308 2360 13416
rect 2409 13379 2467 13385
rect 2409 13345 2421 13379
rect 2455 13376 2467 13379
rect 3513 13379 3571 13385
rect 3513 13376 3525 13379
rect 2455 13348 3525 13376
rect 2455 13345 2467 13348
rect 2409 13339 2467 13345
rect 3513 13345 3525 13348
rect 3559 13345 3571 13379
rect 3513 13339 3571 13345
rect 4893 13379 4951 13385
rect 4893 13345 4905 13379
rect 4939 13376 4951 13379
rect 5905 13379 5963 13385
rect 5905 13376 5917 13379
rect 4939 13348 5917 13376
rect 4939 13345 4951 13348
rect 4893 13339 4951 13345
rect 5905 13345 5917 13348
rect 5951 13345 5963 13379
rect 5905 13339 5963 13345
rect 2501 13311 2559 13317
rect 2501 13308 2513 13311
rect 2188 13280 2513 13308
rect 2188 13268 2194 13280
rect 2501 13277 2513 13280
rect 2547 13277 2559 13311
rect 3326 13308 3332 13320
rect 2501 13271 2559 13277
rect 2976 13280 3188 13308
rect 3287 13280 3332 13308
rect 2317 13243 2375 13249
rect 2317 13209 2329 13243
rect 2363 13240 2375 13243
rect 2774 13240 2780 13252
rect 2363 13212 2780 13240
rect 2363 13209 2375 13212
rect 2317 13203 2375 13209
rect 2774 13200 2780 13212
rect 2832 13200 2838 13252
rect 2866 13200 2872 13252
rect 2924 13240 2930 13252
rect 2976 13249 3004 13280
rect 2961 13243 3019 13249
rect 2961 13240 2973 13243
rect 2924 13212 2973 13240
rect 2924 13200 2930 13212
rect 2961 13209 2973 13212
rect 3007 13209 3019 13243
rect 2961 13203 3019 13209
rect 3053 13243 3111 13249
rect 3053 13209 3065 13243
rect 3099 13209 3111 13243
rect 3160 13240 3188 13280
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 3602 13268 3608 13320
rect 3660 13308 3666 13320
rect 4341 13311 4399 13317
rect 4341 13308 4353 13311
rect 3660 13280 4353 13308
rect 3660 13268 3666 13280
rect 4341 13277 4353 13280
rect 4387 13277 4399 13311
rect 5074 13308 5080 13320
rect 4987 13280 5080 13308
rect 4341 13271 4399 13277
rect 5074 13268 5080 13280
rect 5132 13308 5138 13320
rect 5169 13311 5227 13317
rect 5169 13308 5181 13311
rect 5132 13280 5181 13308
rect 5132 13268 5138 13280
rect 5169 13277 5181 13280
rect 5215 13277 5227 13311
rect 5169 13271 5227 13277
rect 5629 13311 5687 13317
rect 5629 13277 5641 13311
rect 5675 13308 5687 13311
rect 5810 13308 5816 13320
rect 5675 13280 5816 13308
rect 5675 13277 5687 13280
rect 5629 13271 5687 13277
rect 5810 13268 5816 13280
rect 5868 13268 5874 13320
rect 6012 13308 6040 13416
rect 7653 13413 7665 13447
rect 7699 13413 7711 13447
rect 11517 13447 11575 13453
rect 11517 13444 11529 13447
rect 7653 13407 7711 13413
rect 9232 13416 11529 13444
rect 6914 13336 6920 13388
rect 6972 13376 6978 13388
rect 7009 13379 7067 13385
rect 7009 13376 7021 13379
rect 6972 13348 7021 13376
rect 6972 13336 6978 13348
rect 7009 13345 7021 13348
rect 7055 13345 7067 13379
rect 7190 13376 7196 13388
rect 7151 13348 7196 13376
rect 7009 13339 7067 13345
rect 7190 13336 7196 13348
rect 7248 13336 7254 13388
rect 7668 13376 7696 13407
rect 8018 13376 8024 13388
rect 7668 13348 8024 13376
rect 8018 13336 8024 13348
rect 8076 13376 8082 13388
rect 8941 13379 8999 13385
rect 8941 13376 8953 13379
rect 8076 13348 8953 13376
rect 8076 13336 8082 13348
rect 8941 13345 8953 13348
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 9232 13308 9260 13416
rect 11517 13413 11529 13416
rect 11563 13413 11575 13447
rect 11517 13407 11575 13413
rect 10781 13379 10839 13385
rect 10781 13345 10793 13379
rect 10827 13345 10839 13379
rect 10781 13339 10839 13345
rect 6012 13280 9260 13308
rect 9585 13311 9643 13317
rect 9585 13277 9597 13311
rect 9631 13308 9643 13311
rect 9674 13308 9680 13320
rect 9631 13280 9680 13308
rect 9631 13277 9643 13280
rect 9585 13271 9643 13277
rect 9674 13268 9680 13280
rect 9732 13268 9738 13320
rect 10796 13308 10824 13339
rect 10870 13336 10876 13388
rect 10928 13376 10934 13388
rect 11977 13379 12035 13385
rect 11977 13376 11989 13379
rect 10928 13348 11989 13376
rect 10928 13336 10934 13348
rect 11977 13345 11989 13348
rect 12023 13345 12035 13379
rect 11977 13339 12035 13345
rect 12161 13379 12219 13385
rect 12161 13345 12173 13379
rect 12207 13376 12219 13379
rect 12618 13376 12624 13388
rect 12207 13348 12624 13376
rect 12207 13345 12219 13348
rect 12161 13339 12219 13345
rect 10962 13308 10968 13320
rect 10796 13280 10968 13308
rect 10962 13268 10968 13280
rect 11020 13308 11026 13320
rect 12176 13308 12204 13339
rect 12618 13336 12624 13348
rect 12676 13336 12682 13388
rect 12342 13308 12348 13320
rect 11020 13280 12204 13308
rect 12303 13280 12348 13308
rect 11020 13268 11026 13280
rect 12342 13268 12348 13280
rect 12400 13268 12406 13320
rect 3421 13243 3479 13249
rect 3421 13240 3433 13243
rect 3160 13212 3433 13240
rect 3053 13203 3111 13209
rect 3421 13209 3433 13212
rect 3467 13209 3479 13243
rect 4798 13240 4804 13252
rect 4759 13212 4804 13240
rect 3421 13203 3479 13209
rect 3068 13172 3096 13203
rect 4798 13200 4804 13212
rect 4856 13200 4862 13252
rect 5721 13243 5779 13249
rect 5721 13209 5733 13243
rect 5767 13240 5779 13243
rect 6362 13240 6368 13252
rect 5767 13212 6368 13240
rect 5767 13209 5779 13212
rect 5721 13203 5779 13209
rect 6362 13200 6368 13212
rect 6420 13200 6426 13252
rect 9398 13240 9404 13252
rect 9359 13212 9404 13240
rect 9398 13200 9404 13212
rect 9456 13200 9462 13252
rect 9493 13243 9551 13249
rect 9493 13209 9505 13243
rect 9539 13240 9551 13243
rect 9858 13240 9864 13252
rect 9539 13212 9864 13240
rect 9539 13209 9551 13212
rect 9493 13203 9551 13209
rect 9858 13200 9864 13212
rect 9916 13200 9922 13252
rect 10042 13240 10048 13252
rect 10003 13212 10048 13240
rect 10042 13200 10048 13212
rect 10100 13200 10106 13252
rect 10134 13200 10140 13252
rect 10192 13240 10198 13252
rect 10689 13243 10747 13249
rect 10192 13212 10237 13240
rect 10192 13200 10198 13212
rect 10689 13209 10701 13243
rect 10735 13240 10747 13243
rect 12066 13240 12072 13252
rect 10735 13212 12072 13240
rect 10735 13209 10747 13212
rect 10689 13203 10747 13209
rect 12066 13200 12072 13212
rect 12124 13200 12130 13252
rect 12802 13240 12808 13252
rect 12763 13212 12808 13240
rect 12802 13200 12808 13212
rect 12860 13200 12866 13252
rect 12894 13200 12900 13252
rect 12952 13240 12958 13252
rect 12952 13212 12997 13240
rect 12952 13200 12958 13212
rect 3145 13175 3203 13181
rect 3145 13172 3157 13175
rect 3068 13144 3157 13172
rect 3145 13141 3157 13144
rect 3191 13141 3203 13175
rect 7282 13172 7288 13184
rect 7243 13144 7288 13172
rect 3145 13135 3203 13141
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 10594 13172 10600 13184
rect 10555 13144 10600 13172
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 11882 13172 11888 13184
rect 11843 13144 11888 13172
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 1104 13082 13892 13104
rect 1104 13030 8214 13082
rect 8266 13030 8278 13082
rect 8330 13030 8342 13082
rect 8394 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 13892 13082
rect 1104 13008 13892 13030
rect 1670 12928 1676 12980
rect 1728 12968 1734 12980
rect 6362 12968 6368 12980
rect 1728 12940 5948 12968
rect 6323 12940 6368 12968
rect 1728 12928 1734 12940
rect 2774 12860 2780 12912
rect 2832 12900 2838 12912
rect 2961 12903 3019 12909
rect 2961 12900 2973 12903
rect 2832 12872 2973 12900
rect 2832 12860 2838 12872
rect 2961 12869 2973 12872
rect 3007 12900 3019 12903
rect 3237 12903 3295 12909
rect 3237 12900 3249 12903
rect 3007 12872 3249 12900
rect 3007 12869 3019 12872
rect 2961 12863 3019 12869
rect 3237 12869 3249 12872
rect 3283 12869 3295 12903
rect 5810 12900 5816 12912
rect 5771 12872 5816 12900
rect 3237 12863 3295 12869
rect 5810 12860 5816 12872
rect 5868 12860 5874 12912
rect 5920 12900 5948 12940
rect 6362 12928 6368 12940
rect 6420 12928 6426 12980
rect 7377 12971 7435 12977
rect 7377 12937 7389 12971
rect 7423 12968 7435 12971
rect 12342 12968 12348 12980
rect 7423 12940 12348 12968
rect 7423 12937 7435 12940
rect 7377 12931 7435 12937
rect 6917 12903 6975 12909
rect 6917 12900 6929 12903
rect 5920 12872 6929 12900
rect 6917 12869 6929 12872
rect 6963 12869 6975 12903
rect 6917 12863 6975 12869
rect 7929 12903 7987 12909
rect 7929 12869 7941 12903
rect 7975 12900 7987 12903
rect 9950 12900 9956 12912
rect 7975 12872 9956 12900
rect 7975 12869 7987 12872
rect 7929 12863 7987 12869
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12832 2927 12835
rect 3326 12832 3332 12844
rect 2915 12804 3332 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 3513 12835 3571 12841
rect 3513 12801 3525 12835
rect 3559 12832 3571 12835
rect 3602 12832 3608 12844
rect 3559 12804 3608 12832
rect 3559 12801 3571 12804
rect 3513 12795 3571 12801
rect 3602 12792 3608 12804
rect 3660 12792 3666 12844
rect 4433 12835 4491 12841
rect 4433 12801 4445 12835
rect 4479 12801 4491 12835
rect 4433 12795 4491 12801
rect 3421 12767 3479 12773
rect 3421 12733 3433 12767
rect 3467 12764 3479 12767
rect 4448 12764 4476 12795
rect 5074 12792 5080 12844
rect 5132 12832 5138 12844
rect 5169 12835 5227 12841
rect 5169 12832 5181 12835
rect 5132 12804 5181 12832
rect 5132 12792 5138 12804
rect 5169 12801 5181 12804
rect 5215 12801 5227 12835
rect 5169 12795 5227 12801
rect 6089 12835 6147 12841
rect 6089 12801 6101 12835
rect 6135 12832 6147 12835
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6135 12804 6561 12832
rect 6135 12801 6147 12804
rect 6089 12795 6147 12801
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 7006 12832 7012 12844
rect 6967 12804 7012 12832
rect 6549 12795 6607 12801
rect 6104 12764 6132 12795
rect 7006 12792 7012 12804
rect 7064 12792 7070 12844
rect 7742 12832 7748 12844
rect 7703 12804 7748 12832
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 8018 12832 8024 12844
rect 7979 12804 8024 12832
rect 8018 12792 8024 12804
rect 8076 12792 8082 12844
rect 8956 12841 8984 12872
rect 9950 12860 9956 12872
rect 10008 12860 10014 12912
rect 10042 12860 10048 12912
rect 10100 12900 10106 12912
rect 10321 12903 10379 12909
rect 10321 12900 10333 12903
rect 10100 12872 10333 12900
rect 10100 12860 10106 12872
rect 10321 12869 10333 12872
rect 10367 12869 10379 12903
rect 10321 12863 10379 12869
rect 8941 12835 8999 12841
rect 8941 12801 8953 12835
rect 8987 12801 8999 12835
rect 9674 12832 9680 12844
rect 9635 12804 9680 12832
rect 8941 12795 8999 12801
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 9968 12832 9996 12860
rect 11900 12841 11928 12940
rect 12342 12928 12348 12940
rect 12400 12928 12406 12980
rect 10597 12835 10655 12841
rect 10597 12832 10609 12835
rect 9968 12804 10609 12832
rect 10597 12801 10609 12804
rect 10643 12801 10655 12835
rect 11609 12835 11667 12841
rect 11609 12832 11621 12835
rect 10597 12795 10655 12801
rect 10704 12804 11621 12832
rect 3467 12736 6132 12764
rect 6825 12767 6883 12773
rect 3467 12733 3479 12736
rect 3421 12727 3479 12733
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 6914 12764 6920 12776
rect 6871 12736 6920 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 6914 12724 6920 12736
rect 6972 12724 6978 12776
rect 9398 12724 9404 12776
rect 9456 12764 9462 12776
rect 9585 12767 9643 12773
rect 9585 12764 9597 12767
rect 9456 12736 9597 12764
rect 9456 12724 9462 12736
rect 9585 12733 9597 12736
rect 9631 12764 9643 12767
rect 10704 12764 10732 12804
rect 11609 12801 11621 12804
rect 11655 12801 11667 12835
rect 11609 12795 11667 12801
rect 11885 12835 11943 12841
rect 11885 12801 11897 12835
rect 11931 12801 11943 12835
rect 11885 12795 11943 12801
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 12805 12835 12863 12841
rect 12805 12832 12817 12835
rect 12768 12804 12817 12832
rect 12768 12792 12774 12804
rect 12805 12801 12817 12804
rect 12851 12801 12863 12835
rect 12805 12795 12863 12801
rect 9631 12736 10732 12764
rect 10781 12767 10839 12773
rect 9631 12733 9643 12736
rect 9585 12727 9643 12733
rect 10781 12733 10793 12767
rect 10827 12733 10839 12767
rect 11330 12764 11336 12776
rect 11291 12736 11336 12764
rect 10781 12727 10839 12733
rect 4798 12696 4804 12708
rect 4759 12668 4804 12696
rect 4798 12656 4804 12668
rect 4856 12656 4862 12708
rect 3878 12588 3884 12640
rect 3936 12628 3942 12640
rect 5718 12628 5724 12640
rect 3936 12600 5724 12628
rect 3936 12588 3942 12600
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 10796 12628 10824 12727
rect 11330 12724 11336 12736
rect 11388 12724 11394 12776
rect 11793 12767 11851 12773
rect 11793 12733 11805 12767
rect 11839 12764 11851 12767
rect 12728 12764 12756 12792
rect 11839 12736 12756 12764
rect 11839 12733 11851 12736
rect 11793 12727 11851 12733
rect 11241 12699 11299 12705
rect 11241 12665 11253 12699
rect 11287 12696 11299 12699
rect 12066 12696 12072 12708
rect 11287 12668 12072 12696
rect 11287 12665 11299 12668
rect 11241 12659 11299 12665
rect 12066 12656 12072 12668
rect 12124 12656 12130 12708
rect 12802 12656 12808 12708
rect 12860 12696 12866 12708
rect 13170 12696 13176 12708
rect 12860 12668 13176 12696
rect 12860 12656 12866 12668
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 11514 12628 11520 12640
rect 10796 12600 11520 12628
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 1104 12538 13892 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 12214 12538
rect 12266 12486 12278 12538
rect 12330 12486 12342 12538
rect 12394 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 13892 12538
rect 1104 12464 13892 12486
rect 3326 12424 3332 12436
rect 3287 12396 3332 12424
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 3602 12384 3608 12436
rect 3660 12424 3666 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3660 12396 3801 12424
rect 3660 12384 3666 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 6914 12424 6920 12436
rect 3789 12387 3847 12393
rect 5552 12396 6920 12424
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 4249 12291 4307 12297
rect 4249 12288 4261 12291
rect 4212 12260 4261 12288
rect 4212 12248 4218 12260
rect 4249 12257 4261 12260
rect 4295 12257 4307 12291
rect 4249 12251 4307 12257
rect 4338 12248 4344 12300
rect 4396 12288 4402 12300
rect 5552 12297 5580 12396
rect 6914 12384 6920 12396
rect 6972 12424 6978 12436
rect 6972 12396 8524 12424
rect 6972 12384 6978 12396
rect 6181 12359 6239 12365
rect 6181 12325 6193 12359
rect 6227 12325 6239 12359
rect 7742 12356 7748 12368
rect 7703 12328 7748 12356
rect 6181 12319 6239 12325
rect 5537 12291 5595 12297
rect 5537 12288 5549 12291
rect 4396 12260 5549 12288
rect 4396 12248 4402 12260
rect 5537 12257 5549 12260
rect 5583 12257 5595 12291
rect 5718 12288 5724 12300
rect 5679 12260 5724 12288
rect 5537 12251 5595 12257
rect 5718 12248 5724 12260
rect 5776 12248 5782 12300
rect 6196 12288 6224 12319
rect 7742 12316 7748 12328
rect 7800 12356 7806 12368
rect 8389 12359 8447 12365
rect 8389 12356 8401 12359
rect 7800 12328 8401 12356
rect 7800 12316 7806 12328
rect 8389 12325 8401 12328
rect 8435 12325 8447 12359
rect 8389 12319 8447 12325
rect 7929 12291 7987 12297
rect 7929 12288 7941 12291
rect 6196 12260 7941 12288
rect 2130 12220 2136 12232
rect 2091 12192 2136 12220
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 2866 12220 2872 12232
rect 2827 12192 2872 12220
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12220 3111 12223
rect 3326 12220 3332 12232
rect 3099 12192 3332 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 3326 12180 3332 12192
rect 3384 12180 3390 12232
rect 4798 12180 4804 12232
rect 4856 12220 4862 12232
rect 6288 12229 6316 12260
rect 7929 12257 7941 12260
rect 7975 12257 7987 12291
rect 8496 12288 8524 12396
rect 9674 12384 9680 12436
rect 9732 12424 9738 12436
rect 9861 12427 9919 12433
rect 9861 12424 9873 12427
rect 9732 12396 9873 12424
rect 9732 12384 9738 12396
rect 9861 12393 9873 12396
rect 9907 12393 9919 12427
rect 10134 12424 10140 12436
rect 10095 12396 10140 12424
rect 9861 12387 9919 12393
rect 10134 12384 10140 12396
rect 10192 12384 10198 12436
rect 11330 12384 11336 12436
rect 11388 12424 11394 12436
rect 12529 12427 12587 12433
rect 12529 12424 12541 12427
rect 11388 12396 12541 12424
rect 11388 12384 11394 12396
rect 12529 12393 12541 12396
rect 12575 12393 12587 12427
rect 12894 12424 12900 12436
rect 12855 12396 12900 12424
rect 12529 12387 12587 12393
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 14366 12356 14372 12368
rect 10888 12328 14372 12356
rect 9214 12288 9220 12300
rect 8496 12260 9220 12288
rect 7929 12251 7987 12257
rect 9214 12248 9220 12260
rect 9272 12248 9278 12300
rect 9401 12291 9459 12297
rect 9401 12257 9413 12291
rect 9447 12288 9459 12291
rect 10226 12288 10232 12300
rect 9447 12260 10232 12288
rect 9447 12257 9459 12260
rect 9401 12251 9459 12257
rect 10226 12248 10232 12260
rect 10284 12248 10290 12300
rect 10888 12297 10916 12328
rect 14366 12316 14372 12328
rect 14424 12316 14430 12368
rect 10873 12291 10931 12297
rect 10873 12257 10885 12291
rect 10919 12257 10931 12291
rect 10873 12251 10931 12257
rect 10962 12248 10968 12300
rect 11020 12288 11026 12300
rect 11020 12260 11113 12288
rect 11020 12248 11026 12260
rect 4985 12223 5043 12229
rect 4985 12220 4997 12223
rect 4856 12192 4997 12220
rect 4856 12180 4862 12192
rect 4985 12189 4997 12192
rect 5031 12189 5043 12223
rect 4985 12183 5043 12189
rect 6273 12223 6331 12229
rect 6273 12189 6285 12223
rect 6319 12189 6331 12223
rect 7466 12220 7472 12232
rect 7427 12192 7472 12220
rect 6273 12183 6331 12189
rect 7466 12180 7472 12192
rect 7524 12180 7530 12232
rect 9950 12220 9956 12232
rect 9911 12192 9956 12220
rect 9950 12180 9956 12192
rect 10008 12180 10014 12232
rect 10980 12220 11008 12248
rect 11514 12220 11520 12232
rect 10888 12192 11008 12220
rect 11475 12192 11520 12220
rect 3234 12152 3240 12164
rect 3195 12124 3240 12152
rect 3234 12112 3240 12124
rect 3292 12112 3298 12164
rect 4157 12155 4215 12161
rect 4157 12121 4169 12155
rect 4203 12152 4215 12155
rect 5718 12152 5724 12164
rect 4203 12124 5724 12152
rect 4203 12121 4215 12124
rect 4157 12115 4215 12121
rect 5718 12112 5724 12124
rect 5776 12112 5782 12164
rect 8481 12155 8539 12161
rect 8481 12121 8493 12155
rect 8527 12152 8539 12155
rect 8665 12155 8723 12161
rect 8665 12152 8677 12155
rect 8527 12124 8677 12152
rect 8527 12121 8539 12124
rect 8481 12115 8539 12121
rect 8665 12121 8677 12124
rect 8711 12121 8723 12155
rect 8665 12115 8723 12121
rect 9214 12112 9220 12164
rect 9272 12152 9278 12164
rect 10888 12152 10916 12192
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 12161 12223 12219 12229
rect 12161 12220 12173 12223
rect 12124 12192 12173 12220
rect 12124 12180 12130 12192
rect 12161 12189 12173 12192
rect 12207 12189 12219 12223
rect 12161 12183 12219 12189
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12220 12495 12223
rect 12710 12220 12716 12232
rect 12483 12192 12716 12220
rect 12483 12189 12495 12192
rect 12437 12183 12495 12189
rect 9272 12124 10916 12152
rect 12176 12152 12204 12183
rect 12710 12180 12716 12192
rect 12768 12180 12774 12232
rect 13170 12220 13176 12232
rect 13131 12192 13176 12220
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 12805 12155 12863 12161
rect 12805 12152 12817 12155
rect 12176 12124 12817 12152
rect 9272 12112 9278 12124
rect 12805 12121 12817 12124
rect 12851 12121 12863 12155
rect 12805 12115 12863 12121
rect 4890 12044 4896 12096
rect 4948 12084 4954 12096
rect 5077 12087 5135 12093
rect 5077 12084 5089 12087
rect 4948 12056 5089 12084
rect 4948 12044 4954 12056
rect 5077 12053 5089 12056
rect 5123 12053 5135 12087
rect 5077 12047 5135 12053
rect 5813 12087 5871 12093
rect 5813 12053 5825 12087
rect 5859 12084 5871 12087
rect 6362 12084 6368 12096
rect 5859 12056 6368 12084
rect 5859 12053 5871 12056
rect 5813 12047 5871 12053
rect 6362 12044 6368 12056
rect 6420 12044 6426 12096
rect 8570 12084 8576 12096
rect 8531 12056 8576 12084
rect 8570 12044 8576 12056
rect 8628 12044 8634 12096
rect 9030 12044 9036 12096
rect 9088 12084 9094 12096
rect 9493 12087 9551 12093
rect 9493 12084 9505 12087
rect 9088 12056 9505 12084
rect 9088 12044 9094 12056
rect 9493 12053 9505 12056
rect 9539 12053 9551 12087
rect 9493 12047 9551 12053
rect 9950 12044 9956 12096
rect 10008 12084 10014 12096
rect 10413 12087 10471 12093
rect 10413 12084 10425 12087
rect 10008 12056 10425 12084
rect 10008 12044 10014 12056
rect 10413 12053 10425 12056
rect 10459 12053 10471 12087
rect 10413 12047 10471 12053
rect 10781 12087 10839 12093
rect 10781 12053 10793 12087
rect 10827 12084 10839 12087
rect 11054 12084 11060 12096
rect 10827 12056 11060 12084
rect 10827 12053 10839 12056
rect 10781 12047 10839 12053
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 13265 12087 13323 12093
rect 13265 12053 13277 12087
rect 13311 12084 13323 12087
rect 13446 12084 13452 12096
rect 13311 12056 13452 12084
rect 13311 12053 13323 12056
rect 13265 12047 13323 12053
rect 13446 12044 13452 12056
rect 13504 12044 13510 12096
rect 1104 11994 13892 12016
rect 1104 11942 8214 11994
rect 8266 11942 8278 11994
rect 8330 11942 8342 11994
rect 8394 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 13892 11994
rect 1104 11920 13892 11942
rect 1394 11880 1400 11892
rect 1355 11852 1400 11880
rect 1394 11840 1400 11852
rect 1452 11840 1458 11892
rect 1765 11883 1823 11889
rect 1765 11849 1777 11883
rect 1811 11880 1823 11883
rect 3878 11880 3884 11892
rect 1811 11852 3884 11880
rect 1811 11849 1823 11852
rect 1765 11843 1823 11849
rect 3878 11840 3884 11852
rect 3936 11840 3942 11892
rect 4065 11883 4123 11889
rect 4065 11849 4077 11883
rect 4111 11880 4123 11883
rect 4154 11880 4160 11892
rect 4111 11852 4160 11880
rect 4111 11849 4123 11852
rect 4065 11843 4123 11849
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 5258 11840 5264 11892
rect 5316 11880 5322 11892
rect 5905 11883 5963 11889
rect 5905 11880 5917 11883
rect 5316 11852 5917 11880
rect 5316 11840 5322 11852
rect 5905 11849 5917 11852
rect 5951 11849 5963 11883
rect 9217 11883 9275 11889
rect 9217 11880 9229 11883
rect 5905 11843 5963 11849
rect 6012 11852 9229 11880
rect 2685 11815 2743 11821
rect 2685 11781 2697 11815
rect 2731 11812 2743 11815
rect 3234 11812 3240 11824
rect 2731 11784 3240 11812
rect 2731 11781 2743 11784
rect 2685 11775 2743 11781
rect 3234 11772 3240 11784
rect 3292 11772 3298 11824
rect 6012 11812 6040 11852
rect 9217 11849 9229 11852
rect 9263 11849 9275 11883
rect 9217 11843 9275 11849
rect 9677 11883 9735 11889
rect 9677 11849 9689 11883
rect 9723 11880 9735 11883
rect 9766 11880 9772 11892
rect 9723 11852 9772 11880
rect 9723 11849 9735 11852
rect 9677 11843 9735 11849
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 10042 11840 10048 11892
rect 10100 11880 10106 11892
rect 10229 11883 10287 11889
rect 10229 11880 10241 11883
rect 10100 11852 10241 11880
rect 10100 11840 10106 11852
rect 10229 11849 10241 11852
rect 10275 11849 10287 11883
rect 10229 11843 10287 11849
rect 4080 11784 6040 11812
rect 7745 11815 7803 11821
rect 2866 11744 2872 11756
rect 2779 11716 2872 11744
rect 2866 11704 2872 11716
rect 2924 11744 2930 11756
rect 4080 11744 4108 11784
rect 7745 11781 7757 11815
rect 7791 11812 7803 11815
rect 8570 11812 8576 11824
rect 7791 11784 8576 11812
rect 7791 11781 7803 11784
rect 7745 11775 7803 11781
rect 8570 11772 8576 11784
rect 8628 11772 8634 11824
rect 9950 11812 9956 11824
rect 9048 11784 9956 11812
rect 2924 11716 4108 11744
rect 4157 11747 4215 11753
rect 2924 11704 2930 11716
rect 4157 11713 4169 11747
rect 4203 11744 4215 11747
rect 5626 11744 5632 11756
rect 4203 11716 5632 11744
rect 4203 11713 4215 11716
rect 4157 11707 4215 11713
rect 5626 11704 5632 11716
rect 5684 11704 5690 11756
rect 6089 11747 6147 11753
rect 6089 11744 6101 11747
rect 5735 11716 6101 11744
rect 1854 11676 1860 11688
rect 1815 11648 1860 11676
rect 1854 11636 1860 11648
rect 1912 11636 1918 11688
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11645 2007 11679
rect 2222 11676 2228 11688
rect 2183 11648 2228 11676
rect 1949 11639 2007 11645
rect 1486 11568 1492 11620
rect 1544 11608 1550 11620
rect 1964 11608 1992 11639
rect 2222 11636 2228 11648
rect 2280 11636 2286 11688
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 3418 11676 3424 11688
rect 2832 11648 2877 11676
rect 3379 11648 3424 11676
rect 2832 11636 2838 11648
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 3881 11679 3939 11685
rect 3881 11645 3893 11679
rect 3927 11676 3939 11679
rect 4338 11676 4344 11688
rect 3927 11648 4344 11676
rect 3927 11645 3939 11648
rect 3881 11639 3939 11645
rect 3326 11608 3332 11620
rect 1544 11580 1992 11608
rect 3287 11580 3332 11608
rect 1544 11568 1550 11580
rect 1964 11540 1992 11580
rect 3326 11568 3332 11580
rect 3384 11568 3390 11620
rect 3896 11540 3924 11639
rect 4338 11636 4344 11648
rect 4396 11636 4402 11688
rect 4617 11679 4675 11685
rect 4617 11676 4629 11679
rect 4540 11648 4629 11676
rect 1964 11512 3924 11540
rect 3970 11500 3976 11552
rect 4028 11540 4034 11552
rect 4540 11549 4568 11648
rect 4617 11645 4629 11648
rect 4663 11645 4675 11679
rect 5166 11676 5172 11688
rect 5127 11648 5172 11676
rect 4617 11639 4675 11645
rect 5166 11636 5172 11648
rect 5224 11636 5230 11688
rect 5258 11636 5264 11688
rect 5316 11676 5322 11688
rect 5316 11648 5361 11676
rect 5316 11636 5322 11648
rect 4982 11568 4988 11620
rect 5040 11608 5046 11620
rect 5077 11611 5135 11617
rect 5077 11608 5089 11611
rect 5040 11580 5089 11608
rect 5040 11568 5046 11580
rect 5077 11577 5089 11580
rect 5123 11577 5135 11611
rect 5350 11608 5356 11620
rect 5311 11580 5356 11608
rect 5077 11571 5135 11577
rect 5350 11568 5356 11580
rect 5408 11568 5414 11620
rect 4525 11543 4583 11549
rect 4525 11540 4537 11543
rect 4028 11512 4537 11540
rect 4028 11500 4034 11512
rect 4525 11509 4537 11512
rect 4571 11509 4583 11543
rect 4525 11503 4583 11509
rect 4890 11500 4896 11552
rect 4948 11540 4954 11552
rect 5735 11540 5763 11716
rect 6089 11713 6101 11716
rect 6135 11713 6147 11747
rect 6089 11707 6147 11713
rect 6181 11747 6239 11753
rect 6181 11713 6193 11747
rect 6227 11744 6239 11747
rect 6365 11747 6423 11753
rect 6365 11744 6377 11747
rect 6227 11716 6377 11744
rect 6227 11713 6239 11716
rect 6181 11707 6239 11713
rect 6365 11713 6377 11716
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 6454 11704 6460 11756
rect 6512 11744 6518 11756
rect 6641 11747 6699 11753
rect 6641 11744 6653 11747
rect 6512 11716 6653 11744
rect 6512 11704 6518 11716
rect 6641 11713 6653 11716
rect 6687 11713 6699 11747
rect 7098 11744 7104 11756
rect 7059 11716 7104 11744
rect 6641 11707 6699 11713
rect 7098 11704 7104 11716
rect 7156 11704 7162 11756
rect 7285 11747 7343 11753
rect 7285 11713 7297 11747
rect 7331 11744 7343 11747
rect 7466 11744 7472 11756
rect 7331 11716 7472 11744
rect 7331 11713 7343 11716
rect 7285 11707 7343 11713
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 9048 11753 9076 11784
rect 9950 11772 9956 11784
rect 10008 11772 10014 11824
rect 10318 11772 10324 11824
rect 10376 11812 10382 11824
rect 12437 11815 12495 11821
rect 10376 11784 11744 11812
rect 10376 11772 10382 11784
rect 8389 11747 8447 11753
rect 8389 11713 8401 11747
rect 8435 11744 8447 11747
rect 9033 11747 9091 11753
rect 9033 11744 9045 11747
rect 8435 11716 9045 11744
rect 8435 11713 8447 11716
rect 8389 11707 8447 11713
rect 9033 11713 9045 11716
rect 9079 11713 9091 11747
rect 9033 11707 9091 11713
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11744 9643 11747
rect 10134 11744 10140 11756
rect 9631 11716 10140 11744
rect 9631 11713 9643 11716
rect 9585 11707 9643 11713
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 10410 11704 10416 11756
rect 10468 11744 10474 11756
rect 10689 11747 10747 11753
rect 10689 11744 10701 11747
rect 10468 11716 10701 11744
rect 10468 11704 10474 11716
rect 10689 11713 10701 11716
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 10778 11704 10784 11756
rect 10836 11744 10842 11756
rect 11716 11753 11744 11784
rect 12437 11781 12449 11815
rect 12483 11812 12495 11815
rect 13446 11812 13452 11824
rect 12483 11784 13308 11812
rect 13407 11784 13452 11812
rect 12483 11781 12495 11784
rect 12437 11775 12495 11781
rect 13280 11756 13308 11784
rect 13446 11772 13452 11784
rect 13504 11772 13510 11824
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 10836 11716 11529 11744
rect 10836 11704 10842 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 12529 11747 12587 11753
rect 12529 11713 12541 11747
rect 12575 11744 12587 11747
rect 12986 11744 12992 11756
rect 12575 11716 12992 11744
rect 12575 11713 12587 11716
rect 12529 11707 12587 11713
rect 12986 11704 12992 11716
rect 13044 11704 13050 11756
rect 13262 11744 13268 11756
rect 13223 11716 13268 11744
rect 13262 11704 13268 11716
rect 13320 11704 13326 11756
rect 5810 11636 5816 11688
rect 5868 11676 5874 11688
rect 5868 11648 6592 11676
rect 5868 11636 5874 11648
rect 6086 11568 6092 11620
rect 6144 11608 6150 11620
rect 6457 11611 6515 11617
rect 6457 11608 6469 11611
rect 6144 11580 6469 11608
rect 6144 11568 6150 11580
rect 6457 11577 6469 11580
rect 6503 11577 6515 11611
rect 6564 11608 6592 11648
rect 8294 11636 8300 11688
rect 8352 11676 8358 11688
rect 8481 11679 8539 11685
rect 8481 11676 8493 11679
rect 8352 11648 8493 11676
rect 8352 11636 8358 11648
rect 8481 11645 8493 11648
rect 8527 11645 8539 11679
rect 8481 11639 8539 11645
rect 9214 11636 9220 11688
rect 9272 11676 9278 11688
rect 9490 11676 9496 11688
rect 9272 11648 9496 11676
rect 9272 11636 9278 11648
rect 9490 11636 9496 11648
rect 9548 11676 9554 11688
rect 9769 11679 9827 11685
rect 9769 11676 9781 11679
rect 9548 11648 9781 11676
rect 9548 11636 9554 11648
rect 9769 11645 9781 11648
rect 9815 11645 9827 11679
rect 10502 11676 10508 11688
rect 10463 11648 10508 11676
rect 9769 11639 9827 11645
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 13078 11676 13084 11688
rect 10796 11648 13084 11676
rect 8938 11608 8944 11620
rect 6564 11580 8944 11608
rect 6457 11571 6515 11577
rect 8938 11568 8944 11580
rect 8996 11568 9002 11620
rect 9858 11568 9864 11620
rect 9916 11608 9922 11620
rect 10137 11611 10195 11617
rect 10137 11608 10149 11611
rect 9916 11580 10149 11608
rect 9916 11568 9922 11580
rect 10137 11577 10149 11580
rect 10183 11577 10195 11611
rect 10137 11571 10195 11577
rect 4948 11512 5763 11540
rect 4948 11500 4954 11512
rect 5902 11500 5908 11552
rect 5960 11540 5966 11552
rect 6181 11543 6239 11549
rect 6181 11540 6193 11543
rect 5960 11512 6193 11540
rect 5960 11500 5966 11512
rect 6181 11509 6193 11512
rect 6227 11509 6239 11543
rect 6181 11503 6239 11509
rect 6730 11500 6736 11552
rect 6788 11540 6794 11552
rect 6825 11543 6883 11549
rect 6825 11540 6837 11543
rect 6788 11512 6837 11540
rect 6788 11500 6794 11512
rect 6825 11509 6837 11512
rect 6871 11509 6883 11543
rect 6825 11503 6883 11509
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 10796 11540 10824 11648
rect 13078 11636 13084 11648
rect 13136 11636 13142 11688
rect 11054 11568 11060 11620
rect 11112 11608 11118 11620
rect 11609 11611 11667 11617
rect 11609 11608 11621 11611
rect 11112 11580 11621 11608
rect 11112 11568 11118 11580
rect 11609 11577 11621 11580
rect 11655 11577 11667 11611
rect 11609 11571 11667 11577
rect 9456 11512 10824 11540
rect 9456 11500 9462 11512
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11149 11543 11207 11549
rect 11149 11540 11161 11543
rect 10928 11512 11161 11540
rect 10928 11500 10934 11512
rect 11149 11509 11161 11512
rect 11195 11509 11207 11543
rect 11149 11503 11207 11509
rect 12345 11543 12403 11549
rect 12345 11509 12357 11543
rect 12391 11540 12403 11543
rect 12894 11540 12900 11552
rect 12391 11512 12900 11540
rect 12391 11509 12403 11512
rect 12345 11503 12403 11509
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 1104 11450 13892 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 12214 11450
rect 12266 11398 12278 11450
rect 12330 11398 12342 11450
rect 12394 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 13892 11450
rect 1104 11376 13892 11398
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 3329 11339 3387 11345
rect 3329 11336 3341 11339
rect 2832 11308 3341 11336
rect 2832 11296 2838 11308
rect 3329 11305 3341 11308
rect 3375 11305 3387 11339
rect 3329 11299 3387 11305
rect 5626 11296 5632 11348
rect 5684 11336 5690 11348
rect 5813 11339 5871 11345
rect 5813 11336 5825 11339
rect 5684 11308 5825 11336
rect 5684 11296 5690 11308
rect 5813 11305 5825 11308
rect 5859 11305 5871 11339
rect 7098 11336 7104 11348
rect 5813 11299 5871 11305
rect 6104 11308 7104 11336
rect 3053 11271 3111 11277
rect 3053 11237 3065 11271
rect 3099 11268 3111 11271
rect 3234 11268 3240 11280
rect 3099 11240 3240 11268
rect 3099 11237 3111 11240
rect 3053 11231 3111 11237
rect 3234 11228 3240 11240
rect 3292 11228 3298 11280
rect 4982 11228 4988 11280
rect 5040 11268 5046 11280
rect 5258 11268 5264 11280
rect 5040 11240 5264 11268
rect 5040 11228 5046 11240
rect 5258 11228 5264 11240
rect 5316 11268 5322 11280
rect 6104 11268 6132 11308
rect 7098 11296 7104 11308
rect 7156 11296 7162 11348
rect 8294 11336 8300 11348
rect 8255 11308 8300 11336
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 8938 11336 8944 11348
rect 8899 11308 8944 11336
rect 8938 11296 8944 11308
rect 8996 11296 9002 11348
rect 10134 11336 10140 11348
rect 10095 11308 10140 11336
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 11146 11336 11152 11348
rect 10520 11308 11152 11336
rect 5316 11240 6132 11268
rect 6181 11271 6239 11277
rect 5316 11228 5322 11240
rect 6181 11237 6193 11271
rect 6227 11268 6239 11271
rect 6822 11268 6828 11280
rect 6227 11240 6828 11268
rect 6227 11237 6239 11240
rect 6181 11231 6239 11237
rect 6822 11228 6828 11240
rect 6880 11228 6886 11280
rect 7193 11271 7251 11277
rect 7193 11237 7205 11271
rect 7239 11268 7251 11271
rect 10520 11268 10548 11308
rect 11146 11296 11152 11308
rect 11204 11296 11210 11348
rect 11241 11339 11299 11345
rect 11241 11305 11253 11339
rect 11287 11336 11299 11339
rect 11882 11336 11888 11348
rect 11287 11308 11888 11336
rect 11287 11305 11299 11308
rect 11241 11299 11299 11305
rect 11882 11296 11888 11308
rect 11940 11296 11946 11348
rect 11422 11268 11428 11280
rect 7239 11240 10548 11268
rect 10612 11240 11428 11268
rect 7239 11237 7251 11240
rect 7193 11231 7251 11237
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 6454 11200 6460 11212
rect 3936 11172 6460 11200
rect 3936 11160 3942 11172
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11132 1639 11135
rect 2222 11132 2228 11144
rect 1627 11104 2228 11132
rect 1627 11101 1639 11104
rect 1581 11095 1639 11101
rect 2222 11092 2228 11104
rect 2280 11092 2286 11144
rect 3050 11132 3056 11144
rect 3011 11104 3056 11132
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 3326 11132 3332 11144
rect 3283 11104 3332 11132
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 3970 11132 3976 11144
rect 3931 11104 3976 11132
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 4522 11092 4528 11144
rect 4580 11132 4586 11144
rect 4890 11132 4896 11144
rect 4580 11104 4896 11132
rect 4580 11092 4586 11104
rect 4890 11092 4896 11104
rect 4948 11092 4954 11144
rect 5902 11092 5908 11144
rect 5960 11132 5966 11144
rect 5997 11135 6055 11141
rect 5997 11132 6009 11135
rect 5960 11104 6009 11132
rect 5960 11092 5966 11104
rect 5997 11101 6009 11104
rect 6043 11101 6055 11135
rect 5997 11095 6055 11101
rect 6086 11092 6092 11144
rect 6144 11132 6150 11144
rect 6288 11141 6316 11172
rect 6454 11160 6460 11172
rect 6512 11160 6518 11212
rect 6549 11203 6607 11209
rect 6549 11169 6561 11203
rect 6595 11200 6607 11203
rect 7834 11200 7840 11212
rect 6595 11172 7840 11200
rect 6595 11169 6607 11172
rect 6549 11163 6607 11169
rect 6273 11135 6331 11141
rect 6144 11104 6189 11132
rect 6144 11092 6150 11104
rect 6273 11101 6285 11135
rect 6319 11101 6331 11135
rect 6273 11095 6331 11101
rect 5442 11024 5448 11076
rect 5500 11064 5506 11076
rect 6564 11064 6592 11163
rect 7834 11160 7840 11172
rect 7892 11160 7898 11212
rect 9398 11200 9404 11212
rect 8404 11172 8708 11200
rect 9359 11172 9404 11200
rect 7466 11092 7472 11144
rect 7524 11132 7530 11144
rect 8404 11141 8432 11172
rect 8113 11135 8171 11141
rect 8113 11132 8125 11135
rect 7524 11104 8125 11132
rect 7524 11092 7530 11104
rect 8113 11101 8125 11104
rect 8159 11101 8171 11135
rect 8113 11095 8171 11101
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 8570 11132 8576 11144
rect 8531 11104 8576 11132
rect 8389 11095 8447 11101
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 8680 11132 8708 11172
rect 9398 11160 9404 11172
rect 9456 11160 9462 11212
rect 9490 11160 9496 11212
rect 9548 11200 9554 11212
rect 9548 11172 9593 11200
rect 9548 11160 9554 11172
rect 10226 11160 10232 11212
rect 10284 11200 10290 11212
rect 10413 11203 10471 11209
rect 10413 11200 10425 11203
rect 10284 11172 10425 11200
rect 10284 11160 10290 11172
rect 10413 11169 10425 11172
rect 10459 11169 10471 11203
rect 10413 11163 10471 11169
rect 9858 11132 9864 11144
rect 8680 11104 9864 11132
rect 9858 11092 9864 11104
rect 9916 11132 9922 11144
rect 10318 11132 10324 11144
rect 9916 11104 10324 11132
rect 9916 11092 9922 11104
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 10612 11141 10640 11240
rect 11422 11228 11428 11240
rect 11480 11228 11486 11280
rect 12802 11268 12808 11280
rect 12763 11240 12808 11268
rect 12802 11228 12808 11240
rect 12860 11228 12866 11280
rect 10870 11200 10876 11212
rect 10831 11172 10876 11200
rect 10870 11160 10876 11172
rect 10928 11160 10934 11212
rect 10505 11135 10563 11141
rect 10505 11101 10517 11135
rect 10551 11101 10563 11135
rect 10505 11095 10563 11101
rect 10597 11135 10655 11141
rect 10597 11101 10609 11135
rect 10643 11101 10655 11135
rect 10597 11095 10655 11101
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11101 10839 11135
rect 11054 11132 11060 11144
rect 11015 11104 11060 11132
rect 10781 11095 10839 11101
rect 5500 11036 6592 11064
rect 6733 11067 6791 11073
rect 5500 11024 5506 11036
rect 6733 11033 6745 11067
rect 6779 11033 6791 11067
rect 6733 11027 6791 11033
rect 6825 11067 6883 11073
rect 6825 11033 6837 11067
rect 6871 11064 6883 11067
rect 6914 11064 6920 11076
rect 6871 11036 6920 11064
rect 6871 11033 6883 11036
rect 6825 11027 6883 11033
rect 2958 10956 2964 11008
rect 3016 10996 3022 11008
rect 6748 10996 6776 11027
rect 6914 11024 6920 11036
rect 6972 11024 6978 11076
rect 8757 11067 8815 11073
rect 8757 11033 8769 11067
rect 8803 11064 8815 11067
rect 9309 11067 9367 11073
rect 9309 11064 9321 11067
rect 8803 11036 9321 11064
rect 8803 11033 8815 11036
rect 8757 11027 8815 11033
rect 9309 11033 9321 11036
rect 9355 11033 9367 11067
rect 9309 11027 9367 11033
rect 3016 10968 6776 10996
rect 10520 10996 10548 11095
rect 10796 11064 10824 11095
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 11146 11092 11152 11144
rect 11204 11132 11210 11144
rect 11517 11135 11575 11141
rect 11517 11132 11529 11135
rect 11204 11104 11529 11132
rect 11204 11092 11210 11104
rect 11517 11101 11529 11104
rect 11563 11132 11575 11135
rect 12342 11132 12348 11144
rect 11563 11104 12348 11132
rect 11563 11101 11575 11104
rect 11517 11095 11575 11101
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 12989 11135 13047 11141
rect 12989 11101 13001 11135
rect 13035 11132 13047 11135
rect 13173 11135 13231 11141
rect 13173 11132 13185 11135
rect 13035 11104 13185 11132
rect 13035 11101 13047 11104
rect 12989 11095 13047 11101
rect 13173 11101 13185 11104
rect 13219 11132 13231 11135
rect 13446 11132 13452 11144
rect 13219 11104 13452 11132
rect 13219 11101 13231 11104
rect 13173 11095 13231 11101
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 10796 11036 11100 11064
rect 11072 11008 11100 11036
rect 10962 10996 10968 11008
rect 10520 10968 10968 10996
rect 3016 10956 3022 10968
rect 10962 10956 10968 10968
rect 11020 10956 11026 11008
rect 11054 10956 11060 11008
rect 11112 10956 11118 11008
rect 13354 10996 13360 11008
rect 13315 10968 13360 10996
rect 13354 10956 13360 10968
rect 13412 10956 13418 11008
rect 1104 10906 13892 10928
rect 1104 10854 8214 10906
rect 8266 10854 8278 10906
rect 8330 10854 8342 10906
rect 8394 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 13892 10906
rect 1104 10832 13892 10854
rect 2133 10795 2191 10801
rect 2133 10761 2145 10795
rect 2179 10792 2191 10795
rect 2222 10792 2228 10804
rect 2179 10764 2228 10792
rect 2179 10761 2191 10764
rect 2133 10755 2191 10761
rect 2222 10752 2228 10764
rect 2280 10752 2286 10804
rect 3418 10752 3424 10804
rect 3476 10792 3482 10804
rect 3605 10795 3663 10801
rect 3605 10792 3617 10795
rect 3476 10764 3617 10792
rect 3476 10752 3482 10764
rect 3605 10761 3617 10764
rect 3651 10761 3663 10795
rect 3605 10755 3663 10761
rect 4341 10795 4399 10801
rect 4341 10761 4353 10795
rect 4387 10792 4399 10795
rect 5166 10792 5172 10804
rect 4387 10764 5172 10792
rect 4387 10761 4399 10764
rect 4341 10755 4399 10761
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 5810 10752 5816 10804
rect 5868 10752 5874 10804
rect 6178 10752 6184 10804
rect 6236 10792 6242 10804
rect 10318 10792 10324 10804
rect 6236 10764 10324 10792
rect 6236 10752 6242 10764
rect 3326 10724 3332 10736
rect 3287 10696 3332 10724
rect 3326 10684 3332 10696
rect 3384 10684 3390 10736
rect 4433 10727 4491 10733
rect 4433 10693 4445 10727
rect 4479 10724 4491 10727
rect 4801 10727 4859 10733
rect 4801 10724 4813 10727
rect 4479 10696 4813 10724
rect 4479 10693 4491 10696
rect 4433 10687 4491 10693
rect 4801 10693 4813 10696
rect 4847 10724 4859 10727
rect 5350 10724 5356 10736
rect 4847 10696 5356 10724
rect 4847 10693 4859 10696
rect 4801 10687 4859 10693
rect 5350 10684 5356 10696
rect 5408 10684 5414 10736
rect 5828 10724 5856 10752
rect 6362 10724 6368 10736
rect 5460 10696 5856 10724
rect 6323 10696 6368 10724
rect 1670 10656 1676 10668
rect 1631 10628 1676 10656
rect 1670 10616 1676 10628
rect 1728 10616 1734 10668
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10625 1823 10659
rect 1765 10619 1823 10625
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10656 2651 10659
rect 2866 10656 2872 10668
rect 2639 10628 2872 10656
rect 2639 10625 2651 10628
rect 2593 10619 2651 10625
rect 1486 10588 1492 10600
rect 1447 10560 1492 10588
rect 1486 10548 1492 10560
rect 1544 10548 1550 10600
rect 1780 10520 1808 10619
rect 2866 10616 2872 10628
rect 2924 10616 2930 10668
rect 3050 10616 3056 10668
rect 3108 10656 3114 10668
rect 3513 10659 3571 10665
rect 3513 10656 3525 10659
rect 3108 10628 3525 10656
rect 3108 10616 3114 10628
rect 3513 10625 3525 10628
rect 3559 10656 3571 10659
rect 3789 10659 3847 10665
rect 3789 10656 3801 10659
rect 3559 10628 3801 10656
rect 3559 10625 3571 10628
rect 3513 10619 3571 10625
rect 3789 10625 3801 10628
rect 3835 10625 3847 10659
rect 4522 10656 4528 10668
rect 4483 10628 4528 10656
rect 3789 10619 3847 10625
rect 4522 10616 4528 10628
rect 4580 10616 4586 10668
rect 5460 10665 5488 10696
rect 6362 10684 6368 10696
rect 6420 10684 6426 10736
rect 6564 10733 6592 10764
rect 6549 10727 6607 10733
rect 6549 10693 6561 10727
rect 6595 10693 6607 10727
rect 6549 10687 6607 10693
rect 6638 10684 6644 10736
rect 6696 10724 6702 10736
rect 6733 10727 6791 10733
rect 6733 10724 6745 10727
rect 6696 10696 6745 10724
rect 6696 10684 6702 10696
rect 6733 10693 6745 10696
rect 6779 10724 6791 10727
rect 7742 10724 7748 10736
rect 6779 10696 7748 10724
rect 6779 10693 6791 10696
rect 6733 10687 6791 10693
rect 5445 10659 5503 10665
rect 5445 10625 5457 10659
rect 5491 10625 5503 10659
rect 5810 10656 5816 10668
rect 5771 10628 5816 10656
rect 5445 10619 5503 10625
rect 5810 10616 5816 10628
rect 5868 10616 5874 10668
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10656 5963 10659
rect 5994 10656 6000 10668
rect 5951 10628 6000 10656
rect 5951 10625 5963 10628
rect 5905 10619 5963 10625
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 6089 10659 6147 10665
rect 6089 10625 6101 10659
rect 6135 10656 6147 10659
rect 6454 10656 6460 10668
rect 6135 10628 6460 10656
rect 6135 10625 6147 10628
rect 6089 10619 6147 10625
rect 6454 10616 6460 10628
rect 6512 10616 6518 10668
rect 7098 10656 7104 10668
rect 7059 10628 7104 10656
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 7190 10616 7196 10668
rect 7248 10656 7254 10668
rect 7392 10665 7420 10696
rect 7742 10684 7748 10696
rect 7800 10684 7806 10736
rect 7929 10727 7987 10733
rect 7929 10693 7941 10727
rect 7975 10724 7987 10727
rect 8757 10727 8815 10733
rect 8757 10724 8769 10727
rect 7975 10696 8769 10724
rect 7975 10693 7987 10696
rect 7929 10687 7987 10693
rect 8757 10693 8769 10696
rect 8803 10693 8815 10727
rect 8757 10687 8815 10693
rect 7377 10659 7435 10665
rect 7248 10628 7293 10656
rect 7248 10616 7254 10628
rect 7377 10625 7389 10659
rect 7423 10625 7435 10659
rect 7377 10619 7435 10625
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 7616 10628 7849 10656
rect 7616 10616 7622 10628
rect 7837 10625 7849 10628
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10625 8447 10659
rect 8389 10619 8447 10625
rect 7653 10591 7711 10597
rect 7653 10557 7665 10591
rect 7699 10557 7711 10591
rect 7653 10551 7711 10557
rect 5902 10520 5908 10532
rect 1780 10492 5908 10520
rect 5902 10480 5908 10492
rect 5960 10480 5966 10532
rect 5997 10523 6055 10529
rect 5997 10489 6009 10523
rect 6043 10520 6055 10523
rect 6086 10520 6092 10532
rect 6043 10492 6092 10520
rect 6043 10489 6055 10492
rect 5997 10483 6055 10489
rect 6086 10480 6092 10492
rect 6144 10480 6150 10532
rect 6917 10523 6975 10529
rect 6917 10489 6929 10523
rect 6963 10520 6975 10523
rect 7006 10520 7012 10532
rect 6963 10492 7012 10520
rect 6963 10489 6975 10492
rect 6917 10483 6975 10489
rect 7006 10480 7012 10492
rect 7064 10480 7070 10532
rect 7285 10523 7343 10529
rect 7285 10489 7297 10523
rect 7331 10520 7343 10523
rect 7558 10520 7564 10532
rect 7331 10492 7564 10520
rect 7331 10489 7343 10492
rect 7285 10483 7343 10489
rect 7558 10480 7564 10492
rect 7616 10480 7622 10532
rect 7668 10520 7696 10551
rect 7742 10548 7748 10600
rect 7800 10588 7806 10600
rect 8404 10588 8432 10619
rect 8478 10616 8484 10668
rect 8536 10656 8542 10668
rect 8573 10659 8631 10665
rect 8573 10656 8585 10659
rect 8536 10628 8585 10656
rect 8536 10616 8542 10628
rect 8573 10625 8585 10628
rect 8619 10656 8631 10659
rect 9769 10659 9827 10665
rect 8619 10628 9674 10656
rect 8619 10625 8631 10628
rect 8573 10619 8631 10625
rect 9646 10600 9674 10628
rect 9769 10625 9781 10659
rect 9815 10656 9827 10659
rect 10042 10656 10048 10668
rect 9815 10628 10048 10656
rect 9815 10625 9827 10628
rect 9769 10619 9827 10625
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 10152 10665 10180 10764
rect 10318 10752 10324 10764
rect 10376 10792 10382 10804
rect 11054 10792 11060 10804
rect 10376 10764 10916 10792
rect 11015 10764 11060 10792
rect 10376 10752 10382 10764
rect 10226 10684 10232 10736
rect 10284 10724 10290 10736
rect 10284 10696 10732 10724
rect 10284 10684 10290 10696
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10625 10195 10659
rect 10410 10656 10416 10668
rect 10371 10628 10416 10656
rect 10137 10619 10195 10625
rect 10410 10616 10416 10628
rect 10468 10616 10474 10668
rect 10502 10616 10508 10668
rect 10560 10656 10566 10668
rect 10704 10665 10732 10696
rect 10888 10665 10916 10764
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 11514 10792 11520 10804
rect 11475 10764 11520 10792
rect 11514 10752 11520 10764
rect 11572 10752 11578 10804
rect 11974 10792 11980 10804
rect 11935 10764 11980 10792
rect 11974 10752 11980 10764
rect 12032 10752 12038 10804
rect 11072 10724 11100 10752
rect 11885 10727 11943 10733
rect 11885 10724 11897 10727
rect 11072 10696 11897 10724
rect 11885 10693 11897 10696
rect 11931 10693 11943 10727
rect 12894 10724 12900 10736
rect 12855 10696 12900 10724
rect 11885 10687 11943 10693
rect 12894 10684 12900 10696
rect 12952 10684 12958 10736
rect 13354 10684 13360 10736
rect 13412 10724 13418 10736
rect 13541 10727 13599 10733
rect 13541 10724 13553 10727
rect 13412 10696 13553 10724
rect 13412 10684 13418 10696
rect 13541 10693 13553 10696
rect 13587 10693 13599 10727
rect 13541 10687 13599 10693
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 10560 10628 10609 10656
rect 10560 10616 10566 10628
rect 10597 10625 10609 10628
rect 10643 10625 10655 10659
rect 10597 10619 10655 10625
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 10873 10659 10931 10665
rect 10873 10625 10885 10659
rect 10919 10625 10931 10659
rect 12342 10656 12348 10668
rect 12303 10628 12348 10656
rect 10873 10619 10931 10625
rect 12342 10616 12348 10628
rect 12400 10616 12406 10668
rect 12802 10656 12808 10668
rect 12763 10628 12808 10656
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 12986 10656 12992 10668
rect 12947 10628 12992 10656
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 13262 10616 13268 10668
rect 13320 10656 13326 10668
rect 13449 10659 13507 10665
rect 13449 10656 13461 10659
rect 13320 10628 13461 10656
rect 13320 10616 13326 10628
rect 13449 10625 13461 10628
rect 13495 10625 13507 10659
rect 13449 10619 13507 10625
rect 7800 10560 8432 10588
rect 8496 10560 8984 10588
rect 9646 10560 9680 10600
rect 7800 10548 7806 10560
rect 7834 10520 7840 10532
rect 7668 10492 7840 10520
rect 7834 10480 7840 10492
rect 7892 10480 7898 10532
rect 8297 10523 8355 10529
rect 8297 10489 8309 10523
rect 8343 10520 8355 10523
rect 8496 10520 8524 10560
rect 8343 10492 8524 10520
rect 8956 10520 8984 10560
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 9858 10588 9864 10600
rect 9819 10560 9864 10588
rect 9858 10548 9864 10560
rect 9916 10548 9922 10600
rect 10321 10591 10379 10597
rect 10321 10557 10333 10591
rect 10367 10588 10379 10591
rect 10781 10591 10839 10597
rect 10781 10588 10793 10591
rect 10367 10560 10793 10588
rect 10367 10557 10379 10560
rect 10321 10551 10379 10557
rect 10781 10557 10793 10560
rect 10827 10557 10839 10591
rect 10781 10551 10839 10557
rect 12161 10591 12219 10597
rect 12161 10557 12173 10591
rect 12207 10588 12219 10591
rect 12618 10588 12624 10600
rect 12207 10560 12624 10588
rect 12207 10557 12219 10560
rect 12161 10551 12219 10557
rect 12618 10548 12624 10560
rect 12676 10588 12682 10600
rect 12894 10588 12900 10600
rect 12676 10560 12900 10588
rect 12676 10548 12682 10560
rect 12894 10548 12900 10560
rect 12952 10548 12958 10600
rect 11514 10520 11520 10532
rect 8956 10492 11520 10520
rect 8343 10489 8355 10492
rect 8297 10483 8355 10489
rect 11514 10480 11520 10492
rect 11572 10480 11578 10532
rect 5166 10412 5172 10464
rect 5224 10452 5230 10464
rect 5629 10455 5687 10461
rect 5629 10452 5641 10455
rect 5224 10424 5641 10452
rect 5224 10412 5230 10424
rect 5629 10421 5641 10424
rect 5675 10421 5687 10455
rect 5629 10415 5687 10421
rect 5810 10412 5816 10464
rect 5868 10452 5874 10464
rect 6178 10452 6184 10464
rect 5868 10424 6184 10452
rect 5868 10412 5874 10424
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 6822 10412 6828 10464
rect 6880 10452 6886 10464
rect 8478 10452 8484 10464
rect 6880 10424 8484 10452
rect 6880 10412 6886 10424
rect 8478 10412 8484 10424
rect 8536 10412 8542 10464
rect 9493 10455 9551 10461
rect 9493 10421 9505 10455
rect 9539 10452 9551 10455
rect 9674 10452 9680 10464
rect 9539 10424 9680 10452
rect 9539 10421 9551 10424
rect 9493 10415 9551 10421
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 9950 10452 9956 10464
rect 9911 10424 9956 10452
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10042 10412 10048 10464
rect 10100 10452 10106 10464
rect 10321 10455 10379 10461
rect 10321 10452 10333 10455
rect 10100 10424 10333 10452
rect 10100 10412 10106 10424
rect 10321 10421 10333 10424
rect 10367 10421 10379 10455
rect 10321 10415 10379 10421
rect 10686 10412 10692 10464
rect 10744 10452 10750 10464
rect 11146 10452 11152 10464
rect 10744 10424 11152 10452
rect 10744 10412 10750 10424
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 1104 10362 13892 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 12214 10362
rect 12266 10310 12278 10362
rect 12330 10310 12342 10362
rect 12394 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 13892 10362
rect 1104 10288 13892 10310
rect 3050 10248 3056 10260
rect 3011 10220 3056 10248
rect 3050 10208 3056 10220
rect 3108 10208 3114 10260
rect 5718 10248 5724 10260
rect 5679 10220 5724 10248
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 5994 10208 6000 10260
rect 6052 10248 6058 10260
rect 6914 10248 6920 10260
rect 6052 10220 6408 10248
rect 6875 10220 6920 10248
rect 6052 10208 6058 10220
rect 6270 10180 6276 10192
rect 5276 10152 6276 10180
rect 5276 10121 5304 10152
rect 6270 10140 6276 10152
rect 6328 10140 6334 10192
rect 6380 10180 6408 10220
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 7098 10208 7104 10260
rect 7156 10248 7162 10260
rect 7285 10251 7343 10257
rect 7285 10248 7297 10251
rect 7156 10220 7297 10248
rect 7156 10208 7162 10220
rect 7285 10217 7297 10220
rect 7331 10248 7343 10251
rect 7466 10248 7472 10260
rect 7331 10220 7472 10248
rect 7331 10217 7343 10220
rect 7285 10211 7343 10217
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 10321 10251 10379 10257
rect 10321 10217 10333 10251
rect 10367 10248 10379 10251
rect 10594 10248 10600 10260
rect 10367 10220 10600 10248
rect 10367 10217 10379 10220
rect 10321 10211 10379 10217
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 10873 10251 10931 10257
rect 10873 10217 10885 10251
rect 10919 10248 10931 10251
rect 10962 10248 10968 10260
rect 10919 10220 10968 10248
rect 10919 10217 10931 10220
rect 10873 10211 10931 10217
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 11146 10248 11152 10260
rect 11107 10220 11152 10248
rect 11146 10208 11152 10220
rect 11204 10208 11210 10260
rect 11422 10208 11428 10260
rect 11480 10248 11486 10260
rect 11517 10251 11575 10257
rect 11517 10248 11529 10251
rect 11480 10220 11529 10248
rect 11480 10208 11486 10220
rect 11517 10217 11529 10220
rect 11563 10217 11575 10251
rect 11517 10211 11575 10217
rect 12713 10251 12771 10257
rect 12713 10217 12725 10251
rect 12759 10248 12771 10251
rect 12986 10248 12992 10260
rect 12759 10220 12992 10248
rect 12759 10217 12771 10220
rect 12713 10211 12771 10217
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 7190 10180 7196 10192
rect 6380 10152 7196 10180
rect 7190 10140 7196 10152
rect 7248 10180 7254 10192
rect 8110 10180 8116 10192
rect 7248 10152 8116 10180
rect 7248 10140 7254 10152
rect 8110 10140 8116 10152
rect 8168 10180 8174 10192
rect 9309 10183 9367 10189
rect 9309 10180 9321 10183
rect 8168 10152 9321 10180
rect 8168 10140 8174 10152
rect 9309 10149 9321 10152
rect 9355 10180 9367 10183
rect 9950 10180 9956 10192
rect 9355 10152 9956 10180
rect 9355 10149 9367 10152
rect 9309 10143 9367 10149
rect 9950 10140 9956 10152
rect 10008 10180 10014 10192
rect 10686 10180 10692 10192
rect 10008 10152 10692 10180
rect 10008 10140 10014 10152
rect 10686 10140 10692 10152
rect 10744 10140 10750 10192
rect 10796 10152 11192 10180
rect 5261 10115 5319 10121
rect 5261 10081 5273 10115
rect 5307 10081 5319 10115
rect 5442 10112 5448 10124
rect 5403 10084 5448 10112
rect 5261 10075 5319 10081
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 6086 10112 6092 10124
rect 6047 10084 6092 10112
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 7006 10112 7012 10124
rect 6288 10084 7012 10112
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10044 3847 10047
rect 3878 10044 3884 10056
rect 3835 10016 3884 10044
rect 3835 10013 3847 10016
rect 3789 10007 3847 10013
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 5166 10044 5172 10056
rect 5127 10016 5172 10044
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 5902 10004 5908 10056
rect 5960 10044 5966 10056
rect 5997 10047 6055 10053
rect 5997 10044 6009 10047
rect 5960 10016 6009 10044
rect 5960 10004 5966 10016
rect 5997 10013 6009 10016
rect 6043 10013 6055 10047
rect 6178 10044 6184 10056
rect 6139 10016 6184 10044
rect 5997 10007 6055 10013
rect 2958 9976 2964 9988
rect 2919 9948 2964 9976
rect 2958 9936 2964 9948
rect 3016 9936 3022 9988
rect 6012 9976 6040 10007
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 6288 10053 6316 10084
rect 7006 10072 7012 10084
rect 7064 10112 7070 10124
rect 7469 10115 7527 10121
rect 7469 10112 7481 10115
rect 7064 10084 7481 10112
rect 7064 10072 7070 10084
rect 7469 10081 7481 10084
rect 7515 10081 7527 10115
rect 8573 10115 8631 10121
rect 8573 10112 8585 10115
rect 7469 10075 7527 10081
rect 8036 10084 8585 10112
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10013 6331 10047
rect 6273 10007 6331 10013
rect 6457 10047 6515 10053
rect 6457 10013 6469 10047
rect 6503 10044 6515 10047
rect 7098 10044 7104 10056
rect 6503 10016 7104 10044
rect 6503 10013 6515 10016
rect 6457 10007 6515 10013
rect 7098 10004 7104 10016
rect 7156 10004 7162 10056
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10013 7251 10047
rect 7193 10007 7251 10013
rect 7377 10047 7435 10053
rect 7377 10013 7389 10047
rect 7423 10013 7435 10047
rect 7558 10044 7564 10056
rect 7519 10016 7564 10044
rect 7377 10007 7435 10013
rect 6730 9976 6736 9988
rect 6012 9948 6736 9976
rect 6730 9936 6736 9948
rect 6788 9976 6794 9988
rect 7208 9976 7236 10007
rect 6788 9948 7236 9976
rect 7392 9976 7420 10007
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 7834 10004 7840 10056
rect 7892 10044 7898 10056
rect 8036 10044 8064 10084
rect 8573 10081 8585 10084
rect 8619 10081 8631 10115
rect 8573 10075 8631 10081
rect 9401 10115 9459 10121
rect 9401 10081 9413 10115
rect 9447 10112 9459 10115
rect 10137 10115 10195 10121
rect 10137 10112 10149 10115
rect 9447 10084 10149 10112
rect 9447 10081 9459 10084
rect 9401 10075 9459 10081
rect 10137 10081 10149 10084
rect 10183 10081 10195 10115
rect 10137 10075 10195 10081
rect 7892 10016 8064 10044
rect 8389 10047 8447 10053
rect 7892 10004 7898 10016
rect 8389 10013 8401 10047
rect 8435 10044 8447 10047
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8435 10016 8953 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 7650 9976 7656 9988
rect 7392 9948 7656 9976
rect 6788 9936 6794 9948
rect 7650 9936 7656 9948
rect 7708 9936 7714 9988
rect 8481 9979 8539 9985
rect 8481 9945 8493 9979
rect 8527 9976 8539 9979
rect 8662 9976 8668 9988
rect 8527 9948 8668 9976
rect 8527 9945 8539 9948
rect 8481 9939 8539 9945
rect 8662 9936 8668 9948
rect 8720 9936 8726 9988
rect 8846 9936 8852 9988
rect 8904 9976 8910 9988
rect 9232 9976 9260 10007
rect 9490 10004 9496 10056
rect 9548 10044 9554 10056
rect 9548 10016 9593 10044
rect 9548 10004 9554 10016
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 10502 10044 10508 10056
rect 9732 10016 10508 10044
rect 9732 10004 9738 10016
rect 10502 10004 10508 10016
rect 10560 10044 10566 10056
rect 10796 10053 10824 10152
rect 11164 10053 11192 10152
rect 12894 10072 12900 10124
rect 12952 10112 12958 10124
rect 13265 10115 13323 10121
rect 13265 10112 13277 10115
rect 12952 10084 13277 10112
rect 12952 10072 12958 10084
rect 13265 10081 13277 10084
rect 13311 10081 13323 10115
rect 13265 10075 13323 10081
rect 10597 10047 10655 10053
rect 10597 10044 10609 10047
rect 10560 10016 10609 10044
rect 10560 10004 10566 10016
rect 10597 10013 10609 10016
rect 10643 10013 10655 10047
rect 10781 10047 10839 10053
rect 10781 10022 10793 10047
rect 10597 10007 10655 10013
rect 10704 10013 10793 10022
rect 10827 10013 10839 10047
rect 10965 10047 11023 10053
rect 10965 10038 10977 10047
rect 10704 10007 10839 10013
rect 10888 10013 10977 10038
rect 11011 10013 11023 10047
rect 10888 10010 11023 10013
rect 10704 9994 10824 10007
rect 9858 9976 9864 9988
rect 8904 9948 9864 9976
rect 8904 9936 8910 9948
rect 9858 9936 9864 9948
rect 9916 9976 9922 9988
rect 10704 9976 10732 9994
rect 9916 9948 10732 9976
rect 9916 9936 9922 9948
rect 3234 9868 3240 9920
rect 3292 9908 3298 9920
rect 3881 9911 3939 9917
rect 3881 9908 3893 9911
rect 3292 9880 3893 9908
rect 3292 9868 3298 9880
rect 3881 9877 3893 9880
rect 3927 9877 3939 9911
rect 3881 9871 3939 9877
rect 4801 9911 4859 9917
rect 4801 9877 4813 9911
rect 4847 9908 4859 9911
rect 4890 9908 4896 9920
rect 4847 9880 4896 9908
rect 4847 9877 4859 9880
rect 4801 9871 4859 9877
rect 4890 9868 4896 9880
rect 4948 9868 4954 9920
rect 8018 9908 8024 9920
rect 7979 9880 8024 9908
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 10137 9911 10195 9917
rect 10137 9877 10149 9911
rect 10183 9908 10195 9911
rect 10888 9908 10916 10010
rect 10965 10007 11023 10010
rect 11149 10047 11207 10053
rect 11149 10013 11161 10047
rect 11195 10013 11207 10047
rect 11149 10007 11207 10013
rect 11333 10047 11391 10053
rect 11333 10013 11345 10047
rect 11379 10044 11391 10047
rect 12437 10047 12495 10053
rect 11379 10016 11468 10044
rect 11379 10013 11391 10016
rect 11333 10007 11391 10013
rect 11238 9936 11244 9988
rect 11296 9976 11302 9988
rect 11440 9976 11468 10016
rect 12437 10013 12449 10047
rect 12483 10044 12495 10047
rect 12802 10044 12808 10056
rect 12483 10016 12808 10044
rect 12483 10013 12495 10016
rect 12437 10007 12495 10013
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 13078 9976 13084 9988
rect 11296 9948 11468 9976
rect 13039 9948 13084 9976
rect 11296 9936 11302 9948
rect 13078 9936 13084 9948
rect 13136 9936 13142 9988
rect 11330 9908 11336 9920
rect 10183 9880 11336 9908
rect 10183 9877 10195 9880
rect 10137 9871 10195 9877
rect 11330 9868 11336 9880
rect 11388 9868 11394 9920
rect 12526 9908 12532 9920
rect 12487 9880 12532 9908
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 13170 9868 13176 9920
rect 13228 9908 13234 9920
rect 13228 9880 13273 9908
rect 13228 9868 13234 9880
rect 1104 9818 13892 9840
rect 1104 9766 8214 9818
rect 8266 9766 8278 9818
rect 8330 9766 8342 9818
rect 8394 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 13892 9818
rect 1104 9744 13892 9766
rect 1486 9664 1492 9716
rect 1544 9704 1550 9716
rect 1544 9676 4752 9704
rect 1544 9664 1550 9676
rect 3326 9636 3332 9648
rect 3160 9608 3332 9636
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9568 1731 9571
rect 2222 9568 2228 9580
rect 1719 9540 2228 9568
rect 1719 9537 1731 9540
rect 1673 9531 1731 9537
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 3160 9577 3188 9608
rect 3326 9596 3332 9608
rect 3384 9636 3390 9648
rect 3421 9639 3479 9645
rect 3421 9636 3433 9639
rect 3384 9608 3433 9636
rect 3384 9596 3390 9608
rect 3421 9605 3433 9608
rect 3467 9636 3479 9639
rect 3467 9608 4660 9636
rect 3467 9605 3479 9608
rect 3421 9599 3479 9605
rect 3145 9571 3203 9577
rect 3145 9537 3157 9571
rect 3191 9537 3203 9571
rect 3145 9531 3203 9537
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9568 3755 9571
rect 3878 9568 3884 9580
rect 3743 9540 3884 9568
rect 3743 9537 3755 9540
rect 3697 9531 3755 9537
rect 3878 9528 3884 9540
rect 3936 9528 3942 9580
rect 4632 9577 4660 9608
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9568 4399 9571
rect 4617 9571 4675 9577
rect 4387 9540 4568 9568
rect 4387 9537 4399 9540
rect 4341 9531 4399 9537
rect 2958 9432 2964 9444
rect 2919 9404 2964 9432
rect 2958 9392 2964 9404
rect 3016 9392 3022 9444
rect 4540 9432 4568 9540
rect 4617 9537 4629 9571
rect 4663 9537 4675 9571
rect 4617 9531 4675 9537
rect 4724 9500 4752 9676
rect 6178 9664 6184 9716
rect 6236 9704 6242 9716
rect 6914 9704 6920 9716
rect 6236 9676 6920 9704
rect 6236 9664 6242 9676
rect 6914 9664 6920 9676
rect 6972 9704 6978 9716
rect 7650 9704 7656 9716
rect 6972 9676 7656 9704
rect 6972 9664 6978 9676
rect 7650 9664 7656 9676
rect 7708 9704 7714 9716
rect 8757 9707 8815 9713
rect 7708 9676 7788 9704
rect 7708 9664 7714 9676
rect 5074 9636 5080 9648
rect 5035 9608 5080 9636
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 7760 9636 7788 9676
rect 8757 9673 8769 9707
rect 8803 9704 8815 9707
rect 9490 9704 9496 9716
rect 8803 9676 9496 9704
rect 8803 9673 8815 9676
rect 8757 9667 8815 9673
rect 9490 9664 9496 9676
rect 9548 9664 9554 9716
rect 10410 9664 10416 9716
rect 10468 9704 10474 9716
rect 10468 9676 10824 9704
rect 10468 9664 10474 9676
rect 7837 9639 7895 9645
rect 7837 9636 7849 9639
rect 7760 9608 7849 9636
rect 7837 9605 7849 9608
rect 7883 9605 7895 9639
rect 7837 9599 7895 9605
rect 8021 9639 8079 9645
rect 8021 9605 8033 9639
rect 8067 9636 8079 9639
rect 8202 9636 8208 9648
rect 8067 9608 8208 9636
rect 8067 9605 8079 9608
rect 8021 9599 8079 9605
rect 8202 9596 8208 9608
rect 8260 9596 8266 9648
rect 8297 9639 8355 9645
rect 8297 9605 8309 9639
rect 8343 9636 8355 9639
rect 8846 9636 8852 9648
rect 8343 9608 8852 9636
rect 8343 9605 8355 9608
rect 8297 9599 8355 9605
rect 8846 9596 8852 9608
rect 8904 9596 8910 9648
rect 9030 9636 9036 9648
rect 8991 9608 9036 9636
rect 9030 9596 9036 9608
rect 9088 9596 9094 9648
rect 9122 9596 9128 9648
rect 9180 9636 9186 9648
rect 10796 9645 10824 9676
rect 10597 9639 10655 9645
rect 10597 9636 10609 9639
rect 9180 9608 10609 9636
rect 9180 9596 9186 9608
rect 10597 9605 10609 9608
rect 10643 9605 10655 9639
rect 10597 9599 10655 9605
rect 10781 9639 10839 9645
rect 10781 9605 10793 9639
rect 10827 9636 10839 9639
rect 10965 9639 11023 9645
rect 10827 9608 10861 9636
rect 10827 9605 10839 9608
rect 10781 9599 10839 9605
rect 10965 9605 10977 9639
rect 11011 9636 11023 9639
rect 11054 9636 11060 9648
rect 11011 9608 11060 9636
rect 11011 9605 11023 9608
rect 10965 9599 11023 9605
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 6457 9571 6515 9577
rect 6457 9568 6469 9571
rect 5215 9540 6469 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 6457 9537 6469 9540
rect 6503 9537 6515 9571
rect 6730 9568 6736 9580
rect 6691 9540 6736 9568
rect 6457 9531 6515 9537
rect 6730 9528 6736 9540
rect 6788 9528 6794 9580
rect 6822 9528 6828 9580
rect 6880 9568 6886 9580
rect 7190 9568 7196 9580
rect 6880 9540 6925 9568
rect 7151 9540 7196 9568
rect 6880 9528 6886 9540
rect 7190 9528 7196 9540
rect 7248 9568 7254 9580
rect 7558 9568 7564 9580
rect 7248 9540 7564 9568
rect 7248 9528 7254 9540
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 8478 9568 8484 9580
rect 8439 9540 8484 9568
rect 8478 9528 8484 9540
rect 8536 9528 8542 9580
rect 8589 9571 8647 9577
rect 8589 9537 8601 9571
rect 8635 9568 8647 9571
rect 9217 9571 9275 9577
rect 8635 9540 8708 9568
rect 8635 9537 8647 9540
rect 8589 9531 8647 9537
rect 4985 9503 5043 9509
rect 4985 9500 4997 9503
rect 4724 9472 4997 9500
rect 4985 9469 4997 9472
rect 5031 9500 5043 9503
rect 5442 9500 5448 9512
rect 5031 9472 5448 9500
rect 5031 9469 5043 9472
rect 4985 9463 5043 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 6181 9503 6239 9509
rect 6181 9469 6193 9503
rect 6227 9500 6239 9503
rect 8680 9500 8708 9540
rect 9217 9537 9229 9571
rect 9263 9537 9275 9571
rect 9217 9531 9275 9537
rect 8754 9500 8760 9512
rect 6227 9472 8340 9500
rect 8680 9472 8760 9500
rect 6227 9469 6239 9472
rect 6181 9463 6239 9469
rect 4614 9432 4620 9444
rect 4527 9404 4620 9432
rect 4614 9392 4620 9404
rect 4672 9432 4678 9444
rect 8018 9432 8024 9444
rect 4672 9404 8024 9432
rect 4672 9392 4678 9404
rect 8018 9392 8024 9404
rect 8076 9392 8082 9444
rect 8312 9432 8340 9472
rect 8754 9460 8760 9472
rect 8812 9500 8818 9512
rect 9232 9500 9260 9531
rect 9306 9528 9312 9580
rect 9364 9568 9370 9580
rect 9493 9571 9551 9577
rect 9364 9540 9409 9568
rect 9364 9528 9370 9540
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 8812 9472 9260 9500
rect 9508 9500 9536 9531
rect 10226 9528 10232 9580
rect 10284 9568 10290 9580
rect 10413 9571 10471 9577
rect 10413 9568 10425 9571
rect 10284 9540 10425 9568
rect 10284 9528 10290 9540
rect 10413 9537 10425 9540
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 10502 9500 10508 9512
rect 9508 9472 10508 9500
rect 8812 9460 8818 9472
rect 10502 9460 10508 9472
rect 10560 9460 10566 9512
rect 10612 9500 10640 9599
rect 11054 9596 11060 9608
rect 11112 9636 11118 9648
rect 11422 9636 11428 9648
rect 11112 9608 11428 9636
rect 11112 9596 11118 9608
rect 11422 9596 11428 9608
rect 11480 9596 11486 9648
rect 10870 9568 10876 9580
rect 10783 9540 10876 9568
rect 10870 9528 10876 9540
rect 10928 9568 10934 9580
rect 11514 9568 11520 9580
rect 10928 9540 11284 9568
rect 11475 9540 11520 9568
rect 10928 9528 10934 9540
rect 11146 9500 11152 9512
rect 10612 9472 11152 9500
rect 11146 9460 11152 9472
rect 11204 9460 11210 9512
rect 11256 9500 11284 9540
rect 11514 9528 11520 9540
rect 11572 9528 11578 9580
rect 12526 9568 12532 9580
rect 12487 9540 12532 9568
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 13354 9568 13360 9580
rect 13315 9540 13360 9568
rect 13354 9528 13360 9540
rect 13412 9528 13418 9580
rect 11606 9500 11612 9512
rect 11256 9472 11612 9500
rect 11606 9460 11612 9472
rect 11664 9460 11670 9512
rect 9401 9435 9459 9441
rect 8312 9404 9351 9432
rect 3786 9324 3792 9376
rect 3844 9364 3850 9376
rect 4433 9367 4491 9373
rect 4433 9364 4445 9367
rect 3844 9336 4445 9364
rect 3844 9324 3850 9336
rect 4433 9333 4445 9336
rect 4479 9333 4491 9367
rect 4433 9327 4491 9333
rect 5537 9367 5595 9373
rect 5537 9333 5549 9367
rect 5583 9364 5595 9367
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 5583 9336 6193 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 6181 9333 6193 9336
rect 6227 9333 6239 9367
rect 6914 9364 6920 9376
rect 6875 9336 6920 9364
rect 6181 9327 6239 9333
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 7742 9364 7748 9376
rect 7064 9336 7109 9364
rect 7703 9336 7748 9364
rect 7064 9324 7070 9336
rect 7742 9324 7748 9336
rect 7800 9324 7806 9376
rect 7926 9324 7932 9376
rect 7984 9364 7990 9376
rect 8297 9367 8355 9373
rect 8297 9364 8309 9367
rect 7984 9336 8309 9364
rect 7984 9324 7990 9336
rect 8297 9333 8309 9336
rect 8343 9364 8355 9367
rect 9214 9364 9220 9376
rect 8343 9336 9220 9364
rect 8343 9333 8355 9336
rect 8297 9327 8355 9333
rect 9214 9324 9220 9336
rect 9272 9324 9278 9376
rect 9323 9364 9351 9404
rect 9401 9401 9413 9435
rect 9447 9432 9459 9435
rect 9674 9432 9680 9444
rect 9447 9404 9680 9432
rect 9447 9401 9459 9404
rect 9401 9395 9459 9401
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 10134 9392 10140 9444
rect 10192 9432 10198 9444
rect 10778 9432 10784 9444
rect 10192 9404 10784 9432
rect 10192 9392 10198 9404
rect 10778 9392 10784 9404
rect 10836 9392 10842 9444
rect 12802 9432 12808 9444
rect 12763 9404 12808 9432
rect 12802 9392 12808 9404
rect 12860 9392 12866 9444
rect 11330 9364 11336 9376
rect 9323 9336 11336 9364
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 13262 9364 13268 9376
rect 13223 9336 13268 9364
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 1104 9274 13892 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 12214 9274
rect 12266 9222 12278 9274
rect 12330 9222 12342 9274
rect 12394 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 13892 9274
rect 1104 9200 13892 9222
rect 2222 9160 2228 9172
rect 2183 9132 2228 9160
rect 2222 9120 2228 9132
rect 2280 9120 2286 9172
rect 6273 9163 6331 9169
rect 6273 9160 6285 9163
rect 2746 9132 6285 9160
rect 1486 8984 1492 9036
rect 1544 9024 1550 9036
rect 1581 9027 1639 9033
rect 1581 9024 1593 9027
rect 1544 8996 1593 9024
rect 1544 8984 1550 8996
rect 1581 8993 1593 8996
rect 1627 8993 1639 9027
rect 1762 9024 1768 9036
rect 1723 8996 1768 9024
rect 1581 8987 1639 8993
rect 1762 8984 1768 8996
rect 1820 8984 1826 9036
rect 2240 9024 2268 9120
rect 2409 9027 2467 9033
rect 2409 9024 2421 9027
rect 2240 8996 2421 9024
rect 2409 8993 2421 8996
rect 2455 8993 2467 9027
rect 2409 8987 2467 8993
rect 1857 8959 1915 8965
rect 1857 8925 1869 8959
rect 1903 8956 1915 8959
rect 2746 8956 2774 9132
rect 6273 9129 6285 9132
rect 6319 9129 6331 9163
rect 6273 9123 6331 9129
rect 8021 9163 8079 9169
rect 8021 9129 8033 9163
rect 8067 9160 8079 9163
rect 8110 9160 8116 9172
rect 8067 9132 8116 9160
rect 8067 9129 8079 9132
rect 8021 9123 8079 9129
rect 8110 9120 8116 9132
rect 8168 9120 8174 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8938 9160 8944 9172
rect 8352 9132 8944 9160
rect 8352 9120 8358 9132
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 9122 9160 9128 9172
rect 9083 9132 9128 9160
rect 9122 9120 9128 9132
rect 9180 9120 9186 9172
rect 9493 9163 9551 9169
rect 9493 9129 9505 9163
rect 9539 9160 9551 9163
rect 10134 9160 10140 9172
rect 9539 9132 10140 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 10226 9120 10232 9172
rect 10284 9160 10290 9172
rect 10689 9163 10747 9169
rect 10689 9160 10701 9163
rect 10284 9132 10701 9160
rect 10284 9120 10290 9132
rect 10689 9129 10701 9132
rect 10735 9129 10747 9163
rect 10689 9123 10747 9129
rect 11146 9120 11152 9172
rect 11204 9160 11210 9172
rect 11241 9163 11299 9169
rect 11241 9160 11253 9163
rect 11204 9132 11253 9160
rect 11204 9120 11210 9132
rect 11241 9129 11253 9132
rect 11287 9129 11299 9163
rect 11241 9123 11299 9129
rect 2869 9095 2927 9101
rect 2869 9061 2881 9095
rect 2915 9092 2927 9095
rect 2958 9092 2964 9104
rect 2915 9064 2964 9092
rect 2915 9061 2927 9064
rect 2869 9055 2927 9061
rect 2958 9052 2964 9064
rect 3016 9052 3022 9104
rect 3326 9092 3332 9104
rect 3287 9064 3332 9092
rect 3326 9052 3332 9064
rect 3384 9052 3390 9104
rect 3878 9092 3884 9104
rect 3839 9064 3884 9092
rect 3878 9052 3884 9064
rect 3936 9052 3942 9104
rect 6641 9095 6699 9101
rect 6641 9061 6653 9095
rect 6687 9092 6699 9095
rect 6914 9092 6920 9104
rect 6687 9064 6920 9092
rect 6687 9061 6699 9064
rect 6641 9055 6699 9061
rect 6914 9052 6920 9064
rect 6972 9052 6978 9104
rect 7282 9092 7288 9104
rect 7243 9064 7288 9092
rect 7282 9052 7288 9064
rect 7340 9052 7346 9104
rect 7558 9052 7564 9104
rect 7616 9092 7622 9104
rect 9674 9092 9680 9104
rect 7616 9064 9680 9092
rect 7616 9052 7622 9064
rect 9674 9052 9680 9064
rect 9732 9052 9738 9104
rect 9766 9052 9772 9104
rect 9824 9092 9830 9104
rect 10318 9092 10324 9104
rect 9824 9064 10324 9092
rect 9824 9052 9830 9064
rect 10318 9052 10324 9064
rect 10376 9052 10382 9104
rect 12437 9095 12495 9101
rect 12437 9061 12449 9095
rect 12483 9092 12495 9095
rect 12802 9092 12808 9104
rect 12483 9064 12808 9092
rect 12483 9061 12495 9064
rect 12437 9055 12495 9061
rect 3786 9024 3792 9036
rect 3747 8996 3792 9024
rect 3786 8984 3792 8996
rect 3844 8984 3850 9036
rect 4341 9027 4399 9033
rect 4341 8993 4353 9027
rect 4387 9024 4399 9027
rect 4614 9024 4620 9036
rect 4387 8996 4620 9024
rect 4387 8993 4399 8996
rect 4341 8987 4399 8993
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 7190 9024 7196 9036
rect 6472 8996 7196 9024
rect 1903 8928 2774 8956
rect 2961 8959 3019 8965
rect 1903 8925 1915 8928
rect 1857 8919 1915 8925
rect 2961 8925 2973 8959
rect 3007 8956 3019 8959
rect 3234 8956 3240 8968
rect 3007 8928 3240 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 3602 8956 3608 8968
rect 3515 8928 3608 8956
rect 3602 8916 3608 8928
rect 3660 8956 3666 8968
rect 6472 8965 6500 8996
rect 7190 8984 7196 8996
rect 7248 9024 7254 9036
rect 8754 9024 8760 9036
rect 7248 8996 8760 9024
rect 7248 8984 7254 8996
rect 8754 8984 8760 8996
rect 8812 9024 8818 9036
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 8812 8996 9229 9024
rect 8812 8984 8818 8996
rect 9217 8993 9229 8996
rect 9263 8993 9275 9027
rect 9217 8987 9275 8993
rect 10042 8984 10048 9036
rect 10100 9024 10106 9036
rect 10778 9024 10784 9036
rect 10100 8996 10784 9024
rect 10100 8984 10106 8996
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 12452 9024 12480 9055
rect 12802 9052 12808 9064
rect 12860 9052 12866 9104
rect 11716 8996 12480 9024
rect 12529 9027 12587 9033
rect 4433 8959 4491 8965
rect 4433 8956 4445 8959
rect 3660 8928 4445 8956
rect 3660 8916 3666 8928
rect 4433 8925 4445 8928
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8925 6515 8959
rect 6457 8919 6515 8925
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8925 6607 8959
rect 6730 8956 6736 8968
rect 6691 8928 6736 8956
rect 6549 8919 6607 8925
rect 3142 8888 3148 8900
rect 3103 8860 3148 8888
rect 3142 8848 3148 8860
rect 3200 8848 3206 8900
rect 4617 8891 4675 8897
rect 4617 8857 4629 8891
rect 4663 8888 4675 8891
rect 5350 8888 5356 8900
rect 4663 8860 5356 8888
rect 4663 8857 4675 8860
rect 4617 8851 4675 8857
rect 5350 8848 5356 8860
rect 5408 8848 5414 8900
rect 6564 8888 6592 8919
rect 6730 8916 6736 8928
rect 6788 8916 6794 8968
rect 7466 8956 7472 8968
rect 7427 8928 7472 8956
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9125 8919 9183 8925
rect 9692 8928 10149 8956
rect 7006 8888 7012 8900
rect 6564 8860 7012 8888
rect 7006 8848 7012 8860
rect 7064 8888 7070 8900
rect 7064 8860 7236 8888
rect 7064 8848 7070 8860
rect 7208 8832 7236 8860
rect 7742 8848 7748 8900
rect 7800 8888 7806 8900
rect 7837 8891 7895 8897
rect 7837 8888 7849 8891
rect 7800 8860 7849 8888
rect 7800 8848 7806 8860
rect 7837 8857 7849 8860
rect 7883 8857 7895 8891
rect 7837 8851 7895 8857
rect 8018 8848 8024 8900
rect 8076 8888 8082 8900
rect 8113 8891 8171 8897
rect 8113 8888 8125 8891
rect 8076 8860 8125 8888
rect 8076 8848 8082 8860
rect 8113 8857 8125 8860
rect 8159 8857 8171 8891
rect 8113 8851 8171 8857
rect 8297 8891 8355 8897
rect 8297 8857 8309 8891
rect 8343 8888 8355 8891
rect 9030 8888 9036 8900
rect 8343 8860 9036 8888
rect 8343 8857 8355 8860
rect 8297 8851 8355 8857
rect 9030 8848 9036 8860
rect 9088 8848 9094 8900
rect 9140 8888 9168 8919
rect 9692 8897 9720 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 11054 8956 11060 8968
rect 10137 8919 10195 8925
rect 10244 8928 11060 8956
rect 9677 8891 9735 8897
rect 9677 8888 9689 8891
rect 9140 8860 9689 8888
rect 9677 8857 9689 8860
rect 9723 8857 9735 8891
rect 9677 8851 9735 8857
rect 9861 8891 9919 8897
rect 9861 8857 9873 8891
rect 9907 8857 9919 8891
rect 10042 8888 10048 8900
rect 10003 8860 10048 8888
rect 9861 8851 9919 8857
rect 3418 8820 3424 8832
rect 3379 8792 3424 8820
rect 3418 8780 3424 8792
rect 3476 8780 3482 8832
rect 4798 8820 4804 8832
rect 4759 8792 4804 8820
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 7190 8780 7196 8832
rect 7248 8820 7254 8832
rect 7466 8820 7472 8832
rect 7248 8792 7472 8820
rect 7248 8780 7254 8792
rect 7466 8780 7472 8792
rect 7524 8820 7530 8832
rect 7561 8823 7619 8829
rect 7561 8820 7573 8823
rect 7524 8792 7573 8820
rect 7524 8780 7530 8792
rect 7561 8789 7573 8792
rect 7607 8789 7619 8823
rect 7561 8783 7619 8789
rect 7653 8823 7711 8829
rect 7653 8789 7665 8823
rect 7699 8820 7711 8823
rect 8036 8820 8064 8848
rect 7699 8792 8064 8820
rect 9876 8820 9904 8851
rect 10042 8848 10048 8860
rect 10100 8848 10106 8900
rect 10244 8888 10272 8928
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8956 11207 8959
rect 11606 8956 11612 8968
rect 11195 8928 11612 8956
rect 11195 8925 11207 8928
rect 11149 8919 11207 8925
rect 11606 8916 11612 8928
rect 11664 8916 11670 8968
rect 11716 8965 11744 8996
rect 12529 8993 12541 9027
rect 12575 9024 12587 9027
rect 13262 9024 13268 9036
rect 12575 8996 13268 9024
rect 12575 8993 12587 8996
rect 12529 8987 12587 8993
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 11701 8959 11759 8965
rect 11701 8925 11713 8959
rect 11747 8925 11759 8959
rect 11701 8919 11759 8925
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8925 12035 8959
rect 12618 8956 12624 8968
rect 12579 8928 12624 8956
rect 11977 8919 12035 8925
rect 10686 8888 10692 8900
rect 10152 8860 10272 8888
rect 10647 8860 10692 8888
rect 10152 8820 10180 8860
rect 10686 8848 10692 8860
rect 10744 8848 10750 8900
rect 10870 8888 10876 8900
rect 10831 8860 10876 8888
rect 10870 8848 10876 8860
rect 10928 8848 10934 8900
rect 10962 8848 10968 8900
rect 11020 8888 11026 8900
rect 11020 8860 11065 8888
rect 11020 8848 11026 8860
rect 11514 8848 11520 8900
rect 11572 8888 11578 8900
rect 11992 8888 12020 8919
rect 12618 8916 12624 8928
rect 12676 8916 12682 8968
rect 13354 8956 13360 8968
rect 13315 8928 13360 8956
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 11572 8860 12020 8888
rect 11572 8848 11578 8860
rect 12710 8848 12716 8900
rect 12768 8888 12774 8900
rect 13541 8891 13599 8897
rect 13541 8888 13553 8891
rect 12768 8860 13553 8888
rect 12768 8848 12774 8860
rect 13541 8857 13553 8860
rect 13587 8857 13599 8891
rect 13541 8851 13599 8857
rect 9876 8792 10180 8820
rect 10229 8823 10287 8829
rect 7699 8789 7711 8792
rect 7653 8783 7711 8789
rect 10229 8789 10241 8823
rect 10275 8820 10287 8823
rect 10318 8820 10324 8832
rect 10275 8792 10324 8820
rect 10275 8789 10287 8792
rect 10229 8783 10287 8789
rect 10318 8780 10324 8792
rect 10376 8780 10382 8832
rect 10502 8820 10508 8832
rect 10463 8792 10508 8820
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 10594 8780 10600 8832
rect 10652 8820 10658 8832
rect 10888 8820 10916 8848
rect 11790 8820 11796 8832
rect 10652 8792 10916 8820
rect 11751 8792 11796 8820
rect 10652 8780 10658 8792
rect 11790 8780 11796 8792
rect 11848 8780 11854 8832
rect 1104 8730 13892 8752
rect 1104 8678 8214 8730
rect 8266 8678 8278 8730
rect 8330 8678 8342 8730
rect 8394 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 13892 8730
rect 1104 8656 13892 8678
rect 6825 8619 6883 8625
rect 6825 8616 6837 8619
rect 4172 8588 6837 8616
rect 3142 8548 3148 8560
rect 3103 8520 3148 8548
rect 3142 8508 3148 8520
rect 3200 8508 3206 8560
rect 3237 8551 3295 8557
rect 3237 8517 3249 8551
rect 3283 8548 3295 8551
rect 3602 8548 3608 8560
rect 3283 8520 3608 8548
rect 3283 8517 3295 8520
rect 3237 8511 3295 8517
rect 1578 8480 1584 8492
rect 1539 8452 1584 8480
rect 1578 8440 1584 8452
rect 1636 8440 1642 8492
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3252 8480 3280 8511
rect 3602 8508 3608 8520
rect 3660 8508 3666 8560
rect 4172 8492 4200 8588
rect 6825 8585 6837 8588
rect 6871 8585 6883 8619
rect 6825 8579 6883 8585
rect 7285 8619 7343 8625
rect 7285 8585 7297 8619
rect 7331 8616 7343 8619
rect 7374 8616 7380 8628
rect 7331 8588 7380 8616
rect 7331 8585 7343 8588
rect 7285 8579 7343 8585
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 7466 8576 7472 8628
rect 7524 8616 7530 8628
rect 7926 8616 7932 8628
rect 7524 8588 7932 8616
rect 7524 8576 7530 8588
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 8018 8576 8024 8628
rect 8076 8616 8082 8628
rect 8849 8619 8907 8625
rect 8076 8588 8524 8616
rect 8076 8576 8082 8588
rect 5920 8520 7144 8548
rect 3099 8452 3280 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 3421 8483 3479 8489
rect 3421 8480 3433 8483
rect 3384 8452 3433 8480
rect 3384 8440 3390 8452
rect 3421 8449 3433 8452
rect 3467 8449 3479 8483
rect 4154 8480 4160 8492
rect 4067 8452 4160 8480
rect 3421 8443 3479 8449
rect 4154 8440 4160 8452
rect 4212 8440 4218 8492
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 4614 8480 4620 8492
rect 4479 8452 4620 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 5718 8440 5724 8492
rect 5776 8480 5782 8492
rect 5920 8489 5948 8520
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5776 8452 5917 8480
rect 5776 8440 5782 8452
rect 5905 8449 5917 8452
rect 5951 8449 5963 8483
rect 6546 8480 6552 8492
rect 6507 8452 6552 8480
rect 5905 8443 5963 8449
rect 6546 8440 6552 8452
rect 6604 8440 6610 8492
rect 5350 8304 5356 8356
rect 5408 8344 5414 8356
rect 5721 8347 5779 8353
rect 5721 8344 5733 8347
rect 5408 8316 5733 8344
rect 5408 8304 5414 8316
rect 5721 8313 5733 8316
rect 5767 8313 5779 8347
rect 7116 8344 7144 8520
rect 7742 8508 7748 8560
rect 7800 8548 7806 8560
rect 8202 8548 8208 8560
rect 7800 8520 8208 8548
rect 7800 8508 7806 8520
rect 8202 8508 8208 8520
rect 8260 8508 8266 8560
rect 8496 8557 8524 8588
rect 8849 8585 8861 8619
rect 8895 8616 8907 8619
rect 9122 8616 9128 8628
rect 8895 8588 9128 8616
rect 8895 8585 8907 8588
rect 8849 8579 8907 8585
rect 9122 8576 9128 8588
rect 9180 8576 9186 8628
rect 10226 8616 10232 8628
rect 9692 8588 10232 8616
rect 8481 8551 8539 8557
rect 8481 8517 8493 8551
rect 8527 8517 8539 8551
rect 8481 8511 8539 8517
rect 8665 8551 8723 8557
rect 8665 8517 8677 8551
rect 8711 8548 8723 8551
rect 8938 8548 8944 8560
rect 8711 8520 8944 8548
rect 8711 8517 8723 8520
rect 8665 8511 8723 8517
rect 8938 8508 8944 8520
rect 8996 8548 9002 8560
rect 9692 8548 9720 8588
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 8996 8520 9720 8548
rect 8996 8508 9002 8520
rect 7193 8483 7251 8489
rect 7193 8449 7205 8483
rect 7239 8480 7251 8483
rect 7653 8483 7711 8489
rect 7653 8480 7665 8483
rect 7239 8452 7665 8480
rect 7239 8449 7251 8452
rect 7193 8443 7251 8449
rect 7653 8449 7665 8452
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 7466 8412 7472 8424
rect 7427 8384 7472 8412
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 7558 8372 7564 8424
rect 7616 8412 7622 8424
rect 7852 8412 7880 8443
rect 7926 8440 7932 8492
rect 7984 8480 7990 8492
rect 8297 8483 8355 8489
rect 8297 8480 8309 8483
rect 7984 8452 8309 8480
rect 7984 8440 7990 8452
rect 8297 8449 8309 8452
rect 8343 8480 8355 8483
rect 8757 8483 8815 8489
rect 8757 8480 8769 8483
rect 8343 8452 8769 8480
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 8757 8449 8769 8452
rect 8803 8449 8815 8483
rect 9490 8480 9496 8492
rect 9451 8452 9496 8480
rect 8757 8443 8815 8449
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 9692 8489 9720 8520
rect 9858 8508 9864 8560
rect 9916 8508 9922 8560
rect 10410 8548 10416 8560
rect 10060 8520 10416 8548
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8449 9735 8483
rect 9677 8443 9735 8449
rect 9769 8483 9827 8489
rect 9769 8449 9781 8483
rect 9815 8480 9827 8483
rect 9876 8480 9904 8508
rect 9815 8452 9904 8480
rect 9953 8483 10011 8489
rect 9815 8449 9827 8452
rect 9769 8443 9827 8449
rect 9953 8449 9965 8483
rect 9999 8478 10011 8483
rect 10060 8478 10088 8520
rect 10410 8508 10416 8520
rect 10468 8508 10474 8560
rect 10226 8480 10232 8492
rect 9999 8450 10088 8478
rect 10187 8452 10232 8480
rect 9999 8449 10011 8450
rect 9953 8443 10011 8449
rect 10226 8440 10232 8452
rect 10284 8440 10290 8492
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8480 10747 8483
rect 11146 8480 11152 8492
rect 10735 8452 11152 8480
rect 10735 8449 10747 8452
rect 10689 8443 10747 8449
rect 11146 8440 11152 8452
rect 11204 8440 11210 8492
rect 11330 8480 11336 8492
rect 11291 8452 11336 8480
rect 11330 8440 11336 8452
rect 11388 8480 11394 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 11388 8452 11529 8480
rect 11388 8440 11394 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 11790 8440 11796 8492
rect 11848 8480 11854 8492
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 11848 8452 12449 8480
rect 11848 8440 11854 8452
rect 12437 8449 12449 8452
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 12710 8440 12716 8492
rect 12768 8480 12774 8492
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 12768 8452 13185 8480
rect 12768 8440 12774 8452
rect 13173 8449 13185 8452
rect 13219 8449 13231 8483
rect 13173 8443 13231 8449
rect 7616 8384 7880 8412
rect 9585 8415 9643 8421
rect 7616 8372 7622 8384
rect 9585 8381 9597 8415
rect 9631 8412 9643 8415
rect 9858 8412 9864 8424
rect 9631 8384 9864 8412
rect 9631 8381 9643 8384
rect 9585 8375 9643 8381
rect 9858 8372 9864 8384
rect 9916 8412 9922 8424
rect 10597 8415 10655 8421
rect 10597 8412 10609 8415
rect 9916 8384 10609 8412
rect 9916 8372 9922 8384
rect 10597 8381 10609 8384
rect 10643 8381 10655 8415
rect 10778 8412 10784 8424
rect 10739 8384 10784 8412
rect 10597 8375 10655 8381
rect 10778 8372 10784 8384
rect 10836 8372 10842 8424
rect 10873 8347 10931 8353
rect 10873 8344 10885 8347
rect 7116 8316 9628 8344
rect 5721 8307 5779 8313
rect 6454 8276 6460 8288
rect 6415 8248 6460 8276
rect 6454 8236 6460 8248
rect 6512 8236 6518 8288
rect 7466 8236 7472 8288
rect 7524 8276 7530 8288
rect 7834 8276 7840 8288
rect 7524 8248 7840 8276
rect 7524 8236 7530 8248
rect 7834 8236 7840 8248
rect 7892 8276 7898 8288
rect 8846 8276 8852 8288
rect 7892 8248 8852 8276
rect 7892 8236 7898 8248
rect 8846 8236 8852 8248
rect 8904 8236 8910 8288
rect 9306 8276 9312 8288
rect 9267 8248 9312 8276
rect 9306 8236 9312 8248
rect 9364 8236 9370 8288
rect 9600 8276 9628 8316
rect 9784 8316 10885 8344
rect 9784 8276 9812 8316
rect 10873 8313 10885 8316
rect 10919 8344 10931 8347
rect 12805 8347 12863 8353
rect 12805 8344 12817 8347
rect 10919 8316 12817 8344
rect 10919 8313 10931 8316
rect 10873 8307 10931 8313
rect 12805 8313 12817 8316
rect 12851 8313 12863 8347
rect 12805 8307 12863 8313
rect 9600 8248 9812 8276
rect 9950 8236 9956 8288
rect 10008 8276 10014 8288
rect 10137 8279 10195 8285
rect 10137 8276 10149 8279
rect 10008 8248 10149 8276
rect 10008 8236 10014 8248
rect 10137 8245 10149 8248
rect 10183 8245 10195 8279
rect 13354 8276 13360 8288
rect 13315 8248 13360 8276
rect 10137 8239 10195 8245
rect 13354 8236 13360 8248
rect 13412 8236 13418 8288
rect 1104 8186 13892 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 12214 8186
rect 12266 8134 12278 8186
rect 12330 8134 12342 8186
rect 12394 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 13892 8186
rect 1104 8112 13892 8134
rect 1578 8032 1584 8084
rect 1636 8072 1642 8084
rect 2133 8075 2191 8081
rect 2133 8072 2145 8075
rect 1636 8044 2145 8072
rect 1636 8032 1642 8044
rect 2133 8041 2145 8044
rect 2179 8041 2191 8075
rect 2133 8035 2191 8041
rect 4341 8075 4399 8081
rect 4341 8041 4353 8075
rect 4387 8072 4399 8075
rect 4614 8072 4620 8084
rect 4387 8044 4620 8072
rect 4387 8041 4399 8044
rect 4341 8035 4399 8041
rect 1486 7936 1492 7948
rect 1447 7908 1492 7936
rect 1486 7896 1492 7908
rect 1544 7896 1550 7948
rect 1670 7936 1676 7948
rect 1631 7908 1676 7936
rect 1670 7896 1676 7908
rect 1728 7896 1734 7948
rect 2148 7936 2176 8035
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 7469 8075 7527 8081
rect 7469 8041 7481 8075
rect 7515 8072 7527 8075
rect 8570 8072 8576 8084
rect 7515 8044 8576 8072
rect 7515 8041 7527 8044
rect 7469 8035 7527 8041
rect 8570 8032 8576 8044
rect 8628 8072 8634 8084
rect 9122 8072 9128 8084
rect 8628 8044 9128 8072
rect 8628 8032 8634 8044
rect 9122 8032 9128 8044
rect 9180 8032 9186 8084
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 9950 8072 9956 8084
rect 9732 8044 9956 8072
rect 9732 8032 9738 8044
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 10965 8075 11023 8081
rect 10965 8072 10977 8075
rect 10836 8044 10977 8072
rect 10836 8032 10842 8044
rect 10965 8041 10977 8044
rect 11011 8041 11023 8075
rect 10965 8035 11023 8041
rect 3053 8007 3111 8013
rect 3053 7973 3065 8007
rect 3099 8004 3111 8007
rect 3326 8004 3332 8016
rect 3099 7976 3332 8004
rect 3099 7973 3111 7976
rect 3053 7967 3111 7973
rect 3326 7964 3332 7976
rect 3384 7964 3390 8016
rect 4157 8007 4215 8013
rect 4157 7973 4169 8007
rect 4203 8004 4215 8007
rect 4798 8004 4804 8016
rect 4203 7976 4804 8004
rect 4203 7973 4215 7976
rect 4157 7967 4215 7973
rect 4798 7964 4804 7976
rect 4856 7964 4862 8016
rect 5350 8004 5356 8016
rect 5311 7976 5356 8004
rect 5350 7964 5356 7976
rect 5408 7964 5414 8016
rect 8941 8007 8999 8013
rect 8941 8004 8953 8007
rect 7300 7976 8953 8004
rect 2225 7939 2283 7945
rect 2225 7936 2237 7939
rect 2148 7908 2237 7936
rect 2225 7905 2237 7908
rect 2271 7905 2283 7939
rect 2225 7899 2283 7905
rect 2961 7939 3019 7945
rect 2961 7905 2973 7939
rect 3007 7936 3019 7939
rect 3418 7936 3424 7948
rect 3007 7908 3424 7936
rect 3007 7905 3019 7908
rect 2961 7899 3019 7905
rect 3418 7896 3424 7908
rect 3476 7896 3482 7948
rect 3513 7939 3571 7945
rect 3513 7905 3525 7939
rect 3559 7936 3571 7939
rect 4062 7936 4068 7948
rect 3559 7908 4068 7936
rect 3559 7905 3571 7908
rect 3513 7899 3571 7905
rect 4062 7896 4068 7908
rect 4120 7896 4126 7948
rect 4890 7936 4896 7948
rect 4632 7908 4896 7936
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7868 2743 7871
rect 3142 7868 3148 7880
rect 2731 7840 3148 7868
rect 2731 7837 2743 7840
rect 2685 7831 2743 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7868 3847 7871
rect 3878 7868 3884 7880
rect 3835 7840 3884 7868
rect 3835 7837 3847 7840
rect 3789 7831 3847 7837
rect 3878 7828 3884 7840
rect 3936 7868 3942 7880
rect 4632 7877 4660 7908
rect 4890 7896 4896 7908
rect 4948 7896 4954 7948
rect 5445 7939 5503 7945
rect 5445 7905 5457 7939
rect 5491 7936 5503 7939
rect 6454 7936 6460 7948
rect 5491 7908 6460 7936
rect 5491 7905 5503 7908
rect 5445 7899 5503 7905
rect 6454 7896 6460 7908
rect 6512 7896 6518 7948
rect 6546 7896 6552 7948
rect 6604 7936 6610 7948
rect 7300 7945 7328 7976
rect 8941 7973 8953 7976
rect 8987 7973 8999 8007
rect 13262 8004 13268 8016
rect 13223 7976 13268 8004
rect 8941 7967 8999 7973
rect 13262 7964 13268 7976
rect 13320 7964 13326 8016
rect 6825 7939 6883 7945
rect 6825 7936 6837 7939
rect 6604 7908 6837 7936
rect 6604 7896 6610 7908
rect 6825 7905 6837 7908
rect 6871 7905 6883 7939
rect 6825 7899 6883 7905
rect 7285 7939 7343 7945
rect 7285 7905 7297 7939
rect 7331 7905 7343 7939
rect 7285 7899 7343 7905
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7936 7527 7939
rect 7561 7939 7619 7945
rect 7561 7936 7573 7939
rect 7515 7908 7573 7936
rect 7515 7905 7527 7908
rect 7469 7899 7527 7905
rect 7561 7905 7573 7908
rect 7607 7905 7619 7939
rect 7561 7899 7619 7905
rect 4433 7871 4491 7877
rect 4433 7868 4445 7871
rect 3936 7840 4445 7868
rect 3936 7828 3942 7840
rect 4433 7837 4445 7840
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 5718 7868 5724 7880
rect 5679 7840 5724 7868
rect 4617 7831 4675 7837
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 5997 7871 6055 7877
rect 5997 7837 6009 7871
rect 6043 7868 6055 7871
rect 6564 7868 6592 7896
rect 6043 7840 6592 7868
rect 6641 7871 6699 7877
rect 6043 7837 6055 7840
rect 5997 7831 6055 7837
rect 6641 7837 6653 7871
rect 6687 7868 6699 7871
rect 7300 7868 7328 7899
rect 8018 7896 8024 7948
rect 8076 7896 8082 7948
rect 8662 7936 8668 7948
rect 8623 7908 8668 7936
rect 8662 7896 8668 7908
rect 8720 7896 8726 7948
rect 8846 7896 8852 7948
rect 8904 7936 8910 7948
rect 9493 7939 9551 7945
rect 9493 7936 9505 7939
rect 8904 7908 9505 7936
rect 8904 7896 8910 7908
rect 9493 7905 9505 7908
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 9824 7908 10088 7936
rect 9824 7896 9830 7908
rect 6687 7840 7328 7868
rect 7745 7871 7803 7877
rect 6687 7837 6699 7840
rect 6641 7831 6699 7837
rect 7745 7837 7757 7871
rect 7791 7868 7803 7871
rect 7926 7868 7932 7880
rect 7791 7840 7932 7868
rect 7791 7837 7803 7840
rect 7745 7831 7803 7837
rect 7926 7828 7932 7840
rect 7984 7828 7990 7880
rect 8036 7868 8064 7896
rect 8205 7871 8263 7877
rect 8205 7870 8217 7871
rect 8128 7868 8217 7870
rect 8036 7842 8217 7868
rect 8036 7840 8156 7842
rect 8205 7837 8217 7842
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7868 8815 7871
rect 8938 7868 8944 7880
rect 8803 7840 8944 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 9306 7868 9312 7880
rect 9267 7840 9312 7868
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 9858 7868 9864 7880
rect 9819 7840 9864 7868
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 10060 7877 10088 7908
rect 10226 7896 10232 7948
rect 10284 7936 10290 7948
rect 10870 7936 10876 7948
rect 10284 7908 10876 7936
rect 10284 7896 10290 7908
rect 10520 7877 10548 7908
rect 10870 7896 10876 7908
rect 10928 7936 10934 7948
rect 11241 7939 11299 7945
rect 11241 7936 11253 7939
rect 10928 7908 11008 7936
rect 10928 7896 10934 7908
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7837 10103 7871
rect 10045 7831 10103 7837
rect 10505 7871 10563 7877
rect 10505 7837 10517 7871
rect 10551 7837 10563 7871
rect 10505 7831 10563 7837
rect 10594 7828 10600 7880
rect 10652 7828 10658 7880
rect 1762 7800 1768 7812
rect 1723 7772 1768 7800
rect 1762 7760 1768 7772
rect 1820 7760 1826 7812
rect 2777 7803 2835 7809
rect 2777 7769 2789 7803
rect 2823 7800 2835 7803
rect 3050 7800 3056 7812
rect 2823 7772 3056 7800
rect 2823 7769 2835 7772
rect 2777 7763 2835 7769
rect 3050 7760 3056 7772
rect 3108 7760 3114 7812
rect 6730 7800 6736 7812
rect 6691 7772 6736 7800
rect 6730 7760 6736 7772
rect 6788 7760 6794 7812
rect 8021 7803 8079 7809
rect 8021 7769 8033 7803
rect 8067 7769 8079 7803
rect 8021 7763 8079 7769
rect 4157 7735 4215 7741
rect 4157 7701 4169 7735
rect 4203 7732 4215 7735
rect 4430 7732 4436 7744
rect 4203 7704 4436 7732
rect 4203 7701 4215 7704
rect 4157 7695 4215 7701
rect 4430 7692 4436 7704
rect 4488 7732 4494 7744
rect 5350 7732 5356 7744
rect 4488 7704 5356 7732
rect 4488 7692 4494 7704
rect 5350 7692 5356 7704
rect 5408 7692 5414 7744
rect 7558 7692 7564 7744
rect 7616 7732 7622 7744
rect 8036 7732 8064 7763
rect 8110 7760 8116 7812
rect 8168 7800 8174 7812
rect 9214 7800 9220 7812
rect 8168 7772 9220 7800
rect 8168 7760 8174 7772
rect 9214 7760 9220 7772
rect 9272 7760 9278 7812
rect 9401 7803 9459 7809
rect 9401 7769 9413 7803
rect 9447 7800 9459 7803
rect 10612 7800 10640 7828
rect 9447 7772 10640 7800
rect 9447 7769 9459 7772
rect 9401 7763 9459 7769
rect 7616 7704 8064 7732
rect 8297 7735 8355 7741
rect 7616 7692 7622 7704
rect 8297 7701 8309 7735
rect 8343 7732 8355 7735
rect 8754 7732 8760 7744
rect 8343 7704 8760 7732
rect 8343 7701 8355 7704
rect 8297 7695 8355 7701
rect 8754 7692 8760 7704
rect 8812 7692 8818 7744
rect 8846 7692 8852 7744
rect 8904 7732 8910 7744
rect 9674 7732 9680 7744
rect 8904 7704 9680 7732
rect 8904 7692 8910 7704
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 9858 7732 9864 7744
rect 9819 7704 9864 7732
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 10042 7692 10048 7744
rect 10100 7732 10106 7744
rect 10410 7732 10416 7744
rect 10100 7704 10416 7732
rect 10100 7692 10106 7704
rect 10410 7692 10416 7704
rect 10468 7732 10474 7744
rect 10597 7735 10655 7741
rect 10597 7732 10609 7735
rect 10468 7704 10609 7732
rect 10468 7692 10474 7704
rect 10597 7701 10609 7704
rect 10643 7701 10655 7735
rect 10980 7732 11008 7908
rect 11072 7908 11253 7936
rect 11072 7877 11100 7908
rect 11241 7905 11253 7908
rect 11287 7936 11299 7939
rect 11287 7908 12020 7936
rect 11287 7905 11299 7908
rect 11241 7899 11299 7905
rect 11992 7877 12020 7908
rect 12618 7896 12624 7948
rect 12676 7936 12682 7948
rect 12805 7939 12863 7945
rect 12805 7936 12817 7939
rect 12676 7908 12817 7936
rect 12676 7896 12682 7908
rect 12805 7905 12817 7908
rect 12851 7905 12863 7939
rect 13354 7936 13360 7948
rect 13315 7908 13360 7936
rect 12805 7899 12863 7905
rect 13354 7896 13360 7908
rect 13412 7896 13418 7948
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7837 11115 7871
rect 11057 7831 11115 7837
rect 11701 7871 11759 7877
rect 11701 7837 11713 7871
rect 11747 7868 11759 7871
rect 11977 7871 12035 7877
rect 11747 7840 11928 7868
rect 11747 7837 11759 7840
rect 11701 7831 11759 7837
rect 11146 7800 11152 7812
rect 11107 7772 11152 7800
rect 11146 7760 11152 7772
rect 11204 7760 11210 7812
rect 11790 7800 11796 7812
rect 11751 7772 11796 7800
rect 11790 7760 11796 7772
rect 11848 7760 11854 7812
rect 11900 7800 11928 7840
rect 11977 7837 11989 7871
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 12713 7871 12771 7877
rect 12713 7837 12725 7871
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 12250 7800 12256 7812
rect 11900 7772 12256 7800
rect 12250 7760 12256 7772
rect 12308 7800 12314 7812
rect 12728 7800 12756 7831
rect 12308 7772 12756 7800
rect 12308 7760 12314 7772
rect 13354 7732 13360 7744
rect 10980 7704 13360 7732
rect 10597 7695 10655 7701
rect 13354 7692 13360 7704
rect 13412 7692 13418 7744
rect 1104 7642 13892 7664
rect 1104 7590 8214 7642
rect 8266 7590 8278 7642
rect 8330 7590 8342 7642
rect 8394 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 13892 7642
rect 1104 7568 13892 7590
rect 3050 7528 3056 7540
rect 3011 7500 3056 7528
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 3145 7531 3203 7537
rect 3145 7497 3157 7531
rect 3191 7528 3203 7531
rect 3326 7528 3332 7540
rect 3191 7500 3332 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 3326 7488 3332 7500
rect 3384 7488 3390 7540
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 6730 7528 6736 7540
rect 6687 7500 6736 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 7466 7528 7472 7540
rect 6932 7500 7472 7528
rect 5258 7460 5264 7472
rect 2884 7432 5264 7460
rect 2884 7401 2912 7432
rect 5258 7420 5264 7432
rect 5316 7420 5322 7472
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7392 2467 7395
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 2455 7364 2605 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 2593 7361 2605 7364
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 2869 7395 2927 7401
rect 2869 7361 2881 7395
rect 2915 7361 2927 7395
rect 2869 7355 2927 7361
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7361 3663 7395
rect 3878 7392 3884 7404
rect 3839 7364 3884 7392
rect 3605 7355 3663 7361
rect 1486 7284 1492 7336
rect 1544 7324 1550 7336
rect 3620 7324 3648 7355
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 4430 7392 4436 7404
rect 4391 7364 4436 7392
rect 4430 7352 4436 7364
rect 4488 7352 4494 7404
rect 5718 7352 5724 7404
rect 5776 7392 5782 7404
rect 6932 7401 6960 7500
rect 7466 7488 7472 7500
rect 7524 7528 7530 7540
rect 7929 7531 7987 7537
rect 7929 7528 7941 7531
rect 7524 7500 7941 7528
rect 7524 7488 7530 7500
rect 7929 7497 7941 7500
rect 7975 7497 7987 7531
rect 7929 7491 7987 7497
rect 8021 7531 8079 7537
rect 8021 7497 8033 7531
rect 8067 7528 8079 7531
rect 8110 7528 8116 7540
rect 8067 7500 8116 7528
rect 8067 7497 8079 7500
rect 8021 7491 8079 7497
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 10318 7488 10324 7540
rect 10376 7528 10382 7540
rect 10873 7531 10931 7537
rect 10873 7528 10885 7531
rect 10376 7500 10885 7528
rect 10376 7488 10382 7500
rect 10873 7497 10885 7500
rect 10919 7528 10931 7531
rect 10962 7528 10968 7540
rect 10919 7500 10968 7528
rect 10919 7497 10931 7500
rect 10873 7491 10931 7497
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11146 7488 11152 7540
rect 11204 7528 11210 7540
rect 11977 7531 12035 7537
rect 11977 7528 11989 7531
rect 11204 7500 11989 7528
rect 11204 7488 11210 7500
rect 11977 7497 11989 7500
rect 12023 7497 12035 7531
rect 12250 7528 12256 7540
rect 12211 7500 12256 7528
rect 11977 7491 12035 7497
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 7190 7420 7196 7472
rect 7248 7460 7254 7472
rect 8665 7463 8723 7469
rect 8665 7460 8677 7463
rect 7248 7432 8677 7460
rect 7248 7420 7254 7432
rect 6457 7395 6515 7401
rect 6457 7392 6469 7395
rect 5776 7364 6469 7392
rect 5776 7352 5782 7364
rect 6457 7361 6469 7364
rect 6503 7361 6515 7395
rect 6457 7355 6515 7361
rect 6917 7395 6975 7401
rect 6917 7361 6929 7395
rect 6963 7361 6975 7395
rect 7282 7392 7288 7404
rect 7243 7364 7288 7392
rect 6917 7355 6975 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7392 7619 7395
rect 7650 7392 7656 7404
rect 7607 7364 7656 7392
rect 7607 7361 7619 7364
rect 7561 7355 7619 7361
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 1544 7296 3648 7324
rect 7101 7327 7159 7333
rect 1544 7284 1550 7296
rect 7101 7293 7113 7327
rect 7147 7293 7159 7327
rect 7101 7287 7159 7293
rect 7820 7327 7878 7333
rect 7820 7293 7832 7327
rect 7866 7324 7878 7327
rect 7944 7324 7972 7432
rect 8665 7429 8677 7432
rect 8711 7429 8723 7463
rect 8665 7423 8723 7429
rect 9214 7420 9220 7472
rect 9272 7460 9278 7472
rect 9493 7463 9551 7469
rect 9493 7460 9505 7463
rect 9272 7432 9505 7460
rect 9272 7420 9278 7432
rect 9493 7429 9505 7432
rect 9539 7429 9551 7463
rect 9493 7423 9551 7429
rect 9950 7420 9956 7472
rect 10008 7460 10014 7472
rect 10008 7432 10180 7460
rect 10008 7420 10014 7432
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 8570 7392 8576 7404
rect 8444 7364 8489 7392
rect 8531 7364 8576 7392
rect 8444 7352 8450 7364
rect 8570 7352 8576 7364
rect 8628 7352 8634 7404
rect 8846 7401 8852 7404
rect 8809 7395 8852 7401
rect 8809 7361 8821 7395
rect 8809 7355 8852 7361
rect 8846 7352 8852 7355
rect 8904 7352 8910 7404
rect 9030 7352 9036 7404
rect 9088 7392 9094 7404
rect 9125 7395 9183 7401
rect 9125 7392 9137 7395
rect 9088 7364 9137 7392
rect 9088 7352 9094 7364
rect 9125 7361 9137 7364
rect 9171 7361 9183 7395
rect 9125 7355 9183 7361
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7392 9367 7395
rect 9398 7392 9404 7404
rect 9355 7364 9404 7392
rect 9355 7361 9367 7364
rect 9309 7355 9367 7361
rect 9398 7352 9404 7364
rect 9456 7392 9462 7404
rect 9677 7395 9735 7401
rect 9677 7392 9689 7395
rect 9456 7364 9689 7392
rect 9456 7352 9462 7364
rect 9677 7361 9689 7364
rect 9723 7361 9735 7395
rect 9858 7392 9864 7404
rect 9819 7364 9864 7392
rect 9677 7355 9735 7361
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 10152 7401 10180 7432
rect 10502 7420 10508 7472
rect 10560 7460 10566 7472
rect 12621 7463 12679 7469
rect 12621 7460 12633 7463
rect 10560 7432 12633 7460
rect 10560 7420 10566 7432
rect 12621 7429 12633 7432
rect 12667 7429 12679 7463
rect 12621 7423 12679 7429
rect 10137 7395 10195 7401
rect 10137 7361 10149 7395
rect 10183 7361 10195 7395
rect 10137 7355 10195 7361
rect 10226 7352 10232 7404
rect 10284 7392 10290 7404
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 10284 7364 10333 7392
rect 10284 7352 10290 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 10870 7352 10876 7404
rect 10928 7392 10934 7404
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 10928 7364 11529 7392
rect 10928 7352 10934 7364
rect 11517 7361 11529 7364
rect 11563 7361 11575 7395
rect 11517 7355 11575 7361
rect 11790 7352 11796 7404
rect 11848 7392 11854 7404
rect 12161 7395 12219 7401
rect 12161 7392 12173 7395
rect 11848 7364 12173 7392
rect 11848 7352 11854 7364
rect 12161 7361 12173 7364
rect 12207 7361 12219 7395
rect 12161 7355 12219 7361
rect 12713 7395 12771 7401
rect 12713 7361 12725 7395
rect 12759 7392 12771 7395
rect 12894 7392 12900 7404
rect 12759 7364 12900 7392
rect 12759 7361 12771 7364
rect 12713 7355 12771 7361
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 13354 7392 13360 7404
rect 13315 7364 13360 7392
rect 13354 7352 13360 7364
rect 13412 7352 13418 7404
rect 7866 7296 7972 7324
rect 8113 7327 8171 7333
rect 7866 7293 7878 7296
rect 7820 7287 7878 7293
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8938 7324 8944 7336
rect 8159 7296 8944 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 2409 7259 2467 7265
rect 2409 7225 2421 7259
rect 2455 7256 2467 7259
rect 3142 7256 3148 7268
rect 2455 7228 3148 7256
rect 2455 7225 2467 7228
rect 2409 7219 2467 7225
rect 3142 7216 3148 7228
rect 3200 7216 3206 7268
rect 3881 7259 3939 7265
rect 3881 7225 3893 7259
rect 3927 7256 3939 7259
rect 5350 7256 5356 7268
rect 3927 7228 5356 7256
rect 3927 7225 3939 7228
rect 3881 7219 3939 7225
rect 2590 7148 2596 7200
rect 2648 7188 2654 7200
rect 3896 7188 3924 7219
rect 5350 7216 5356 7228
rect 5408 7216 5414 7268
rect 7006 7256 7012 7268
rect 6967 7228 7012 7256
rect 7006 7216 7012 7228
rect 7064 7216 7070 7268
rect 7116 7256 7144 7287
rect 8938 7284 8944 7296
rect 8996 7284 9002 7336
rect 9950 7324 9956 7336
rect 9911 7296 9956 7324
rect 9950 7284 9956 7296
rect 10008 7284 10014 7336
rect 10045 7327 10103 7333
rect 10045 7293 10057 7327
rect 10091 7293 10103 7327
rect 10045 7287 10103 7293
rect 10413 7327 10471 7333
rect 10413 7293 10425 7327
rect 10459 7324 10471 7327
rect 10965 7327 11023 7333
rect 10965 7324 10977 7327
rect 10459 7296 10977 7324
rect 10459 7293 10471 7296
rect 10413 7287 10471 7293
rect 10965 7293 10977 7296
rect 11011 7293 11023 7327
rect 10965 7287 11023 7293
rect 11057 7327 11115 7333
rect 11057 7293 11069 7327
rect 11103 7293 11115 7327
rect 12802 7324 12808 7336
rect 12763 7296 12808 7324
rect 11057 7287 11115 7293
rect 8754 7256 8760 7268
rect 7116 7228 8760 7256
rect 8754 7216 8760 7228
rect 8812 7216 8818 7268
rect 8846 7216 8852 7268
rect 8904 7256 8910 7268
rect 8904 7228 9536 7256
rect 8904 7216 8910 7228
rect 9508 7200 9536 7228
rect 9766 7216 9772 7268
rect 9824 7256 9830 7268
rect 10060 7256 10088 7287
rect 10870 7256 10876 7268
rect 9824 7228 10876 7256
rect 9824 7216 9830 7228
rect 10870 7216 10876 7228
rect 10928 7256 10934 7268
rect 11072 7256 11100 7287
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 10928 7228 11100 7256
rect 10928 7216 10934 7228
rect 2648 7160 3924 7188
rect 4433 7191 4491 7197
rect 2648 7148 2654 7160
rect 4433 7157 4445 7191
rect 4479 7188 4491 7191
rect 4614 7188 4620 7200
rect 4479 7160 4620 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 5074 7148 5080 7200
rect 5132 7188 5138 7200
rect 7377 7191 7435 7197
rect 7377 7188 7389 7191
rect 5132 7160 7389 7188
rect 5132 7148 5138 7160
rect 7377 7157 7389 7160
rect 7423 7157 7435 7191
rect 7377 7151 7435 7157
rect 8941 7191 8999 7197
rect 8941 7157 8953 7191
rect 8987 7188 8999 7191
rect 9030 7188 9036 7200
rect 8987 7160 9036 7188
rect 8987 7157 8999 7160
rect 8941 7151 8999 7157
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 9490 7148 9496 7200
rect 9548 7188 9554 7200
rect 10413 7191 10471 7197
rect 10413 7188 10425 7191
rect 9548 7160 10425 7188
rect 9548 7148 9554 7160
rect 10413 7157 10425 7160
rect 10459 7157 10471 7191
rect 10413 7151 10471 7157
rect 10505 7191 10563 7197
rect 10505 7157 10517 7191
rect 10551 7188 10563 7191
rect 10778 7188 10784 7200
rect 10551 7160 10784 7188
rect 10551 7157 10563 7160
rect 10505 7151 10563 7157
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 11330 7148 11336 7200
rect 11388 7188 11394 7200
rect 11609 7191 11667 7197
rect 11609 7188 11621 7191
rect 11388 7160 11621 7188
rect 11388 7148 11394 7160
rect 11609 7157 11621 7160
rect 11655 7157 11667 7191
rect 13170 7188 13176 7200
rect 13131 7160 13176 7188
rect 11609 7151 11667 7157
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 1104 7098 13892 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 12214 7098
rect 12266 7046 12278 7098
rect 12330 7046 12342 7098
rect 12394 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 13892 7098
rect 1104 7024 13892 7046
rect 3878 6984 3884 6996
rect 3839 6956 3884 6984
rect 3878 6944 3884 6956
rect 3936 6944 3942 6996
rect 5074 6993 5080 6996
rect 5064 6987 5080 6993
rect 5064 6953 5076 6987
rect 5064 6947 5080 6953
rect 5074 6944 5080 6947
rect 5132 6944 5138 6996
rect 6549 6987 6607 6993
rect 6549 6953 6561 6987
rect 6595 6984 6607 6987
rect 7190 6984 7196 6996
rect 6595 6956 7196 6984
rect 6595 6953 6607 6956
rect 6549 6947 6607 6953
rect 7190 6944 7196 6956
rect 7248 6944 7254 6996
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 7377 6987 7435 6993
rect 7377 6984 7389 6987
rect 7340 6956 7389 6984
rect 7340 6944 7346 6956
rect 7377 6953 7389 6956
rect 7423 6953 7435 6987
rect 7377 6947 7435 6953
rect 8662 6944 8668 6996
rect 8720 6944 8726 6996
rect 9858 6944 9864 6996
rect 9916 6984 9922 6996
rect 10410 6984 10416 6996
rect 9916 6956 10416 6984
rect 9916 6944 9922 6956
rect 10410 6944 10416 6956
rect 10468 6944 10474 6996
rect 12618 6944 12624 6996
rect 12676 6984 12682 6996
rect 12805 6987 12863 6993
rect 12805 6984 12817 6987
rect 12676 6956 12817 6984
rect 12676 6944 12682 6956
rect 12805 6953 12817 6956
rect 12851 6953 12863 6987
rect 12805 6947 12863 6953
rect 6914 6876 6920 6928
rect 6972 6916 6978 6928
rect 7558 6916 7564 6928
rect 6972 6888 7564 6916
rect 6972 6876 6978 6888
rect 7558 6876 7564 6888
rect 7616 6876 7622 6928
rect 7926 6876 7932 6928
rect 7984 6916 7990 6928
rect 8386 6916 8392 6928
rect 7984 6888 8392 6916
rect 7984 6876 7990 6888
rect 8386 6876 8392 6888
rect 8444 6876 8450 6928
rect 8680 6916 8708 6944
rect 10042 6916 10048 6928
rect 8680 6888 9536 6916
rect 10003 6888 10048 6916
rect 6825 6851 6883 6857
rect 6825 6817 6837 6851
rect 6871 6848 6883 6851
rect 6871 6820 7696 6848
rect 6871 6817 6883 6820
rect 6825 6811 6883 6817
rect 2590 6780 2596 6792
rect 2551 6752 2596 6780
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6780 3387 6783
rect 3418 6780 3424 6792
rect 3375 6752 3424 6780
rect 3375 6749 3387 6752
rect 3329 6743 3387 6749
rect 3418 6740 3424 6752
rect 3476 6740 3482 6792
rect 3694 6740 3700 6792
rect 3752 6780 3758 6792
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 3752 6752 3801 6780
rect 3752 6740 3758 6752
rect 3789 6749 3801 6752
rect 3835 6749 3847 6783
rect 3970 6780 3976 6792
rect 3931 6752 3976 6780
rect 3789 6743 3847 6749
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4798 6780 4804 6792
rect 4759 6752 4804 6780
rect 4798 6740 4804 6752
rect 4856 6740 4862 6792
rect 6914 6780 6920 6792
rect 6875 6752 6920 6780
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 7558 6789 7564 6792
rect 7193 6783 7251 6789
rect 7193 6780 7205 6783
rect 7024 6752 7205 6780
rect 5810 6672 5816 6724
rect 5868 6672 5874 6724
rect 2774 6604 2780 6656
rect 2832 6644 2838 6656
rect 2832 6616 2877 6644
rect 2832 6604 2838 6616
rect 2958 6604 2964 6656
rect 3016 6644 3022 6656
rect 3237 6647 3295 6653
rect 3237 6644 3249 6647
rect 3016 6616 3249 6644
rect 3016 6604 3022 6616
rect 3237 6613 3249 6616
rect 3283 6613 3295 6647
rect 7024 6644 7052 6752
rect 7193 6749 7205 6752
rect 7239 6749 7251 6783
rect 7556 6780 7564 6789
rect 7519 6752 7564 6780
rect 7193 6743 7251 6749
rect 7556 6743 7564 6752
rect 7558 6740 7564 6743
rect 7616 6740 7622 6792
rect 7668 6780 7696 6820
rect 7742 6808 7748 6860
rect 7800 6848 7806 6860
rect 8404 6848 8432 6876
rect 7800 6820 8064 6848
rect 8404 6820 8524 6848
rect 7800 6808 7806 6820
rect 8036 6789 8064 6820
rect 7873 6783 7931 6789
rect 7873 6780 7885 6783
rect 7668 6752 7885 6780
rect 7873 6749 7885 6752
rect 7919 6749 7931 6783
rect 7873 6743 7931 6749
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 8110 6740 8116 6792
rect 8168 6780 8174 6792
rect 8496 6789 8524 6820
rect 8570 6808 8576 6860
rect 8628 6848 8634 6860
rect 8665 6851 8723 6857
rect 8665 6848 8677 6851
rect 8628 6820 8677 6848
rect 8628 6808 8634 6820
rect 8665 6817 8677 6820
rect 8711 6817 8723 6851
rect 8665 6811 8723 6817
rect 8754 6808 8760 6860
rect 8812 6848 8818 6860
rect 9398 6848 9404 6860
rect 8812 6820 8857 6848
rect 8956 6820 9404 6848
rect 8812 6808 8818 6820
rect 8389 6783 8447 6789
rect 8389 6780 8401 6783
rect 8168 6752 8401 6780
rect 8168 6740 8174 6752
rect 8389 6749 8401 6752
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 8481 6783 8539 6789
rect 8481 6749 8493 6783
rect 8527 6749 8539 6783
rect 8481 6743 8539 6749
rect 8846 6740 8852 6792
rect 8904 6780 8910 6792
rect 8956 6780 8984 6820
rect 9398 6808 9404 6820
rect 9456 6808 9462 6860
rect 9508 6857 9536 6888
rect 10042 6876 10048 6888
rect 10100 6876 10106 6928
rect 10226 6876 10232 6928
rect 10284 6916 10290 6928
rect 11793 6919 11851 6925
rect 10284 6888 11100 6916
rect 10284 6876 10290 6888
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6817 9551 6851
rect 10244 6848 10272 6876
rect 9493 6811 9551 6817
rect 9692 6820 10272 6848
rect 8904 6752 8984 6780
rect 8904 6740 8910 6752
rect 9030 6740 9036 6792
rect 9088 6780 9094 6792
rect 9692 6789 9720 6820
rect 9217 6783 9275 6789
rect 9217 6780 9229 6783
rect 9088 6752 9229 6780
rect 9088 6740 9094 6752
rect 9217 6749 9229 6752
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 9309 6783 9367 6789
rect 9309 6749 9321 6783
rect 9355 6749 9367 6783
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9309 6743 9367 6749
rect 9416 6752 9689 6780
rect 7101 6715 7159 6721
rect 7101 6681 7113 6715
rect 7147 6712 7159 6715
rect 7653 6715 7711 6721
rect 7653 6712 7665 6715
rect 7147 6684 7665 6712
rect 7147 6681 7159 6684
rect 7101 6675 7159 6681
rect 7653 6681 7665 6684
rect 7699 6681 7711 6715
rect 7653 6675 7711 6681
rect 7745 6715 7803 6721
rect 7745 6681 7757 6715
rect 7791 6712 7803 6715
rect 8205 6715 8263 6721
rect 8205 6712 8217 6715
rect 7791 6684 8217 6712
rect 7791 6681 7803 6684
rect 7745 6675 7803 6681
rect 8205 6681 8217 6684
rect 8251 6712 8263 6715
rect 9324 6712 9352 6743
rect 9416 6724 9444 6752
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 10177 6783 10235 6789
rect 10177 6780 10189 6783
rect 9677 6743 9735 6749
rect 9784 6752 10189 6780
rect 8251 6684 9352 6712
rect 8251 6681 8263 6684
rect 8205 6675 8263 6681
rect 7760 6644 7788 6675
rect 9398 6672 9404 6724
rect 9456 6672 9462 6724
rect 9490 6672 9496 6724
rect 9548 6712 9554 6724
rect 9784 6712 9812 6752
rect 10177 6749 10189 6752
rect 10223 6749 10235 6783
rect 10177 6743 10235 6749
rect 10318 6740 10324 6792
rect 10376 6780 10382 6792
rect 10612 6789 10640 6888
rect 10689 6851 10747 6857
rect 10689 6817 10701 6851
rect 10735 6848 10747 6851
rect 10735 6820 10916 6848
rect 10735 6817 10747 6820
rect 10689 6811 10747 6817
rect 10597 6783 10655 6789
rect 10376 6752 10421 6780
rect 10376 6740 10382 6752
rect 10597 6749 10609 6783
rect 10643 6749 10655 6783
rect 10778 6780 10784 6792
rect 10739 6752 10784 6780
rect 10597 6743 10655 6749
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 10888 6780 10916 6820
rect 11072 6789 11100 6888
rect 11793 6885 11805 6919
rect 11839 6885 11851 6919
rect 11793 6879 11851 6885
rect 11425 6851 11483 6857
rect 11425 6817 11437 6851
rect 11471 6848 11483 6851
rect 11808 6848 11836 6879
rect 11471 6820 11836 6848
rect 11471 6817 11483 6820
rect 11425 6811 11483 6817
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 10888 6752 10977 6780
rect 10965 6749 10977 6752
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 11183 6783 11241 6789
rect 11183 6749 11195 6783
rect 11229 6780 11241 6783
rect 11330 6780 11336 6792
rect 11229 6752 11336 6780
rect 11229 6749 11241 6752
rect 11183 6743 11241 6749
rect 11330 6740 11336 6752
rect 11388 6740 11394 6792
rect 9548 6684 9812 6712
rect 10413 6715 10471 6721
rect 9548 6672 9554 6684
rect 10413 6681 10425 6715
rect 10459 6712 10471 6715
rect 10459 6684 10824 6712
rect 10459 6681 10471 6684
rect 10413 6675 10471 6681
rect 10796 6656 10824 6684
rect 7024 6616 7788 6644
rect 9033 6647 9091 6653
rect 3237 6607 3295 6613
rect 9033 6613 9045 6647
rect 9079 6644 9091 6647
rect 9214 6644 9220 6656
rect 9079 6616 9220 6644
rect 9079 6613 9091 6616
rect 9033 6607 9091 6613
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 9950 6644 9956 6656
rect 9732 6616 9956 6644
rect 9732 6604 9738 6616
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 10226 6604 10232 6656
rect 10284 6644 10290 6656
rect 10689 6647 10747 6653
rect 10689 6644 10701 6647
rect 10284 6616 10701 6644
rect 10284 6604 10290 6616
rect 10689 6613 10701 6616
rect 10735 6613 10747 6647
rect 10689 6607 10747 6613
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 11348 6644 11376 6740
rect 10836 6616 11376 6644
rect 11532 6644 11560 6820
rect 12802 6808 12808 6860
rect 12860 6848 12866 6860
rect 13357 6851 13415 6857
rect 13357 6848 13369 6851
rect 12860 6820 13369 6848
rect 12860 6808 12866 6820
rect 13357 6817 13369 6820
rect 13403 6817 13415 6851
rect 13357 6811 13415 6817
rect 11606 6740 11612 6792
rect 11664 6780 11670 6792
rect 11701 6783 11759 6789
rect 11701 6780 11713 6783
rect 11664 6752 11713 6780
rect 11664 6740 11670 6752
rect 11701 6749 11713 6752
rect 11747 6780 11759 6783
rect 12223 6783 12281 6789
rect 12223 6780 12235 6783
rect 11747 6752 12235 6780
rect 11747 6749 11759 6752
rect 11701 6743 11759 6749
rect 12223 6749 12235 6752
rect 12269 6780 12281 6783
rect 12342 6780 12348 6792
rect 12269 6752 12348 6780
rect 12269 6749 12281 6752
rect 12223 6743 12281 6749
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 12529 6783 12587 6789
rect 12529 6749 12541 6783
rect 12575 6780 12587 6783
rect 12618 6780 12624 6792
rect 12575 6752 12624 6780
rect 12575 6749 12587 6752
rect 12529 6743 12587 6749
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 13170 6780 13176 6792
rect 13131 6752 13176 6780
rect 13170 6740 13176 6752
rect 13228 6740 13234 6792
rect 12161 6647 12219 6653
rect 12161 6644 12173 6647
rect 11532 6616 12173 6644
rect 10836 6604 10842 6616
rect 12161 6613 12173 6616
rect 12207 6613 12219 6647
rect 12161 6607 12219 6613
rect 12250 6604 12256 6656
rect 12308 6644 12314 6656
rect 12345 6647 12403 6653
rect 12345 6644 12357 6647
rect 12308 6616 12357 6644
rect 12308 6604 12314 6616
rect 12345 6613 12357 6616
rect 12391 6613 12403 6647
rect 12710 6644 12716 6656
rect 12671 6616 12716 6644
rect 12345 6607 12403 6613
rect 12710 6604 12716 6616
rect 12768 6604 12774 6656
rect 13262 6644 13268 6656
rect 13223 6616 13268 6644
rect 13262 6604 13268 6616
rect 13320 6604 13326 6656
rect 1104 6554 13892 6576
rect 1104 6502 8214 6554
rect 8266 6502 8278 6554
rect 8330 6502 8342 6554
rect 8394 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 13892 6554
rect 1104 6480 13892 6502
rect 2774 6400 2780 6452
rect 2832 6400 2838 6452
rect 5810 6440 5816 6452
rect 5771 6412 5816 6440
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6409 6239 6443
rect 8110 6440 8116 6452
rect 8071 6412 8116 6440
rect 6181 6403 6239 6409
rect 2792 6358 2820 6400
rect 6196 6372 6224 6403
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 8570 6400 8576 6452
rect 8628 6440 8634 6452
rect 9490 6440 9496 6452
rect 8628 6412 9496 6440
rect 8628 6400 8634 6412
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 10042 6400 10048 6452
rect 10100 6400 10106 6452
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 10413 6443 10471 6449
rect 10413 6440 10425 6443
rect 10284 6412 10425 6440
rect 10284 6400 10290 6412
rect 10413 6409 10425 6412
rect 10459 6409 10471 6443
rect 10413 6403 10471 6409
rect 12342 6400 12348 6452
rect 12400 6440 12406 6452
rect 13449 6443 13507 6449
rect 13449 6440 13461 6443
rect 12400 6412 13461 6440
rect 12400 6400 12406 6412
rect 13449 6409 13461 6412
rect 13495 6409 13507 6443
rect 13449 6403 13507 6409
rect 9674 6372 9680 6384
rect 6196 6344 7130 6372
rect 9600 6344 9680 6372
rect 3878 6304 3884 6316
rect 3839 6276 3884 6304
rect 3878 6264 3884 6276
rect 3936 6264 3942 6316
rect 4614 6304 4620 6316
rect 4575 6276 4620 6304
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 5350 6304 5356 6316
rect 5311 6276 5356 6304
rect 5350 6264 5356 6276
rect 5408 6304 5414 6316
rect 5629 6307 5687 6313
rect 5629 6304 5641 6307
rect 5408 6276 5641 6304
rect 5408 6264 5414 6276
rect 5629 6273 5641 6276
rect 5675 6304 5687 6307
rect 5902 6304 5908 6316
rect 5675 6276 5908 6304
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 5902 6264 5908 6276
rect 5960 6304 5966 6316
rect 5997 6307 6055 6313
rect 5997 6304 6009 6307
rect 5960 6276 6009 6304
rect 5960 6264 5966 6276
rect 5997 6273 6009 6276
rect 6043 6273 6055 6307
rect 5997 6267 6055 6273
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6304 8447 6307
rect 8662 6304 8668 6316
rect 8435 6276 8668 6304
rect 8435 6273 8447 6276
rect 8389 6267 8447 6273
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 8846 6304 8852 6316
rect 8807 6276 8852 6304
rect 8846 6264 8852 6276
rect 8904 6264 8910 6316
rect 9030 6304 9036 6316
rect 8991 6276 9036 6304
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9600 6313 9628 6344
rect 9674 6332 9680 6344
rect 9732 6332 9738 6384
rect 10060 6372 10088 6400
rect 10505 6375 10563 6381
rect 9968 6344 10439 6372
rect 9968 6328 9996 6344
rect 9784 6313 9996 6328
rect 9585 6307 9643 6313
rect 9585 6273 9597 6307
rect 9631 6273 9643 6307
rect 9585 6267 9643 6273
rect 9769 6307 9996 6313
rect 9769 6273 9781 6307
rect 9815 6300 9996 6307
rect 9815 6273 9827 6300
rect 9769 6267 9827 6273
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 10318 6313 10324 6316
rect 10301 6307 10324 6313
rect 10100 6276 10145 6304
rect 10100 6264 10106 6276
rect 10301 6273 10313 6307
rect 10301 6267 10324 6273
rect 10318 6264 10324 6267
rect 10376 6264 10382 6316
rect 10411 6304 10439 6344
rect 10505 6341 10517 6375
rect 10551 6372 10563 6375
rect 11057 6375 11115 6381
rect 11057 6372 11069 6375
rect 10551 6344 11069 6372
rect 10551 6341 10563 6344
rect 10505 6335 10563 6341
rect 11057 6341 11069 6344
rect 11103 6341 11115 6375
rect 11057 6335 11115 6341
rect 11977 6375 12035 6381
rect 11977 6341 11989 6375
rect 12023 6372 12035 6375
rect 12250 6372 12256 6384
rect 12023 6344 12256 6372
rect 12023 6341 12035 6344
rect 11977 6335 12035 6341
rect 12250 6332 12256 6344
rect 12308 6332 12314 6384
rect 12710 6332 12716 6384
rect 12768 6332 12774 6384
rect 10689 6307 10747 6313
rect 10689 6304 10701 6307
rect 10411 6276 10701 6304
rect 10689 6273 10701 6276
rect 10735 6273 10747 6307
rect 10689 6267 10747 6273
rect 10778 6264 10784 6316
rect 10836 6304 10842 6316
rect 10873 6307 10931 6313
rect 10873 6304 10885 6307
rect 10836 6276 10885 6304
rect 10836 6264 10842 6276
rect 10873 6273 10885 6276
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 11333 6307 11391 6313
rect 11333 6273 11345 6307
rect 11379 6273 11391 6307
rect 11333 6267 11391 6273
rect 1670 6236 1676 6248
rect 1631 6208 1676 6236
rect 1670 6196 1676 6208
rect 1728 6196 1734 6248
rect 1949 6239 2007 6245
rect 1949 6205 1961 6239
rect 1995 6236 2007 6239
rect 3234 6236 3240 6248
rect 1995 6208 3240 6236
rect 1995 6205 2007 6208
rect 1949 6199 2007 6205
rect 3234 6196 3240 6208
rect 3292 6196 3298 6248
rect 4798 6236 4804 6248
rect 4080 6208 4804 6236
rect 3050 6128 3056 6180
rect 3108 6168 3114 6180
rect 3789 6171 3847 6177
rect 3789 6168 3801 6171
rect 3108 6140 3801 6168
rect 3108 6128 3114 6140
rect 3789 6137 3801 6140
rect 3835 6137 3847 6171
rect 3789 6131 3847 6137
rect 3418 6100 3424 6112
rect 3379 6072 3424 6100
rect 3418 6060 3424 6072
rect 3476 6060 3482 6112
rect 3970 6060 3976 6112
rect 4028 6100 4034 6112
rect 4080 6109 4108 6208
rect 4798 6196 4804 6208
rect 4856 6236 4862 6248
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 4856 6208 6377 6236
rect 4856 6196 4862 6208
rect 6365 6205 6377 6208
rect 6411 6205 6423 6239
rect 6365 6199 6423 6205
rect 6641 6239 6699 6245
rect 6641 6205 6653 6239
rect 6687 6236 6699 6239
rect 7006 6236 7012 6248
rect 6687 6208 7012 6236
rect 6687 6205 6699 6208
rect 6641 6199 6699 6205
rect 7006 6196 7012 6208
rect 7064 6196 7070 6248
rect 7650 6196 7656 6248
rect 7708 6236 7714 6248
rect 7708 6208 9076 6236
rect 7708 6196 7714 6208
rect 9048 6180 9076 6208
rect 9490 6196 9496 6248
rect 9548 6236 9554 6248
rect 9674 6236 9680 6248
rect 9548 6208 9680 6236
rect 9548 6196 9554 6208
rect 9674 6196 9680 6208
rect 9732 6196 9738 6248
rect 10597 6239 10655 6245
rect 10597 6205 10609 6239
rect 10643 6205 10655 6239
rect 10597 6199 10655 6205
rect 8938 6168 8944 6180
rect 8899 6140 8944 6168
rect 8938 6128 8944 6140
rect 8996 6128 9002 6180
rect 9030 6128 9036 6180
rect 9088 6168 9094 6180
rect 9508 6168 9536 6196
rect 10612 6168 10640 6199
rect 9088 6140 9536 6168
rect 9876 6140 10640 6168
rect 9088 6128 9094 6140
rect 4065 6103 4123 6109
rect 4065 6100 4077 6103
rect 4028 6072 4077 6100
rect 4028 6060 4034 6072
rect 4065 6069 4077 6072
rect 4111 6069 4123 6103
rect 5166 6100 5172 6112
rect 5127 6072 5172 6100
rect 4065 6063 4123 6069
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 8481 6103 8539 6109
rect 8481 6069 8493 6103
rect 8527 6100 8539 6103
rect 8846 6100 8852 6112
rect 8527 6072 8852 6100
rect 8527 6069 8539 6072
rect 8481 6063 8539 6069
rect 8846 6060 8852 6072
rect 8904 6060 8910 6112
rect 9677 6103 9735 6109
rect 9677 6069 9689 6103
rect 9723 6100 9735 6103
rect 9876 6100 9904 6140
rect 10042 6100 10048 6112
rect 9723 6072 9904 6100
rect 10003 6072 10048 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 10042 6060 10048 6072
rect 10100 6060 10106 6112
rect 11146 6100 11152 6112
rect 11107 6072 11152 6100
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 11348 6100 11376 6267
rect 11698 6236 11704 6248
rect 11659 6208 11704 6236
rect 11698 6196 11704 6208
rect 11756 6196 11762 6248
rect 12618 6100 12624 6112
rect 11348 6072 12624 6100
rect 12618 6060 12624 6072
rect 12676 6060 12682 6112
rect 1104 6010 13892 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 12214 6010
rect 12266 5958 12278 6010
rect 12330 5958 12342 6010
rect 12394 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 13892 6010
rect 1104 5936 13892 5958
rect 2958 5856 2964 5908
rect 3016 5896 3022 5908
rect 3602 5896 3608 5908
rect 3016 5868 3608 5896
rect 3016 5856 3022 5868
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 7650 5896 7656 5908
rect 7611 5868 7656 5896
rect 7650 5856 7656 5868
rect 7708 5856 7714 5908
rect 8662 5896 8668 5908
rect 8623 5868 8668 5896
rect 8662 5856 8668 5868
rect 8720 5896 8726 5908
rect 8720 5868 9444 5896
rect 8720 5856 8726 5868
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5828 2835 5831
rect 7929 5831 7987 5837
rect 2823 5800 4016 5828
rect 2823 5797 2835 5800
rect 2777 5791 2835 5797
rect 2225 5763 2283 5769
rect 2225 5760 2237 5763
rect 1688 5732 2237 5760
rect 1688 5704 1716 5732
rect 2225 5729 2237 5732
rect 2271 5729 2283 5763
rect 3145 5763 3203 5769
rect 3145 5760 3157 5763
rect 2225 5723 2283 5729
rect 2424 5732 3157 5760
rect 1670 5692 1676 5704
rect 1631 5664 1676 5692
rect 1670 5652 1676 5664
rect 1728 5652 1734 5704
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 1581 5627 1639 5633
rect 1581 5593 1593 5627
rect 1627 5593 1639 5627
rect 1581 5587 1639 5593
rect 1596 5556 1624 5587
rect 1964 5568 1992 5655
rect 2038 5652 2044 5704
rect 2096 5692 2102 5704
rect 2424 5692 2452 5732
rect 3145 5729 3157 5732
rect 3191 5729 3203 5763
rect 3988 5760 4016 5800
rect 7929 5797 7941 5831
rect 7975 5828 7987 5831
rect 7975 5800 9352 5828
rect 7975 5797 7987 5800
rect 7929 5791 7987 5797
rect 7190 5760 7196 5772
rect 3988 5732 7196 5760
rect 3145 5723 3203 5729
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 7834 5720 7840 5772
rect 7892 5760 7898 5772
rect 8113 5763 8171 5769
rect 8113 5760 8125 5763
rect 7892 5732 8125 5760
rect 7892 5720 7898 5732
rect 8113 5729 8125 5732
rect 8159 5729 8171 5763
rect 8113 5723 8171 5729
rect 8205 5763 8263 5769
rect 8205 5729 8217 5763
rect 8251 5760 8263 5763
rect 8570 5760 8576 5772
rect 8251 5732 8576 5760
rect 8251 5729 8263 5732
rect 8205 5723 8263 5729
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 8846 5720 8852 5772
rect 8904 5760 8910 5772
rect 8904 5732 9076 5760
rect 8904 5720 8910 5732
rect 2096 5664 2452 5692
rect 2501 5695 2559 5701
rect 2096 5652 2102 5664
rect 2501 5661 2513 5695
rect 2547 5661 2559 5695
rect 2501 5655 2559 5661
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5692 2927 5695
rect 2958 5692 2964 5704
rect 2915 5664 2964 5692
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 1670 5556 1676 5568
rect 1596 5528 1676 5556
rect 1670 5516 1676 5528
rect 1728 5516 1734 5568
rect 1946 5556 1952 5568
rect 1859 5528 1952 5556
rect 1946 5516 1952 5528
rect 2004 5556 2010 5568
rect 2516 5556 2544 5655
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 3050 5652 3056 5704
rect 3108 5692 3114 5704
rect 3881 5695 3939 5701
rect 3108 5664 3153 5692
rect 3108 5652 3114 5664
rect 3881 5661 3893 5695
rect 3927 5661 3939 5695
rect 3881 5655 3939 5661
rect 3326 5624 3332 5636
rect 3287 5596 3332 5624
rect 3326 5584 3332 5596
rect 3384 5584 3390 5636
rect 3510 5624 3516 5636
rect 3471 5596 3516 5624
rect 3510 5584 3516 5596
rect 3568 5584 3574 5636
rect 3896 5624 3924 5655
rect 7466 5652 7472 5704
rect 7524 5692 7530 5704
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 7524 5664 7573 5692
rect 7524 5652 7530 5664
rect 7561 5661 7573 5664
rect 7607 5661 7619 5695
rect 7561 5655 7619 5661
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 4154 5624 4160 5636
rect 3896 5596 4016 5624
rect 4115 5596 4160 5624
rect 3988 5568 4016 5596
rect 4154 5584 4160 5596
rect 4212 5584 4218 5636
rect 5166 5584 5172 5636
rect 5224 5584 5230 5636
rect 2004 5528 2544 5556
rect 2004 5516 2010 5528
rect 2958 5516 2964 5568
rect 3016 5556 3022 5568
rect 3878 5556 3884 5568
rect 3016 5528 3884 5556
rect 3016 5516 3022 5528
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 3970 5516 3976 5568
rect 4028 5516 4034 5568
rect 5074 5516 5080 5568
rect 5132 5556 5138 5568
rect 5629 5559 5687 5565
rect 5629 5556 5641 5559
rect 5132 5528 5641 5556
rect 5132 5516 5138 5528
rect 5629 5525 5641 5528
rect 5675 5525 5687 5559
rect 7576 5556 7604 5655
rect 8036 5624 8064 5655
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 8389 5695 8447 5701
rect 8389 5692 8401 5695
rect 8352 5664 8401 5692
rect 8352 5652 8358 5664
rect 8389 5661 8401 5664
rect 8435 5661 8447 5695
rect 8389 5655 8447 5661
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 8754 5692 8760 5704
rect 8527 5664 8760 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 8754 5652 8760 5664
rect 8812 5652 8818 5704
rect 8938 5692 8944 5704
rect 8899 5664 8944 5692
rect 8938 5652 8944 5664
rect 8996 5652 9002 5704
rect 9048 5701 9076 5732
rect 9034 5695 9092 5701
rect 9034 5661 9046 5695
rect 9080 5661 9092 5695
rect 9214 5692 9220 5704
rect 9175 5664 9220 5692
rect 9034 5655 9092 5661
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 9324 5701 9352 5800
rect 9416 5701 9444 5868
rect 10410 5856 10416 5908
rect 10468 5896 10474 5908
rect 11517 5899 11575 5905
rect 11517 5896 11529 5899
rect 10468 5868 11529 5896
rect 10468 5856 10474 5868
rect 11517 5865 11529 5868
rect 11563 5865 11575 5899
rect 11517 5859 11575 5865
rect 13354 5856 13360 5908
rect 13412 5896 13418 5908
rect 13449 5899 13507 5905
rect 13449 5896 13461 5899
rect 13412 5868 13461 5896
rect 13412 5856 13418 5868
rect 13449 5865 13461 5868
rect 13495 5865 13507 5899
rect 13449 5859 13507 5865
rect 10042 5760 10048 5772
rect 10003 5732 10048 5760
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 9309 5695 9367 5701
rect 9309 5661 9321 5695
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 9406 5695 9464 5701
rect 9406 5661 9418 5695
rect 9452 5661 9464 5695
rect 9406 5655 9464 5661
rect 9769 5695 9827 5701
rect 9769 5661 9781 5695
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 9232 5624 9260 5652
rect 8036 5596 9260 5624
rect 8938 5556 8944 5568
rect 7576 5528 8944 5556
rect 5629 5519 5687 5525
rect 8938 5516 8944 5528
rect 8996 5516 9002 5568
rect 9582 5556 9588 5568
rect 9543 5528 9588 5556
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 9784 5556 9812 5655
rect 11146 5652 11152 5704
rect 11204 5652 11210 5704
rect 11698 5692 11704 5704
rect 11611 5664 11704 5692
rect 11698 5652 11704 5664
rect 11756 5652 11762 5704
rect 11514 5556 11520 5568
rect 9784 5528 11520 5556
rect 11514 5516 11520 5528
rect 11572 5556 11578 5568
rect 11716 5556 11744 5652
rect 11974 5624 11980 5636
rect 11935 5596 11980 5624
rect 11974 5584 11980 5596
rect 12032 5584 12038 5636
rect 12710 5584 12716 5636
rect 12768 5584 12774 5636
rect 11572 5528 11744 5556
rect 11572 5516 11578 5528
rect 1104 5466 13892 5488
rect 1104 5414 8214 5466
rect 8266 5414 8278 5466
rect 8330 5414 8342 5466
rect 8394 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 13892 5466
rect 1104 5392 13892 5414
rect 1946 5352 1952 5364
rect 1907 5324 1952 5352
rect 1946 5312 1952 5324
rect 2004 5312 2010 5364
rect 3602 5312 3608 5364
rect 3660 5312 3666 5364
rect 4154 5352 4160 5364
rect 4115 5324 4160 5352
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 5626 5352 5632 5364
rect 4540 5324 5632 5352
rect 2958 5284 2964 5296
rect 2919 5256 2964 5284
rect 2958 5244 2964 5256
rect 3016 5244 3022 5296
rect 3620 5284 3648 5312
rect 3252 5256 3648 5284
rect 1394 5216 1400 5228
rect 1355 5188 1400 5216
rect 1394 5176 1400 5188
rect 1452 5176 1458 5228
rect 1578 5216 1584 5228
rect 1539 5188 1584 5216
rect 1578 5176 1584 5188
rect 1636 5176 1642 5228
rect 2038 5176 2044 5228
rect 2096 5216 2102 5228
rect 2864 5219 2922 5225
rect 2096 5188 2141 5216
rect 2096 5176 2102 5188
rect 2864 5185 2876 5219
rect 2910 5185 2922 5219
rect 2864 5179 2922 5185
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5117 2467 5151
rect 2409 5111 2467 5117
rect 2501 5151 2559 5157
rect 2501 5117 2513 5151
rect 2547 5148 2559 5151
rect 2774 5148 2780 5160
rect 2547 5120 2780 5148
rect 2547 5117 2559 5120
rect 2501 5111 2559 5117
rect 2424 5080 2452 5111
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 2879 5148 2907 5179
rect 3050 5176 3056 5228
rect 3108 5216 3114 5228
rect 3252 5225 3280 5256
rect 3602 5225 3608 5228
rect 3237 5219 3295 5225
rect 3108 5188 3153 5216
rect 3108 5176 3114 5188
rect 3237 5185 3249 5219
rect 3283 5185 3295 5219
rect 3600 5216 3608 5225
rect 3563 5188 3608 5216
rect 3237 5179 3295 5185
rect 3600 5179 3608 5188
rect 3602 5176 3608 5179
rect 3660 5176 3666 5228
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5185 3755 5219
rect 3697 5179 3755 5185
rect 3789 5219 3847 5225
rect 3789 5185 3801 5219
rect 3835 5216 3847 5219
rect 3878 5216 3884 5228
rect 3835 5188 3884 5216
rect 3835 5185 3847 5188
rect 3789 5179 3847 5185
rect 3418 5148 3424 5160
rect 2879 5120 3424 5148
rect 3418 5108 3424 5120
rect 3476 5148 3482 5160
rect 3712 5148 3740 5179
rect 3878 5176 3884 5188
rect 3936 5176 3942 5228
rect 3973 5219 4031 5225
rect 3973 5185 3985 5219
rect 4019 5185 4031 5219
rect 4430 5216 4436 5228
rect 4391 5188 4436 5216
rect 3973 5179 4031 5185
rect 3476 5120 3740 5148
rect 3476 5108 3482 5120
rect 2685 5083 2743 5089
rect 2685 5080 2697 5083
rect 2424 5052 2697 5080
rect 2685 5049 2697 5052
rect 2731 5080 2743 5083
rect 3326 5080 3332 5092
rect 2731 5052 3332 5080
rect 2731 5049 2743 5052
rect 2685 5043 2743 5049
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 3896 5080 3924 5176
rect 3988 5148 4016 5179
rect 4430 5176 4436 5188
rect 4488 5176 4494 5228
rect 4062 5148 4068 5160
rect 3975 5120 4068 5148
rect 4062 5108 4068 5120
rect 4120 5148 4126 5160
rect 4540 5148 4568 5324
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 6457 5355 6515 5361
rect 6457 5321 6469 5355
rect 6503 5321 6515 5355
rect 11974 5352 11980 5364
rect 6457 5315 6515 5321
rect 9232 5324 11980 5352
rect 5442 5284 5448 5296
rect 5000 5256 5448 5284
rect 5000 5225 5028 5256
rect 5442 5244 5448 5256
rect 5500 5244 5506 5296
rect 6472 5284 6500 5315
rect 9232 5293 9260 5324
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 12710 5352 12716 5364
rect 12671 5324 12716 5352
rect 12710 5312 12716 5324
rect 12768 5312 12774 5364
rect 9217 5287 9275 5293
rect 5552 5256 6500 5284
rect 8312 5256 9076 5284
rect 5552 5228 5580 5256
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5185 5043 5219
rect 5166 5216 5172 5228
rect 5127 5188 5172 5216
rect 4985 5179 5043 5185
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 5534 5216 5540 5228
rect 5495 5188 5540 5216
rect 5534 5176 5540 5188
rect 5592 5176 5598 5228
rect 6012 5225 6040 5256
rect 8312 5228 8340 5256
rect 5813 5219 5871 5225
rect 5813 5216 5825 5219
rect 5644 5188 5825 5216
rect 4120 5120 4568 5148
rect 4617 5151 4675 5157
rect 4120 5108 4126 5120
rect 4617 5117 4629 5151
rect 4663 5148 4675 5151
rect 5261 5151 5319 5157
rect 5261 5148 5273 5151
rect 4663 5120 5273 5148
rect 4663 5117 4675 5120
rect 4617 5111 4675 5117
rect 5261 5117 5273 5120
rect 5307 5117 5319 5151
rect 5261 5111 5319 5117
rect 5166 5080 5172 5092
rect 3896 5052 5172 5080
rect 5166 5040 5172 5052
rect 5224 5040 5230 5092
rect 5276 5080 5304 5111
rect 5350 5108 5356 5160
rect 5408 5148 5414 5160
rect 5644 5148 5672 5188
rect 5813 5185 5825 5188
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 5997 5219 6055 5225
rect 5997 5185 6009 5219
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 6822 5176 6828 5228
rect 6880 5176 6886 5228
rect 8294 5216 8300 5228
rect 8255 5188 8300 5216
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 8754 5216 8760 5228
rect 8715 5188 8760 5216
rect 8754 5176 8760 5188
rect 8812 5176 8818 5228
rect 8938 5216 8944 5228
rect 8899 5188 8944 5216
rect 8938 5176 8944 5188
rect 8996 5176 9002 5228
rect 9048 5216 9076 5256
rect 9217 5253 9229 5287
rect 9263 5253 9275 5287
rect 9217 5247 9275 5253
rect 9309 5287 9367 5293
rect 9309 5253 9321 5287
rect 9355 5284 9367 5287
rect 9582 5284 9588 5296
rect 9355 5256 9588 5284
rect 9355 5253 9367 5256
rect 9309 5247 9367 5253
rect 9582 5244 9588 5256
rect 9640 5244 9646 5296
rect 10410 5284 10416 5296
rect 10060 5256 10416 5284
rect 9398 5216 9404 5228
rect 9048 5188 9404 5216
rect 9398 5176 9404 5188
rect 9456 5216 9462 5228
rect 10060 5216 10088 5256
rect 10410 5244 10416 5256
rect 10468 5244 10474 5296
rect 10778 5284 10784 5296
rect 10739 5256 10784 5284
rect 10778 5244 10784 5256
rect 10836 5244 10842 5296
rect 10870 5244 10876 5296
rect 10928 5284 10934 5296
rect 10928 5256 11744 5284
rect 10928 5244 10934 5256
rect 9456 5188 10088 5216
rect 9456 5176 9462 5188
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 10505 5219 10563 5225
rect 10505 5216 10517 5219
rect 10192 5188 10517 5216
rect 10192 5176 10198 5188
rect 10505 5185 10517 5188
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5216 10655 5219
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10643 5188 10977 5216
rect 10643 5185 10655 5188
rect 10597 5179 10655 5185
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 10965 5179 11023 5185
rect 11057 5219 11115 5225
rect 11057 5185 11069 5219
rect 11103 5216 11115 5219
rect 11606 5216 11612 5228
rect 11103 5188 11612 5216
rect 11103 5185 11115 5188
rect 11057 5179 11115 5185
rect 11606 5176 11612 5188
rect 11664 5176 11670 5228
rect 11716 5225 11744 5256
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 12529 5219 12587 5225
rect 12529 5185 12541 5219
rect 12575 5216 12587 5219
rect 12618 5216 12624 5228
rect 12575 5188 12624 5216
rect 12575 5185 12587 5188
rect 12529 5179 12587 5185
rect 12618 5176 12624 5188
rect 12676 5176 12682 5228
rect 5408 5120 5672 5148
rect 5721 5151 5779 5157
rect 5408 5108 5414 5120
rect 5721 5117 5733 5151
rect 5767 5148 5779 5151
rect 7929 5151 7987 5157
rect 7929 5148 7941 5151
rect 5767 5120 7941 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 7929 5117 7941 5120
rect 7975 5117 7987 5151
rect 8205 5151 8263 5157
rect 8205 5148 8217 5151
rect 7929 5111 7987 5117
rect 8128 5120 8217 5148
rect 5905 5083 5963 5089
rect 5905 5080 5917 5083
rect 5276 5052 5917 5080
rect 5905 5049 5917 5052
rect 5951 5049 5963 5083
rect 5905 5043 5963 5049
rect 1673 5015 1731 5021
rect 1673 4981 1685 5015
rect 1719 5012 1731 5015
rect 2406 5012 2412 5024
rect 1719 4984 2412 5012
rect 1719 4981 1731 4984
rect 1673 4975 1731 4981
rect 2406 4972 2412 4984
rect 2464 4972 2470 5024
rect 3234 4972 3240 5024
rect 3292 5012 3298 5024
rect 3421 5015 3479 5021
rect 3421 5012 3433 5015
rect 3292 4984 3433 5012
rect 3292 4972 3298 4984
rect 3421 4981 3433 4984
rect 3467 4981 3479 5015
rect 3421 4975 3479 4981
rect 3602 4972 3608 5024
rect 3660 5012 3666 5024
rect 5442 5012 5448 5024
rect 3660 4984 5448 5012
rect 3660 4972 3666 4984
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 8128 5012 8156 5120
rect 8205 5117 8217 5120
rect 8251 5117 8263 5151
rect 8772 5148 8800 5176
rect 9858 5148 9864 5160
rect 8772 5120 9864 5148
rect 8205 5111 8263 5117
rect 9858 5108 9864 5120
rect 9916 5108 9922 5160
rect 10413 5151 10471 5157
rect 10413 5117 10425 5151
rect 10459 5148 10471 5151
rect 10686 5148 10692 5160
rect 10459 5120 10692 5148
rect 10459 5117 10471 5120
rect 10413 5111 10471 5117
rect 10686 5108 10692 5120
rect 10744 5148 10750 5160
rect 11333 5151 11391 5157
rect 11333 5148 11345 5151
rect 10744 5120 11345 5148
rect 10744 5108 10750 5120
rect 11333 5117 11345 5120
rect 11379 5117 11391 5151
rect 11333 5111 11391 5117
rect 9214 5040 9220 5092
rect 9272 5080 9278 5092
rect 10597 5083 10655 5089
rect 10597 5080 10609 5083
rect 9272 5052 10609 5080
rect 9272 5040 9278 5052
rect 8386 5012 8392 5024
rect 7524 4984 8156 5012
rect 8347 4984 8392 5012
rect 7524 4972 7530 4984
rect 8386 4972 8392 4984
rect 8444 4972 8450 5024
rect 10042 4972 10048 5024
rect 10100 5012 10106 5024
rect 10336 5021 10364 5052
rect 10597 5049 10609 5052
rect 10643 5049 10655 5083
rect 11348 5080 11376 5111
rect 11609 5083 11667 5089
rect 11609 5080 11621 5083
rect 11348 5052 11621 5080
rect 10597 5043 10655 5049
rect 11609 5049 11621 5052
rect 11655 5049 11667 5083
rect 11609 5043 11667 5049
rect 10137 5015 10195 5021
rect 10137 5012 10149 5015
rect 10100 4984 10149 5012
rect 10100 4972 10106 4984
rect 10137 4981 10149 4984
rect 10183 4981 10195 5015
rect 10137 4975 10195 4981
rect 10321 5015 10379 5021
rect 10321 4981 10333 5015
rect 10367 4981 10379 5015
rect 10321 4975 10379 4981
rect 10410 4972 10416 5024
rect 10468 5012 10474 5024
rect 11241 5015 11299 5021
rect 11241 5012 11253 5015
rect 10468 4984 11253 5012
rect 10468 4972 10474 4984
rect 11241 4981 11253 4984
rect 11287 4981 11299 5015
rect 11241 4975 11299 4981
rect 1104 4922 13892 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 12214 4922
rect 12266 4870 12278 4922
rect 12330 4870 12342 4922
rect 12394 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 13892 4922
rect 1104 4848 13892 4870
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3510 4808 3516 4820
rect 2832 4780 3516 4808
rect 2832 4768 2838 4780
rect 3510 4768 3516 4780
rect 3568 4808 3574 4820
rect 4433 4811 4491 4817
rect 4433 4808 4445 4811
rect 3568 4780 4445 4808
rect 3568 4768 3574 4780
rect 4433 4777 4445 4780
rect 4479 4777 4491 4811
rect 4433 4771 4491 4777
rect 4890 4768 4896 4820
rect 4948 4808 4954 4820
rect 5902 4808 5908 4820
rect 4948 4780 5908 4808
rect 4948 4768 4954 4780
rect 5902 4768 5908 4780
rect 5960 4768 5966 4820
rect 6733 4811 6791 4817
rect 6733 4777 6745 4811
rect 6779 4808 6791 4811
rect 6822 4808 6828 4820
rect 6779 4780 6828 4808
rect 6779 4777 6791 4780
rect 6733 4771 6791 4777
rect 6822 4768 6828 4780
rect 6880 4768 6886 4820
rect 8938 4768 8944 4820
rect 8996 4808 9002 4820
rect 9398 4808 9404 4820
rect 8996 4780 9404 4808
rect 8996 4768 9002 4780
rect 9398 4768 9404 4780
rect 9456 4808 9462 4820
rect 9677 4811 9735 4817
rect 9677 4808 9689 4811
rect 9456 4780 9689 4808
rect 9456 4768 9462 4780
rect 9677 4777 9689 4780
rect 9723 4808 9735 4811
rect 10226 4808 10232 4820
rect 9723 4780 10232 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 10226 4768 10232 4780
rect 10284 4808 10290 4820
rect 10284 4780 10916 4808
rect 10284 4768 10290 4780
rect 1394 4700 1400 4752
rect 1452 4740 1458 4752
rect 2869 4743 2927 4749
rect 2869 4740 2881 4743
rect 1452 4712 2881 4740
rect 1452 4700 1458 4712
rect 1504 4613 1532 4712
rect 2869 4709 2881 4712
rect 2915 4709 2927 4743
rect 2869 4703 2927 4709
rect 3881 4743 3939 4749
rect 3881 4709 3893 4743
rect 3927 4740 3939 4743
rect 4706 4740 4712 4752
rect 3927 4712 4712 4740
rect 3927 4709 3939 4712
rect 3881 4703 3939 4709
rect 2314 4672 2320 4684
rect 2275 4644 2320 4672
rect 2314 4632 2320 4644
rect 2372 4632 2378 4684
rect 3033 4675 3091 4681
rect 3033 4641 3045 4675
rect 3079 4672 3091 4675
rect 3510 4672 3516 4684
rect 3079 4644 3516 4672
rect 3079 4641 3091 4644
rect 3033 4635 3091 4641
rect 3510 4632 3516 4644
rect 3568 4632 3574 4684
rect 3896 4672 3924 4703
rect 4706 4700 4712 4712
rect 4764 4700 4770 4752
rect 5166 4740 5172 4752
rect 5079 4712 5172 4740
rect 5166 4700 5172 4712
rect 5224 4740 5230 4752
rect 5994 4740 6000 4752
rect 5224 4712 6000 4740
rect 5224 4700 5230 4712
rect 5994 4700 6000 4712
rect 6052 4700 6058 4752
rect 7561 4743 7619 4749
rect 7561 4709 7573 4743
rect 7607 4740 7619 4743
rect 8294 4740 8300 4752
rect 7607 4712 8300 4740
rect 7607 4709 7619 4712
rect 7561 4703 7619 4709
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 10042 4740 10048 4752
rect 10003 4712 10048 4740
rect 10042 4700 10048 4712
rect 10100 4700 10106 4752
rect 3620 4644 3924 4672
rect 1489 4607 1547 4613
rect 1489 4573 1501 4607
rect 1535 4573 1547 4607
rect 1489 4567 1547 4573
rect 1578 4564 1584 4616
rect 1636 4604 1642 4616
rect 1765 4607 1823 4613
rect 1765 4604 1777 4607
rect 1636 4576 1777 4604
rect 1636 4564 1642 4576
rect 1765 4573 1777 4576
rect 1811 4573 1823 4607
rect 1765 4567 1823 4573
rect 1854 4564 1860 4616
rect 1912 4604 1918 4616
rect 2041 4607 2099 4613
rect 2041 4604 2053 4607
rect 1912 4576 2053 4604
rect 1912 4564 1918 4576
rect 2041 4573 2053 4576
rect 2087 4573 2099 4607
rect 2041 4567 2099 4573
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4573 2283 4607
rect 2406 4604 2412 4616
rect 2367 4576 2412 4604
rect 2225 4567 2283 4573
rect 2240 4536 2268 4567
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 3145 4607 3203 4613
rect 3145 4573 3157 4607
rect 3191 4604 3203 4607
rect 3421 4607 3479 4613
rect 3421 4604 3433 4607
rect 3191 4576 3433 4604
rect 3191 4573 3203 4576
rect 3145 4567 3203 4573
rect 3421 4573 3433 4576
rect 3467 4604 3479 4607
rect 3620 4604 3648 4644
rect 3970 4632 3976 4684
rect 4028 4672 4034 4684
rect 4338 4672 4344 4684
rect 4028 4644 4344 4672
rect 4028 4632 4034 4644
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 3786 4604 3792 4616
rect 3467 4576 3648 4604
rect 3747 4576 3792 4604
rect 3467 4573 3479 4576
rect 3421 4567 3479 4573
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 3878 4564 3884 4616
rect 3936 4604 3942 4616
rect 5184 4613 5212 4700
rect 5810 4672 5816 4684
rect 5460 4644 5816 4672
rect 5460 4613 5488 4644
rect 5810 4632 5816 4644
rect 5868 4672 5874 4684
rect 6365 4675 6423 4681
rect 6365 4672 6377 4675
rect 5868 4644 6377 4672
rect 5868 4632 5874 4644
rect 6365 4641 6377 4644
rect 6411 4641 6423 4675
rect 6365 4635 6423 4641
rect 8386 4632 8392 4684
rect 8444 4672 8450 4684
rect 10778 4672 10784 4684
rect 8444 4644 10784 4672
rect 8444 4632 8450 4644
rect 4251 4607 4309 4613
rect 4251 4604 4263 4607
rect 3936 4576 4263 4604
rect 3936 4564 3942 4576
rect 4251 4573 4263 4576
rect 4297 4604 4309 4607
rect 5169 4607 5227 4613
rect 4297 4576 4844 4604
rect 4297 4573 4309 4576
rect 4251 4567 4309 4573
rect 2958 4536 2964 4548
rect 2240 4508 2964 4536
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 4816 4536 4844 4576
rect 5169 4573 5181 4607
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 5626 4564 5632 4616
rect 5684 4604 5690 4616
rect 5902 4604 5908 4616
rect 5684 4576 5777 4604
rect 5863 4576 5908 4604
rect 5684 4564 5690 4576
rect 5902 4564 5908 4576
rect 5960 4604 5966 4616
rect 6270 4604 6276 4616
rect 5960 4576 6276 4604
rect 5960 4564 5966 4576
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 6457 4607 6515 4613
rect 6457 4573 6469 4607
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 5258 4536 5264 4548
rect 4816 4508 5120 4536
rect 5219 4508 5264 4536
rect 2130 4428 2136 4480
rect 2188 4468 2194 4480
rect 2501 4471 2559 4477
rect 2501 4468 2513 4471
rect 2188 4440 2513 4468
rect 2188 4428 2194 4440
rect 2501 4437 2513 4440
rect 2547 4437 2559 4471
rect 2501 4431 2559 4437
rect 3970 4428 3976 4480
rect 4028 4468 4034 4480
rect 4249 4471 4307 4477
rect 4249 4468 4261 4471
rect 4028 4440 4261 4468
rect 4028 4428 4034 4440
rect 4249 4437 4261 4440
rect 4295 4437 4307 4471
rect 4249 4431 4307 4437
rect 4614 4428 4620 4480
rect 4672 4468 4678 4480
rect 4985 4471 5043 4477
rect 4985 4468 4997 4471
rect 4672 4440 4997 4468
rect 4672 4428 4678 4440
rect 4985 4437 4997 4440
rect 5031 4437 5043 4471
rect 5092 4468 5120 4508
rect 5258 4496 5264 4508
rect 5316 4496 5322 4548
rect 5353 4539 5411 4545
rect 5353 4505 5365 4539
rect 5399 4505 5411 4539
rect 5644 4536 5672 4564
rect 6472 4536 6500 4567
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 7190 4604 7196 4616
rect 6604 4576 6649 4604
rect 7151 4576 7196 4604
rect 6604 4564 6610 4576
rect 7190 4564 7196 4576
rect 7248 4604 7254 4616
rect 8110 4604 8116 4616
rect 7248 4576 8116 4604
rect 7248 4564 7254 4576
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4573 9183 4607
rect 9490 4604 9496 4616
rect 9451 4576 9496 4604
rect 9125 4567 9183 4573
rect 6638 4536 6644 4548
rect 5644 4508 5856 4536
rect 6472 4508 6644 4536
rect 5353 4499 5411 4505
rect 5368 4468 5396 4499
rect 5534 4468 5540 4480
rect 5092 4440 5540 4468
rect 4985 4431 5043 4437
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 5626 4428 5632 4480
rect 5684 4468 5690 4480
rect 5721 4471 5779 4477
rect 5721 4468 5733 4471
rect 5684 4440 5733 4468
rect 5684 4428 5690 4440
rect 5721 4437 5733 4440
rect 5767 4437 5779 4471
rect 5828 4468 5856 4508
rect 6638 4496 6644 4508
rect 6696 4496 6702 4548
rect 7374 4536 7380 4548
rect 7335 4508 7380 4536
rect 7374 4496 7380 4508
rect 7432 4496 7438 4548
rect 8754 4536 8760 4548
rect 7576 4508 8760 4536
rect 7576 4480 7604 4508
rect 8754 4496 8760 4508
rect 8812 4536 8818 4548
rect 9140 4536 9168 4567
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 9858 4604 9864 4616
rect 9819 4576 9864 4604
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 9968 4613 9996 4644
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 9953 4607 10011 4613
rect 9953 4573 9965 4607
rect 9999 4573 10011 4607
rect 10134 4604 10140 4616
rect 10095 4576 10140 4604
rect 9953 4567 10011 4573
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 10686 4604 10692 4616
rect 10647 4576 10692 4604
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 10888 4613 10916 4780
rect 12161 4743 12219 4749
rect 12161 4740 12173 4743
rect 10980 4712 12173 4740
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4573 10931 4607
rect 10980 4604 11008 4712
rect 12161 4709 12173 4712
rect 12207 4709 12219 4743
rect 12161 4703 12219 4709
rect 11057 4675 11115 4681
rect 11057 4641 11069 4675
rect 11103 4672 11115 4675
rect 11790 4672 11796 4684
rect 11103 4644 11796 4672
rect 11103 4641 11115 4644
rect 11057 4635 11115 4641
rect 11790 4632 11796 4644
rect 11848 4632 11854 4684
rect 11149 4607 11207 4613
rect 11149 4604 11161 4607
rect 10980 4576 11161 4604
rect 10873 4567 10931 4573
rect 11149 4573 11161 4576
rect 11195 4573 11207 4607
rect 11149 4567 11207 4573
rect 11333 4607 11391 4613
rect 11333 4573 11345 4607
rect 11379 4573 11391 4607
rect 11606 4604 11612 4616
rect 11567 4576 11612 4604
rect 11333 4567 11391 4573
rect 11054 4536 11060 4548
rect 8812 4508 9168 4536
rect 9416 4508 11060 4536
rect 8812 4496 8818 4508
rect 6454 4468 6460 4480
rect 5828 4440 6460 4468
rect 5721 4431 5779 4437
rect 6454 4428 6460 4440
rect 6512 4428 6518 4480
rect 6546 4428 6552 4480
rect 6604 4468 6610 4480
rect 7558 4468 7564 4480
rect 6604 4440 7564 4468
rect 6604 4428 6610 4440
rect 7558 4428 7564 4440
rect 7616 4428 7622 4480
rect 8846 4428 8852 4480
rect 8904 4468 8910 4480
rect 8941 4471 8999 4477
rect 8941 4468 8953 4471
rect 8904 4440 8953 4468
rect 8904 4428 8910 4440
rect 8941 4437 8953 4440
rect 8987 4437 8999 4471
rect 8941 4431 8999 4437
rect 9214 4428 9220 4480
rect 9272 4468 9278 4480
rect 9416 4477 9444 4508
rect 11054 4496 11060 4508
rect 11112 4496 11118 4548
rect 9401 4471 9459 4477
rect 9401 4468 9413 4471
rect 9272 4440 9413 4468
rect 9272 4428 9278 4440
rect 9401 4437 9413 4440
rect 9447 4437 9459 4471
rect 9401 4431 9459 4437
rect 9582 4428 9588 4480
rect 9640 4468 9646 4480
rect 11348 4468 11376 4567
rect 11606 4564 11612 4576
rect 11664 4604 11670 4616
rect 11885 4607 11943 4613
rect 11885 4604 11897 4607
rect 11664 4576 11897 4604
rect 11664 4564 11670 4576
rect 11885 4573 11897 4576
rect 11931 4573 11943 4607
rect 11885 4567 11943 4573
rect 11997 4607 12055 4613
rect 11997 4573 12009 4607
rect 12043 4573 12055 4607
rect 11997 4567 12055 4573
rect 11422 4496 11428 4548
rect 11480 4536 11486 4548
rect 11517 4539 11575 4545
rect 11517 4536 11529 4539
rect 11480 4508 11529 4536
rect 11480 4496 11486 4508
rect 11517 4505 11529 4508
rect 11563 4536 11575 4539
rect 12012 4536 12040 4567
rect 11563 4508 12040 4536
rect 11563 4505 11575 4508
rect 11517 4499 11575 4505
rect 9640 4440 11376 4468
rect 9640 4428 9646 4440
rect 1104 4378 13892 4400
rect 1104 4326 8214 4378
rect 8266 4326 8278 4378
rect 8330 4326 8342 4378
rect 8394 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 13892 4378
rect 1104 4304 13892 4326
rect 3878 4264 3884 4276
rect 3068 4236 3884 4264
rect 3068 4140 3096 4236
rect 3878 4224 3884 4236
rect 3936 4224 3942 4276
rect 7374 4264 7380 4276
rect 6380 4236 7380 4264
rect 3510 4196 3516 4208
rect 3471 4168 3516 4196
rect 3510 4156 3516 4168
rect 3568 4156 3574 4208
rect 3970 4196 3976 4208
rect 3931 4168 3976 4196
rect 3970 4156 3976 4168
rect 4028 4156 4034 4208
rect 4614 4196 4620 4208
rect 4575 4168 4620 4196
rect 4614 4156 4620 4168
rect 4672 4156 4678 4208
rect 5626 4156 5632 4208
rect 5684 4156 5690 4208
rect 1670 4088 1676 4140
rect 1728 4128 1734 4140
rect 1765 4131 1823 4137
rect 1765 4128 1777 4131
rect 1728 4100 1777 4128
rect 1728 4088 1734 4100
rect 1765 4097 1777 4100
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 1948 4131 2006 4137
rect 1948 4097 1960 4131
rect 1994 4097 2006 4131
rect 2130 4128 2136 4140
rect 2091 4100 2136 4128
rect 1948 4091 2006 4097
rect 1964 3924 1992 4091
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2314 4128 2320 4140
rect 2275 4100 2320 4128
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 2590 4128 2596 4140
rect 2551 4100 2596 4128
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 3050 4128 3056 4140
rect 3011 4100 3056 4128
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 3237 4131 3295 4137
rect 3237 4097 3249 4131
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4128 3387 4131
rect 3697 4131 3755 4137
rect 3697 4128 3709 4131
rect 3375 4100 3709 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 3697 4097 3709 4100
rect 3743 4128 3755 4131
rect 3786 4128 3792 4140
rect 3743 4100 3792 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 2038 4020 2044 4072
rect 2096 4060 2102 4072
rect 3252 4060 3280 4091
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 6380 4128 6408 4236
rect 7374 4224 7380 4236
rect 7432 4224 7438 4276
rect 8110 4224 8116 4276
rect 8168 4264 8174 4276
rect 8168 4236 9444 4264
rect 8168 4224 8174 4236
rect 6733 4199 6791 4205
rect 6733 4165 6745 4199
rect 6779 4196 6791 4199
rect 6779 4168 7420 4196
rect 6779 4165 6791 4168
rect 6733 4159 6791 4165
rect 7392 4140 7420 4168
rect 8846 4156 8852 4208
rect 8904 4156 8910 4208
rect 9416 4196 9444 4236
rect 9490 4224 9496 4276
rect 9548 4264 9554 4276
rect 9585 4267 9643 4273
rect 9585 4264 9597 4267
rect 9548 4236 9597 4264
rect 9548 4224 9554 4236
rect 9585 4233 9597 4236
rect 9631 4233 9643 4267
rect 9585 4227 9643 4233
rect 9861 4267 9919 4273
rect 9861 4233 9873 4267
rect 9907 4264 9919 4267
rect 10134 4264 10140 4276
rect 9907 4236 10140 4264
rect 9907 4233 9919 4236
rect 9861 4227 9919 4233
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 10502 4224 10508 4276
rect 10560 4264 10566 4276
rect 9416 4168 9996 4196
rect 5828 4100 6408 4128
rect 3970 4060 3976 4072
rect 2096 4032 2141 4060
rect 3252 4032 3976 4060
rect 2096 4020 2102 4032
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 4338 4060 4344 4072
rect 4299 4032 4344 4060
rect 4338 4020 4344 4032
rect 4396 4020 4402 4072
rect 5828 4060 5856 4100
rect 6454 4088 6460 4140
rect 6512 4128 6518 4140
rect 6512 4100 6557 4128
rect 6512 4088 6518 4100
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 6696 4100 6741 4128
rect 6696 4088 6702 4100
rect 6822 4088 6828 4140
rect 6880 4137 6886 4140
rect 6880 4128 6888 4137
rect 7374 4128 7380 4140
rect 6880 4100 6925 4128
rect 7335 4100 7380 4128
rect 6880 4091 6888 4100
rect 6880 4088 6886 4091
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 7558 4128 7564 4140
rect 7519 4100 7564 4128
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 9968 4137 9996 4168
rect 9953 4131 10011 4137
rect 9953 4097 9965 4131
rect 9999 4097 10011 4131
rect 9953 4091 10011 4097
rect 10318 4088 10324 4140
rect 10376 4128 10382 4140
rect 10560 4137 10588 4264
rect 10686 4224 10692 4276
rect 10744 4264 10750 4276
rect 10744 4236 10916 4264
rect 10744 4224 10750 4236
rect 10888 4205 10916 4236
rect 10873 4199 10931 4205
rect 10873 4165 10885 4199
rect 10919 4165 10931 4199
rect 11790 4196 11796 4208
rect 11751 4168 11796 4196
rect 10873 4159 10931 4165
rect 11790 4156 11796 4168
rect 11848 4156 11854 4208
rect 12802 4156 12808 4208
rect 12860 4156 12866 4208
rect 10517 4131 10588 4137
rect 10376 4100 10439 4128
rect 10376 4088 10382 4100
rect 4448 4032 5856 4060
rect 6656 4032 7420 4060
rect 2501 3995 2559 4001
rect 2501 3961 2513 3995
rect 2547 3992 2559 3995
rect 4448 3992 4476 4032
rect 6656 3992 6684 4032
rect 2547 3964 4476 3992
rect 5644 3964 6684 3992
rect 2547 3961 2559 3964
rect 2501 3955 2559 3961
rect 2685 3927 2743 3933
rect 2685 3924 2697 3927
rect 1964 3896 2697 3924
rect 2685 3893 2697 3896
rect 2731 3893 2743 3927
rect 2685 3887 2743 3893
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 5644 3924 5672 3964
rect 6730 3952 6736 4004
rect 6788 3992 6794 4004
rect 7285 3995 7343 4001
rect 7285 3992 7297 3995
rect 6788 3964 7297 3992
rect 6788 3952 6794 3964
rect 7285 3961 7297 3964
rect 7331 3961 7343 3995
rect 7392 3992 7420 4032
rect 7466 4020 7472 4072
rect 7524 4060 7530 4072
rect 7837 4063 7895 4069
rect 7837 4060 7849 4063
rect 7524 4032 7849 4060
rect 7524 4020 7530 4032
rect 7837 4029 7849 4032
rect 7883 4029 7895 4063
rect 8110 4060 8116 4072
rect 8071 4032 8116 4060
rect 7837 4023 7895 4029
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 10137 4063 10195 4069
rect 10137 4029 10149 4063
rect 10183 4029 10195 4063
rect 10137 4023 10195 4029
rect 7392 3964 7880 3992
rect 7285 3955 7343 3961
rect 3844 3896 5672 3924
rect 6089 3927 6147 3933
rect 3844 3884 3850 3896
rect 6089 3893 6101 3927
rect 6135 3924 6147 3927
rect 6178 3924 6184 3936
rect 6135 3896 6184 3924
rect 6135 3893 6147 3896
rect 6089 3887 6147 3893
rect 6178 3884 6184 3896
rect 6236 3924 6242 3936
rect 6638 3924 6644 3936
rect 6236 3896 6644 3924
rect 6236 3884 6242 3896
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 7009 3927 7067 3933
rect 7009 3924 7021 3927
rect 6972 3896 7021 3924
rect 6972 3884 6978 3896
rect 7009 3893 7021 3896
rect 7055 3893 7067 3927
rect 7009 3887 7067 3893
rect 7650 3884 7656 3936
rect 7708 3924 7714 3936
rect 7745 3927 7803 3933
rect 7745 3924 7757 3927
rect 7708 3896 7757 3924
rect 7708 3884 7714 3896
rect 7745 3893 7757 3896
rect 7791 3893 7803 3927
rect 7852 3924 7880 3964
rect 10152 3924 10180 4023
rect 10226 4020 10232 4072
rect 10284 4060 10290 4072
rect 10411 4060 10439 4100
rect 10517 4097 10529 4131
rect 10563 4100 10588 4131
rect 10689 4131 10747 4137
rect 10563 4097 10575 4100
rect 10517 4091 10575 4097
rect 10689 4097 10701 4131
rect 10735 4097 10747 4131
rect 10962 4128 10968 4140
rect 10923 4100 10968 4128
rect 10689 4091 10747 4097
rect 10704 4060 10732 4091
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 11062 4131 11120 4137
rect 11062 4097 11074 4131
rect 11108 4097 11120 4131
rect 11514 4128 11520 4140
rect 11475 4100 11520 4128
rect 11062 4091 11120 4097
rect 10284 4032 10329 4060
rect 10411 4032 10732 4060
rect 10284 4020 10290 4032
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 11072 4060 11100 4091
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 13265 4063 13323 4069
rect 13265 4060 13277 4063
rect 10836 4032 11100 4060
rect 11624 4032 13277 4060
rect 10836 4020 10842 4032
rect 10962 3952 10968 4004
rect 11020 3992 11026 4004
rect 11624 3992 11652 4032
rect 13265 4029 13277 4032
rect 13311 4029 13323 4063
rect 13265 4023 13323 4029
rect 11020 3964 11652 3992
rect 11020 3952 11026 3964
rect 7852 3896 10180 3924
rect 11241 3927 11299 3933
rect 7745 3887 7803 3893
rect 11241 3893 11253 3927
rect 11287 3924 11299 3927
rect 11606 3924 11612 3936
rect 11287 3896 11612 3924
rect 11287 3893 11299 3896
rect 11241 3887 11299 3893
rect 11606 3884 11612 3896
rect 11664 3884 11670 3936
rect 1104 3834 13892 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 12214 3834
rect 12266 3782 12278 3834
rect 12330 3782 12342 3834
rect 12394 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 13892 3834
rect 1104 3760 13892 3782
rect 2958 3720 2964 3732
rect 1964 3692 2964 3720
rect 1762 3476 1768 3528
rect 1820 3516 1826 3528
rect 1964 3525 1992 3692
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3881 3723 3939 3729
rect 3881 3720 3893 3723
rect 3252 3692 3893 3720
rect 2038 3612 2044 3664
rect 2096 3652 2102 3664
rect 2409 3655 2467 3661
rect 2409 3652 2421 3655
rect 2096 3624 2421 3652
rect 2096 3612 2102 3624
rect 2409 3621 2421 3624
rect 2455 3621 2467 3655
rect 2409 3615 2467 3621
rect 2130 3544 2136 3596
rect 2188 3584 2194 3596
rect 2547 3587 2605 3593
rect 2547 3584 2559 3587
rect 2188 3556 2559 3584
rect 2188 3544 2194 3556
rect 2547 3553 2559 3556
rect 2593 3553 2605 3587
rect 2547 3547 2605 3553
rect 1856 3519 1914 3525
rect 1856 3516 1868 3519
rect 1820 3488 1868 3516
rect 1820 3476 1826 3488
rect 1856 3485 1868 3488
rect 1902 3485 1914 3519
rect 1856 3479 1914 3485
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3485 2007 3519
rect 1949 3479 2007 3485
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3485 2099 3519
rect 2222 3516 2228 3528
rect 2183 3488 2228 3516
rect 2041 3479 2099 3485
rect 1581 3451 1639 3457
rect 1581 3417 1593 3451
rect 1627 3417 1639 3451
rect 2056 3448 2084 3479
rect 2222 3476 2228 3488
rect 2280 3476 2286 3528
rect 2317 3519 2375 3525
rect 2317 3485 2329 3519
rect 2363 3516 2375 3519
rect 2406 3516 2412 3528
rect 2363 3488 2412 3516
rect 2363 3485 2375 3488
rect 2317 3479 2375 3485
rect 2406 3476 2412 3488
rect 2464 3476 2470 3528
rect 2682 3516 2688 3528
rect 2643 3488 2688 3516
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3485 3019 3519
rect 2961 3479 3019 3485
rect 2498 3448 2504 3460
rect 2056 3420 2504 3448
rect 1581 3411 1639 3417
rect 1596 3380 1624 3411
rect 2498 3408 2504 3420
rect 2556 3408 2562 3460
rect 2976 3448 3004 3479
rect 3050 3476 3056 3528
rect 3108 3516 3114 3528
rect 3252 3525 3280 3692
rect 3881 3689 3893 3692
rect 3927 3720 3939 3723
rect 3970 3720 3976 3732
rect 3927 3692 3976 3720
rect 3927 3689 3939 3692
rect 3881 3683 3939 3689
rect 3970 3680 3976 3692
rect 4028 3680 4034 3732
rect 4614 3680 4620 3732
rect 4672 3720 4678 3732
rect 4672 3692 5580 3720
rect 4672 3680 4678 3692
rect 3513 3655 3571 3661
rect 3513 3621 3525 3655
rect 3559 3621 3571 3655
rect 5552 3652 5580 3692
rect 5626 3680 5632 3732
rect 5684 3720 5690 3732
rect 7466 3720 7472 3732
rect 5684 3692 5764 3720
rect 5684 3680 5690 3692
rect 5736 3661 5764 3692
rect 6656 3692 7472 3720
rect 5721 3655 5779 3661
rect 5552 3624 5672 3652
rect 3513 3615 3571 3621
rect 3528 3584 3556 3615
rect 5644 3593 5672 3624
rect 5721 3621 5733 3655
rect 5767 3621 5779 3655
rect 5721 3615 5779 3621
rect 5353 3587 5411 3593
rect 5353 3584 5365 3587
rect 3528 3556 5365 3584
rect 5353 3553 5365 3556
rect 5399 3553 5411 3587
rect 5353 3547 5411 3553
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3584 5687 3587
rect 5902 3584 5908 3596
rect 5675 3556 5908 3584
rect 5675 3553 5687 3556
rect 5629 3547 5687 3553
rect 5902 3544 5908 3556
rect 5960 3584 5966 3596
rect 6656 3593 6684 3692
rect 7466 3680 7472 3692
rect 7524 3680 7530 3732
rect 8110 3680 8116 3732
rect 8168 3720 8174 3732
rect 9033 3723 9091 3729
rect 9033 3720 9045 3723
rect 8168 3692 9045 3720
rect 8168 3680 8174 3692
rect 9033 3689 9045 3692
rect 9079 3689 9091 3723
rect 9033 3683 9091 3689
rect 9490 3680 9496 3732
rect 9548 3720 9554 3732
rect 9677 3723 9735 3729
rect 9677 3720 9689 3723
rect 9548 3692 9689 3720
rect 9548 3680 9554 3692
rect 6641 3587 6699 3593
rect 6641 3584 6653 3587
rect 5960 3556 6653 3584
rect 5960 3544 5966 3556
rect 6641 3553 6653 3556
rect 6687 3553 6699 3587
rect 6914 3584 6920 3596
rect 6875 3556 6920 3584
rect 6641 3547 6699 3553
rect 6914 3544 6920 3556
rect 6972 3544 6978 3596
rect 7374 3544 7380 3596
rect 7432 3584 7438 3596
rect 8389 3587 8447 3593
rect 8389 3584 8401 3587
rect 7432 3556 8401 3584
rect 7432 3544 7438 3556
rect 8389 3553 8401 3556
rect 8435 3553 8447 3587
rect 8389 3547 8447 3553
rect 9398 3544 9404 3596
rect 9456 3584 9462 3596
rect 9600 3593 9628 3692
rect 9677 3689 9689 3692
rect 9723 3689 9735 3723
rect 9677 3683 9735 3689
rect 10045 3723 10103 3729
rect 10045 3689 10057 3723
rect 10091 3720 10103 3723
rect 10226 3720 10232 3732
rect 10091 3692 10232 3720
rect 10091 3689 10103 3692
rect 10045 3683 10103 3689
rect 10226 3680 10232 3692
rect 10284 3680 10290 3732
rect 12621 3723 12679 3729
rect 12621 3689 12633 3723
rect 12667 3720 12679 3723
rect 12802 3720 12808 3732
rect 12667 3692 12808 3720
rect 12667 3689 12679 3692
rect 12621 3683 12679 3689
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 9493 3587 9551 3593
rect 9493 3584 9505 3587
rect 9456 3556 9505 3584
rect 9456 3544 9462 3556
rect 9493 3553 9505 3556
rect 9539 3553 9551 3587
rect 9493 3547 9551 3553
rect 9585 3587 9643 3593
rect 9585 3553 9597 3587
rect 9631 3553 9643 3587
rect 9585 3547 9643 3553
rect 9769 3587 9827 3593
rect 9769 3553 9781 3587
rect 9815 3584 9827 3587
rect 10962 3584 10968 3596
rect 9815 3556 10968 3584
rect 9815 3553 9827 3556
rect 9769 3547 9827 3553
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 3145 3519 3203 3525
rect 3145 3516 3157 3519
rect 3108 3488 3157 3516
rect 3108 3476 3114 3488
rect 3145 3485 3157 3488
rect 3191 3485 3203 3519
rect 3145 3479 3203 3485
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3485 3295 3519
rect 3237 3479 3295 3485
rect 3381 3519 3439 3525
rect 3381 3485 3393 3519
rect 3427 3516 3439 3519
rect 3602 3516 3608 3528
rect 3427 3488 3608 3516
rect 3427 3485 3439 3488
rect 3381 3479 3439 3485
rect 3602 3476 3608 3488
rect 3660 3476 3666 3528
rect 5994 3516 6000 3528
rect 5955 3488 6000 3516
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 9214 3516 9220 3528
rect 9175 3488 9220 3516
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9677 3519 9735 3525
rect 9355 3488 9628 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9600 3460 9628 3488
rect 9677 3485 9689 3519
rect 9723 3516 9735 3519
rect 9858 3516 9864 3528
rect 9723 3488 9864 3516
rect 9723 3485 9735 3488
rect 9677 3479 9735 3485
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10229 3519 10287 3525
rect 10229 3516 10241 3519
rect 10008 3488 10241 3516
rect 10008 3476 10014 3488
rect 10229 3485 10241 3488
rect 10275 3485 10287 3519
rect 10229 3479 10287 3485
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3516 12495 3519
rect 12618 3516 12624 3528
rect 12483 3488 12624 3516
rect 12483 3485 12495 3488
rect 12437 3479 12495 3485
rect 12618 3476 12624 3488
rect 12676 3516 12682 3528
rect 12713 3519 12771 3525
rect 12713 3516 12725 3519
rect 12676 3488 12725 3516
rect 12676 3476 12682 3488
rect 12713 3485 12725 3488
rect 12759 3485 12771 3519
rect 12713 3479 12771 3485
rect 3878 3448 3884 3460
rect 2976 3420 3884 3448
rect 3878 3408 3884 3420
rect 3936 3448 3942 3460
rect 4062 3448 4068 3460
rect 3936 3420 4068 3448
rect 3936 3408 3942 3420
rect 4062 3408 4068 3420
rect 4120 3408 4126 3460
rect 4890 3408 4896 3460
rect 4948 3408 4954 3460
rect 5442 3408 5448 3460
rect 5500 3448 5506 3460
rect 6089 3451 6147 3457
rect 6089 3448 6101 3451
rect 5500 3420 6101 3448
rect 5500 3408 5506 3420
rect 6089 3417 6101 3420
rect 6135 3448 6147 3451
rect 6822 3448 6828 3460
rect 6135 3420 6828 3448
rect 6135 3417 6147 3420
rect 6089 3411 6147 3417
rect 6822 3408 6828 3420
rect 6880 3408 6886 3460
rect 7650 3408 7656 3460
rect 7708 3408 7714 3460
rect 9582 3408 9588 3460
rect 9640 3408 9646 3460
rect 10410 3408 10416 3460
rect 10468 3448 10474 3460
rect 10505 3451 10563 3457
rect 10505 3448 10517 3451
rect 10468 3420 10517 3448
rect 10468 3408 10474 3420
rect 10505 3417 10517 3420
rect 10551 3417 10563 3451
rect 11882 3448 11888 3460
rect 11730 3420 11888 3448
rect 10505 3411 10563 3417
rect 11882 3408 11888 3420
rect 11940 3408 11946 3460
rect 2590 3380 2596 3392
rect 1596 3352 2596 3380
rect 2590 3340 2596 3352
rect 2648 3340 2654 3392
rect 4706 3340 4712 3392
rect 4764 3380 4770 3392
rect 5258 3380 5264 3392
rect 4764 3352 5264 3380
rect 4764 3340 4770 3352
rect 5258 3340 5264 3352
rect 5316 3380 5322 3392
rect 5905 3383 5963 3389
rect 5905 3380 5917 3383
rect 5316 3352 5917 3380
rect 5316 3340 5322 3352
rect 5905 3349 5917 3352
rect 5951 3349 5963 3383
rect 5905 3343 5963 3349
rect 6273 3383 6331 3389
rect 6273 3349 6285 3383
rect 6319 3380 6331 3383
rect 6546 3380 6552 3392
rect 6319 3352 6552 3380
rect 6319 3349 6331 3352
rect 6273 3343 6331 3349
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 11974 3380 11980 3392
rect 11935 3352 11980 3380
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 12897 3383 12955 3389
rect 12897 3349 12909 3383
rect 12943 3380 12955 3383
rect 12986 3380 12992 3392
rect 12943 3352 12992 3380
rect 12943 3349 12955 3352
rect 12897 3343 12955 3349
rect 12986 3340 12992 3352
rect 13044 3340 13050 3392
rect 1104 3290 13892 3312
rect 1104 3238 8214 3290
rect 8266 3238 8278 3290
rect 8330 3238 8342 3290
rect 8394 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 13892 3290
rect 1104 3216 13892 3238
rect 2590 3136 2596 3188
rect 2648 3136 2654 3188
rect 4706 3176 4712 3188
rect 4667 3148 4712 3176
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 5261 3179 5319 3185
rect 5261 3145 5273 3179
rect 5307 3176 5319 3179
rect 5350 3176 5356 3188
rect 5307 3148 5356 3176
rect 5307 3145 5319 3148
rect 5261 3139 5319 3145
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 5537 3179 5595 3185
rect 5537 3145 5549 3179
rect 5583 3176 5595 3179
rect 6730 3176 6736 3188
rect 5583 3148 6736 3176
rect 5583 3145 5595 3148
rect 5537 3139 5595 3145
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 10502 3136 10508 3188
rect 10560 3176 10566 3188
rect 10689 3179 10747 3185
rect 10689 3176 10701 3179
rect 10560 3148 10701 3176
rect 10560 3136 10566 3148
rect 10689 3145 10701 3148
rect 10735 3145 10747 3179
rect 10689 3139 10747 3145
rect 10965 3179 11023 3185
rect 10965 3145 10977 3179
rect 11011 3176 11023 3179
rect 11974 3176 11980 3188
rect 11011 3148 11980 3176
rect 11011 3145 11023 3148
rect 10965 3139 11023 3145
rect 1670 3068 1676 3120
rect 1728 3108 1734 3120
rect 2608 3108 2636 3136
rect 3145 3111 3203 3117
rect 3145 3108 3157 3111
rect 1728 3080 1992 3108
rect 1728 3068 1734 3080
rect 1578 3040 1584 3052
rect 1539 3012 1584 3040
rect 1578 3000 1584 3012
rect 1636 3000 1642 3052
rect 1964 3049 1992 3080
rect 2240 3080 2636 3108
rect 2884 3080 3157 3108
rect 2240 3049 2268 3080
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3009 2283 3043
rect 2406 3040 2412 3052
rect 2367 3012 2412 3040
rect 2225 3003 2283 3009
rect 1872 2972 1900 3003
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 2498 3000 2504 3052
rect 2556 3040 2562 3052
rect 2884 3049 2912 3080
rect 3145 3077 3157 3080
rect 3191 3077 3203 3111
rect 5179 3111 5237 3117
rect 5179 3108 5191 3111
rect 3145 3071 3203 3077
rect 5000 3080 5191 3108
rect 2593 3043 2651 3049
rect 2593 3040 2605 3043
rect 2556 3012 2605 3040
rect 2556 3000 2562 3012
rect 2593 3009 2605 3012
rect 2639 3009 2651 3043
rect 2593 3003 2651 3009
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3009 2927 3043
rect 3050 3040 3056 3052
rect 3011 3012 3056 3040
rect 2869 3003 2927 3009
rect 3050 3000 3056 3012
rect 3108 3000 3114 3052
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3040 3939 3043
rect 4062 3040 4068 3052
rect 3927 3012 4068 3040
rect 3927 3009 3939 3012
rect 3881 3003 3939 3009
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 4801 3043 4859 3049
rect 4801 3009 4813 3043
rect 4847 3009 4859 3043
rect 4801 3003 4859 3009
rect 2038 2972 2044 2984
rect 1872 2944 2044 2972
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 4816 2972 4844 3003
rect 5000 2984 5028 3080
rect 5179 3077 5191 3080
rect 5225 3077 5237 3111
rect 5179 3071 5237 3077
rect 5445 3111 5503 3117
rect 5445 3077 5457 3111
rect 5491 3108 5503 3111
rect 6546 3108 6552 3120
rect 5491 3080 6552 3108
rect 5491 3077 5503 3080
rect 5445 3071 5503 3077
rect 6546 3068 6552 3080
rect 6604 3068 6610 3120
rect 7282 3108 7288 3120
rect 7243 3080 7288 3108
rect 7282 3068 7288 3080
rect 7340 3068 7346 3120
rect 8662 3068 8668 3120
rect 8720 3068 8726 3120
rect 9950 3108 9956 3120
rect 9692 3080 9956 3108
rect 5074 3000 5080 3052
rect 5132 3040 5138 3052
rect 5537 3043 5595 3049
rect 5132 3012 5177 3040
rect 5132 3000 5138 3012
rect 5537 3009 5549 3043
rect 5583 3040 5595 3043
rect 5629 3043 5687 3049
rect 5629 3040 5641 3043
rect 5583 3012 5641 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 5629 3009 5641 3012
rect 5675 3009 5687 3043
rect 5810 3040 5816 3052
rect 5771 3012 5816 3040
rect 5629 3003 5687 3009
rect 5810 3000 5816 3012
rect 5868 3040 5874 3052
rect 5994 3040 6000 3052
rect 5868 3012 6000 3040
rect 5868 3000 5874 3012
rect 5994 3000 6000 3012
rect 6052 3040 6058 3052
rect 6457 3043 6515 3049
rect 6457 3040 6469 3043
rect 6052 3012 6469 3040
rect 6052 3000 6058 3012
rect 6457 3009 6469 3012
rect 6503 3009 6515 3043
rect 6730 3040 6736 3052
rect 6691 3012 6736 3040
rect 6457 3003 6515 3009
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 7188 3043 7246 3049
rect 7188 3009 7200 3043
rect 7234 3040 7246 3043
rect 7234 3012 7328 3040
rect 7234 3009 7246 3012
rect 7188 3003 7246 3009
rect 4982 2972 4988 2984
rect 4816 2944 4988 2972
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 5258 2932 5264 2984
rect 5316 2972 5322 2984
rect 5828 2972 5856 3000
rect 6086 2972 6092 2984
rect 5316 2944 5856 2972
rect 6047 2944 6092 2972
rect 5316 2932 5322 2944
rect 6086 2932 6092 2944
rect 6144 2932 6150 2984
rect 6181 2975 6239 2981
rect 6181 2941 6193 2975
rect 6227 2972 6239 2975
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6227 2944 6837 2972
rect 6227 2941 6239 2944
rect 6181 2935 6239 2941
rect 6825 2941 6837 2944
rect 6871 2972 6883 2975
rect 6914 2972 6920 2984
rect 6871 2944 6920 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 6914 2932 6920 2944
rect 6972 2932 6978 2984
rect 7300 2972 7328 3012
rect 7374 3000 7380 3052
rect 7432 3040 7438 3052
rect 7432 3012 7477 3040
rect 7432 3000 7438 3012
rect 7558 3000 7564 3052
rect 7616 3040 7622 3052
rect 9692 3049 9720 3080
rect 9950 3068 9956 3080
rect 10008 3068 10014 3120
rect 10045 3111 10103 3117
rect 10045 3077 10057 3111
rect 10091 3108 10103 3111
rect 10980 3108 11008 3139
rect 11974 3136 11980 3148
rect 12032 3136 12038 3188
rect 10091 3080 11008 3108
rect 10091 3077 10103 3080
rect 10045 3071 10103 3077
rect 12986 3068 12992 3120
rect 13044 3068 13050 3120
rect 9677 3043 9735 3049
rect 7616 3012 7661 3040
rect 7616 3000 7622 3012
rect 9677 3009 9689 3043
rect 9723 3009 9735 3043
rect 9858 3040 9864 3052
rect 9819 3012 9864 3040
rect 9677 3003 9735 3009
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 10137 3043 10195 3049
rect 10137 3009 10149 3043
rect 10183 3009 10195 3043
rect 10137 3003 10195 3009
rect 9398 2972 9404 2984
rect 7300 2944 7972 2972
rect 9359 2944 9404 2972
rect 7944 2916 7972 2944
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 10152 2972 10180 3003
rect 10226 3000 10232 3052
rect 10284 3049 10290 3052
rect 10284 3043 10339 3049
rect 10284 3009 10293 3043
rect 10327 3040 10339 3043
rect 10686 3040 10692 3052
rect 10327 3012 10692 3040
rect 10327 3009 10339 3012
rect 10284 3003 10339 3009
rect 10284 3000 10290 3003
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 10870 3040 10876 3052
rect 10831 3012 10876 3040
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 10962 3000 10968 3052
rect 11020 3040 11026 3052
rect 11057 3043 11115 3049
rect 11057 3040 11069 3043
rect 11020 3012 11069 3040
rect 11020 3000 11026 3012
rect 11057 3009 11069 3012
rect 11103 3009 11115 3043
rect 11057 3003 11115 3009
rect 11514 3000 11520 3052
rect 11572 3040 11578 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11572 3012 11713 3040
rect 11572 3000 11578 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 11146 2972 11152 2984
rect 10152 2944 11152 2972
rect 11146 2932 11152 2944
rect 11204 2972 11210 2984
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 11204 2944 11253 2972
rect 11204 2932 11210 2944
rect 11241 2941 11253 2944
rect 11287 2941 11299 2975
rect 11241 2935 11299 2941
rect 11977 2975 12035 2981
rect 11977 2941 11989 2975
rect 12023 2972 12035 2975
rect 12710 2972 12716 2984
rect 12023 2944 12716 2972
rect 12023 2941 12035 2944
rect 11977 2935 12035 2941
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 4893 2907 4951 2913
rect 4893 2873 4905 2907
rect 4939 2904 4951 2907
rect 5718 2904 5724 2916
rect 4939 2876 5724 2904
rect 4939 2873 4951 2876
rect 4893 2867 4951 2873
rect 5718 2864 5724 2876
rect 5776 2864 5782 2916
rect 7006 2904 7012 2916
rect 6967 2876 7012 2904
rect 7006 2864 7012 2876
rect 7064 2864 7070 2916
rect 7926 2904 7932 2916
rect 7887 2876 7932 2904
rect 7926 2864 7932 2876
rect 7984 2864 7990 2916
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 10226 2904 10232 2916
rect 9732 2876 10232 2904
rect 9732 2864 9738 2876
rect 10226 2864 10232 2876
rect 10284 2864 10290 2916
rect 10410 2904 10416 2916
rect 10371 2876 10416 2904
rect 10410 2864 10416 2876
rect 10468 2864 10474 2916
rect 1670 2796 1676 2848
rect 1728 2836 1734 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 1728 2808 1777 2836
rect 1728 2796 1734 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 1765 2799 1823 2805
rect 2041 2839 2099 2845
rect 2041 2805 2053 2839
rect 2087 2836 2099 2839
rect 3786 2836 3792 2848
rect 2087 2808 3792 2836
rect 2087 2805 2099 2808
rect 2041 2799 2099 2805
rect 3786 2796 3792 2808
rect 3844 2796 3850 2848
rect 3970 2836 3976 2848
rect 3931 2808 3976 2836
rect 3970 2796 3976 2808
rect 4028 2796 4034 2848
rect 6454 2796 6460 2848
rect 6512 2836 6518 2848
rect 9692 2836 9720 2864
rect 13446 2836 13452 2848
rect 6512 2808 9720 2836
rect 13407 2808 13452 2836
rect 6512 2796 6518 2808
rect 13446 2796 13452 2808
rect 13504 2796 13510 2848
rect 1104 2746 13892 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 12214 2746
rect 12266 2694 12278 2746
rect 12330 2694 12342 2746
rect 12394 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 13892 2746
rect 1104 2672 13892 2694
rect 2958 2632 2964 2644
rect 1872 2604 2774 2632
rect 2919 2604 2964 2632
rect 1670 2428 1676 2440
rect 1631 2400 1676 2428
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 1762 2388 1768 2440
rect 1820 2428 1826 2440
rect 1872 2437 1900 2604
rect 2406 2564 2412 2576
rect 2367 2536 2412 2564
rect 2406 2524 2412 2536
rect 2464 2524 2470 2576
rect 2746 2564 2774 2604
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 3881 2635 3939 2641
rect 3881 2601 3893 2635
rect 3927 2632 3939 2635
rect 3970 2632 3976 2644
rect 3927 2604 3976 2632
rect 3927 2601 3939 2604
rect 3881 2595 3939 2601
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 4433 2635 4491 2641
rect 4433 2601 4445 2635
rect 4479 2632 4491 2635
rect 4798 2632 4804 2644
rect 4479 2604 4804 2632
rect 4479 2601 4491 2604
rect 4433 2595 4491 2601
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 5626 2592 5632 2644
rect 5684 2632 5690 2644
rect 7282 2632 7288 2644
rect 5684 2604 7288 2632
rect 5684 2592 5690 2604
rect 7282 2592 7288 2604
rect 7340 2632 7346 2644
rect 7558 2632 7564 2644
rect 7340 2604 7420 2632
rect 7519 2604 7564 2632
rect 7340 2592 7346 2604
rect 3050 2564 3056 2576
rect 2746 2536 3056 2564
rect 3050 2524 3056 2536
rect 3108 2524 3114 2576
rect 3142 2524 3148 2576
rect 3200 2564 3206 2576
rect 4890 2564 4896 2576
rect 3200 2536 4896 2564
rect 3200 2524 3206 2536
rect 4890 2524 4896 2536
rect 4948 2524 4954 2576
rect 5074 2564 5080 2576
rect 5035 2536 5080 2564
rect 5074 2524 5080 2536
rect 5132 2524 5138 2576
rect 7392 2564 7420 2604
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 8573 2635 8631 2641
rect 8573 2601 8585 2635
rect 8619 2632 8631 2635
rect 8662 2632 8668 2644
rect 8619 2604 8668 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 9033 2635 9091 2641
rect 9033 2601 9045 2635
rect 9079 2632 9091 2635
rect 9398 2632 9404 2644
rect 9079 2604 9404 2632
rect 9079 2601 9091 2604
rect 9033 2595 9091 2601
rect 9398 2592 9404 2604
rect 9456 2592 9462 2644
rect 11882 2632 11888 2644
rect 11843 2604 11888 2632
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 5460 2536 6132 2564
rect 7392 2536 7696 2564
rect 5460 2508 5488 2536
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 2593 2499 2651 2505
rect 2593 2496 2605 2499
rect 1995 2468 2605 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 2593 2465 2605 2468
rect 2639 2465 2651 2499
rect 3605 2499 3663 2505
rect 3605 2496 3617 2499
rect 2593 2459 2651 2465
rect 3140 2468 3617 2496
rect 1856 2431 1914 2437
rect 1856 2428 1868 2431
rect 1820 2400 1868 2428
rect 1820 2388 1826 2400
rect 1856 2397 1868 2400
rect 1902 2397 1914 2431
rect 2038 2428 2044 2440
rect 1999 2400 2044 2428
rect 1856 2391 1914 2397
rect 2038 2388 2044 2400
rect 2096 2388 2102 2440
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2397 2283 2431
rect 2225 2391 2283 2397
rect 1578 2320 1584 2372
rect 1636 2360 1642 2372
rect 2240 2360 2268 2391
rect 2498 2388 2504 2440
rect 2556 2428 2562 2440
rect 3140 2437 3168 2468
rect 3605 2465 3617 2468
rect 3651 2496 3663 2499
rect 4062 2496 4068 2508
rect 3651 2468 4068 2496
rect 3651 2465 3663 2468
rect 3605 2459 3663 2465
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 5442 2496 5448 2508
rect 5403 2468 5448 2496
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2465 5871 2499
rect 5813 2459 5871 2465
rect 5905 2499 5963 2505
rect 5905 2465 5917 2499
rect 5951 2496 5963 2499
rect 5994 2496 6000 2508
rect 5951 2468 6000 2496
rect 5951 2465 5963 2468
rect 5905 2459 5963 2465
rect 2685 2431 2743 2437
rect 2685 2428 2697 2431
rect 2556 2400 2697 2428
rect 2556 2388 2562 2400
rect 2685 2397 2697 2400
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 3125 2431 3183 2437
rect 3125 2397 3137 2431
rect 3171 2397 3183 2431
rect 3125 2391 3183 2397
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2397 3295 2431
rect 3786 2428 3792 2440
rect 3747 2400 3792 2428
rect 3237 2391 3295 2397
rect 1636 2332 2268 2360
rect 3252 2360 3280 2391
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 4311 2431 4369 2437
rect 4311 2397 4323 2431
rect 4357 2428 4369 2431
rect 4614 2428 4620 2440
rect 4357 2400 4620 2428
rect 4357 2397 4369 2400
rect 4311 2391 4369 2397
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 5258 2428 5264 2440
rect 5219 2400 5264 2428
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5534 2428 5540 2440
rect 5495 2400 5540 2428
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 5626 2388 5632 2440
rect 5684 2428 5690 2440
rect 5720 2431 5778 2437
rect 5720 2428 5732 2431
rect 5684 2400 5732 2428
rect 5684 2388 5690 2400
rect 5720 2397 5732 2400
rect 5766 2397 5778 2431
rect 5720 2391 5778 2397
rect 3510 2360 3516 2372
rect 3252 2332 3516 2360
rect 1636 2320 1642 2332
rect 3510 2320 3516 2332
rect 3568 2320 3574 2372
rect 4709 2363 4767 2369
rect 4080 2332 4384 2360
rect 2038 2252 2044 2304
rect 2096 2292 2102 2304
rect 4080 2292 4108 2332
rect 4246 2292 4252 2304
rect 2096 2264 4108 2292
rect 4207 2264 4252 2292
rect 2096 2252 2102 2264
rect 4246 2252 4252 2264
rect 4304 2252 4310 2304
rect 4356 2292 4384 2332
rect 4709 2329 4721 2363
rect 4755 2360 4767 2363
rect 4890 2360 4896 2372
rect 4755 2332 4896 2360
rect 4755 2329 4767 2332
rect 4709 2323 4767 2329
rect 4890 2320 4896 2332
rect 4948 2320 4954 2372
rect 5828 2360 5856 2459
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6104 2437 6132 2536
rect 6641 2499 6699 2505
rect 6641 2465 6653 2499
rect 6687 2496 6699 2499
rect 6914 2496 6920 2508
rect 6687 2468 6920 2496
rect 6687 2465 6699 2468
rect 6641 2459 6699 2465
rect 6914 2456 6920 2468
rect 6972 2496 6978 2508
rect 7101 2499 7159 2505
rect 7101 2496 7113 2499
rect 6972 2468 7113 2496
rect 6972 2456 6978 2468
rect 7101 2465 7113 2468
rect 7147 2496 7159 2499
rect 7374 2496 7380 2508
rect 7147 2468 7380 2496
rect 7147 2465 7159 2468
rect 7101 2459 7159 2465
rect 7374 2456 7380 2468
rect 7432 2456 7438 2508
rect 6089 2431 6147 2437
rect 6089 2397 6101 2431
rect 6135 2397 6147 2431
rect 6089 2391 6147 2397
rect 6270 2388 6276 2440
rect 6328 2428 6334 2440
rect 6549 2431 6607 2437
rect 6328 2400 6373 2428
rect 6328 2388 6334 2400
rect 6549 2397 6561 2431
rect 6595 2428 6607 2431
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 6595 2400 7205 2428
rect 6595 2397 6607 2400
rect 6549 2391 6607 2397
rect 7193 2397 7205 2400
rect 7239 2428 7251 2431
rect 7558 2428 7564 2440
rect 7239 2400 7564 2428
rect 7239 2397 7251 2400
rect 7193 2391 7251 2397
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 7668 2437 7696 2536
rect 7926 2524 7932 2576
rect 7984 2564 7990 2576
rect 8113 2567 8171 2573
rect 8113 2564 8125 2567
rect 7984 2536 8125 2564
rect 7984 2524 7990 2536
rect 8113 2533 8125 2536
rect 8159 2564 8171 2567
rect 12713 2567 12771 2573
rect 12713 2564 12725 2567
rect 8159 2536 9444 2564
rect 8159 2533 8171 2536
rect 8113 2527 8171 2533
rect 7668 2431 7741 2437
rect 7668 2400 7695 2431
rect 7683 2397 7695 2400
rect 7729 2428 7741 2431
rect 8110 2428 8116 2440
rect 7729 2400 8116 2428
rect 7729 2397 7741 2400
rect 7683 2391 7741 2397
rect 8110 2388 8116 2400
rect 8168 2428 8174 2440
rect 8205 2431 8263 2437
rect 8205 2428 8217 2431
rect 8168 2400 8217 2428
rect 8168 2388 8174 2400
rect 8205 2397 8217 2400
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 6178 2360 6184 2372
rect 5828 2332 6184 2360
rect 6178 2320 6184 2332
rect 6236 2320 6242 2372
rect 6825 2363 6883 2369
rect 6825 2329 6837 2363
rect 6871 2329 6883 2363
rect 6825 2323 6883 2329
rect 6840 2292 6868 2323
rect 4356 2264 6868 2292
rect 7745 2295 7803 2301
rect 7745 2261 7757 2295
rect 7791 2292 7803 2295
rect 8312 2292 8340 2536
rect 9416 2448 9444 2536
rect 12406 2536 12725 2564
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 8754 2428 8760 2440
rect 8715 2400 8760 2428
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 9323 2437 9444 2448
rect 9600 2468 9781 2496
rect 9600 2440 9628 2468
rect 9769 2465 9781 2468
rect 9815 2465 9827 2499
rect 9769 2459 9827 2465
rect 9858 2456 9864 2508
rect 9916 2496 9922 2508
rect 12406 2496 12434 2536
rect 12713 2533 12725 2536
rect 12759 2533 12771 2567
rect 12713 2527 12771 2533
rect 13265 2499 13323 2505
rect 13265 2496 13277 2499
rect 9916 2468 12434 2496
rect 13004 2468 13277 2496
rect 9916 2456 9922 2468
rect 9212 2431 9270 2437
rect 9212 2397 9224 2431
rect 9258 2397 9270 2431
rect 9212 2391 9270 2397
rect 9308 2431 9444 2437
rect 9308 2397 9320 2431
rect 9354 2420 9444 2431
rect 9582 2428 9588 2440
rect 9354 2397 9366 2420
rect 9495 2400 9588 2428
rect 9308 2391 9366 2397
rect 7791 2264 8340 2292
rect 9232 2292 9260 2391
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2397 9735 2431
rect 9950 2428 9956 2440
rect 9911 2400 9956 2428
rect 9677 2391 9735 2397
rect 9398 2360 9404 2372
rect 9359 2332 9404 2360
rect 9398 2320 9404 2332
rect 9456 2320 9462 2372
rect 9692 2360 9720 2391
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 11514 2388 11520 2440
rect 11572 2428 11578 2440
rect 12069 2431 12127 2437
rect 12069 2428 12081 2431
rect 11572 2400 12081 2428
rect 11572 2388 11578 2400
rect 12069 2397 12081 2400
rect 12115 2428 12127 2431
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12115 2400 12357 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 12345 2397 12357 2400
rect 12391 2428 12403 2431
rect 12618 2428 12624 2440
rect 12391 2400 12624 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 12618 2388 12624 2400
rect 12676 2388 12682 2440
rect 12710 2388 12716 2440
rect 12768 2428 12774 2440
rect 13004 2437 13032 2468
rect 13265 2465 13277 2468
rect 13311 2496 13323 2499
rect 13446 2496 13452 2508
rect 13311 2468 13452 2496
rect 13311 2465 13323 2468
rect 13265 2459 13323 2465
rect 13446 2456 13452 2468
rect 13504 2456 13510 2508
rect 12877 2431 12935 2437
rect 12877 2428 12889 2431
rect 12768 2400 12889 2428
rect 12768 2388 12774 2400
rect 12877 2397 12889 2400
rect 12923 2428 12935 2431
rect 12989 2431 13047 2437
rect 12923 2397 12940 2428
rect 12877 2391 12940 2397
rect 12989 2397 13001 2431
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 9858 2360 9864 2372
rect 9692 2332 9864 2360
rect 9692 2292 9720 2332
rect 9858 2320 9864 2332
rect 9916 2320 9922 2372
rect 10226 2360 10232 2372
rect 10187 2332 10232 2360
rect 10226 2320 10232 2332
rect 10284 2320 10290 2372
rect 12912 2360 12940 2391
rect 13357 2363 13415 2369
rect 13357 2360 13369 2363
rect 11072 2304 11100 2346
rect 12912 2332 13369 2360
rect 13357 2329 13369 2332
rect 13403 2360 13415 2363
rect 13446 2360 13452 2372
rect 13403 2332 13452 2360
rect 13403 2329 13415 2332
rect 13357 2323 13415 2329
rect 13446 2320 13452 2332
rect 13504 2320 13510 2372
rect 9232 2264 9720 2292
rect 7791 2261 7803 2264
rect 7745 2255 7803 2261
rect 11054 2252 11060 2304
rect 11112 2252 11118 2304
rect 11146 2252 11152 2304
rect 11204 2292 11210 2304
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 11204 2264 11713 2292
rect 11204 2252 11210 2264
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 11701 2255 11759 2261
rect 12529 2295 12587 2301
rect 12529 2261 12541 2295
rect 12575 2292 12587 2295
rect 12618 2292 12624 2304
rect 12575 2264 12624 2292
rect 12575 2261 12587 2264
rect 12529 2255 12587 2261
rect 12618 2252 12624 2264
rect 12676 2252 12682 2304
rect 1104 2202 13892 2224
rect 1104 2150 8214 2202
rect 8266 2150 8278 2202
rect 8330 2150 8342 2202
rect 8394 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 13892 2202
rect 1104 2128 13892 2150
rect 1578 2048 1584 2100
rect 1636 2088 1642 2100
rect 1636 2060 3464 2088
rect 1636 2048 1642 2060
rect 2866 1980 2872 2032
rect 2924 1980 2930 2032
rect 3436 2020 3464 2060
rect 3510 2048 3516 2100
rect 3568 2088 3574 2100
rect 3605 2091 3663 2097
rect 3605 2088 3617 2091
rect 3568 2060 3617 2088
rect 3568 2048 3574 2060
rect 3605 2057 3617 2060
rect 3651 2057 3663 2091
rect 8110 2088 8116 2100
rect 3605 2051 3663 2057
rect 6380 2060 7972 2088
rect 8071 2060 8116 2088
rect 3436 1992 4476 2020
rect 3513 1955 3571 1961
rect 3513 1921 3525 1955
rect 3559 1952 3571 1955
rect 3786 1952 3792 1964
rect 3559 1924 3792 1952
rect 3559 1921 3571 1924
rect 3513 1915 3571 1921
rect 3786 1912 3792 1924
rect 3844 1912 3850 1964
rect 3881 1955 3939 1961
rect 3881 1921 3893 1955
rect 3927 1921 3939 1955
rect 3881 1915 3939 1921
rect 4065 1955 4123 1961
rect 4065 1921 4077 1955
rect 4111 1952 4123 1955
rect 4246 1952 4252 1964
rect 4111 1924 4252 1952
rect 4111 1921 4123 1924
rect 4065 1915 4123 1921
rect 1578 1884 1584 1896
rect 1539 1856 1584 1884
rect 1578 1844 1584 1856
rect 1636 1844 1642 1896
rect 1857 1887 1915 1893
rect 1857 1853 1869 1887
rect 1903 1884 1915 1887
rect 3326 1884 3332 1896
rect 1903 1856 3332 1884
rect 1903 1853 1915 1856
rect 1857 1847 1915 1853
rect 3326 1844 3332 1856
rect 3384 1844 3390 1896
rect 3896 1884 3924 1915
rect 4246 1912 4252 1924
rect 4304 1912 4310 1964
rect 4448 1884 4476 1992
rect 5258 1980 5264 2032
rect 5316 1980 5322 2032
rect 5718 2020 5724 2032
rect 5679 1992 5724 2020
rect 5718 1980 5724 1992
rect 5776 1980 5782 2032
rect 5994 1884 6000 1896
rect 3896 1856 4292 1884
rect 4448 1856 6000 1884
rect 3329 1751 3387 1757
rect 3329 1717 3341 1751
rect 3375 1748 3387 1751
rect 4062 1748 4068 1760
rect 3375 1720 4068 1748
rect 3375 1717 3387 1720
rect 3329 1711 3387 1717
rect 4062 1708 4068 1720
rect 4120 1708 4126 1760
rect 4264 1757 4292 1856
rect 5994 1844 6000 1856
rect 6052 1884 6058 1896
rect 6380 1893 6408 2060
rect 7374 1980 7380 2032
rect 7432 1980 7438 2032
rect 7944 1952 7972 2060
rect 8110 2048 8116 2060
rect 8168 2048 8174 2100
rect 9950 2088 9956 2100
rect 8404 2060 9956 2088
rect 8404 1961 8432 2060
rect 9950 2048 9956 2060
rect 10008 2048 10014 2100
rect 10226 2048 10232 2100
rect 10284 2088 10290 2100
rect 10396 2091 10454 2097
rect 10396 2088 10408 2091
rect 10284 2060 10408 2088
rect 10284 2048 10290 2060
rect 10396 2057 10408 2060
rect 10442 2057 10454 2091
rect 11054 2088 11060 2100
rect 11015 2060 11060 2088
rect 10396 2051 10454 2057
rect 11054 2048 11060 2060
rect 11112 2048 11118 2100
rect 9398 1980 9404 2032
rect 9456 1980 9462 2032
rect 10689 2023 10747 2029
rect 10689 1989 10701 2023
rect 10735 2020 10747 2023
rect 11146 2020 11152 2032
rect 10735 1992 11152 2020
rect 10735 1989 10747 1992
rect 10689 1983 10747 1989
rect 11146 1980 11152 1992
rect 11204 1980 11210 2032
rect 11330 1980 11336 2032
rect 11388 2020 11394 2032
rect 11388 1992 12282 2020
rect 11388 1980 11394 1992
rect 8389 1955 8447 1961
rect 8389 1952 8401 1955
rect 7944 1924 8401 1952
rect 8389 1921 8401 1924
rect 8435 1921 8447 1955
rect 10545 1955 10603 1961
rect 10545 1952 10557 1955
rect 8389 1915 8447 1921
rect 9876 1924 10557 1952
rect 9876 1896 9904 1924
rect 10545 1921 10557 1924
rect 10591 1921 10603 1955
rect 10545 1915 10603 1921
rect 10781 1955 10839 1961
rect 10781 1921 10793 1955
rect 10827 1921 10839 1955
rect 10962 1952 10968 1964
rect 10923 1924 10968 1952
rect 10781 1915 10839 1921
rect 6365 1887 6423 1893
rect 6365 1884 6377 1887
rect 6052 1856 6377 1884
rect 6052 1844 6058 1856
rect 6365 1853 6377 1856
rect 6411 1853 6423 1887
rect 6638 1884 6644 1896
rect 6599 1856 6644 1884
rect 6365 1847 6423 1853
rect 6638 1844 6644 1856
rect 6696 1844 6702 1896
rect 8662 1884 8668 1896
rect 8623 1856 8668 1884
rect 8662 1844 8668 1856
rect 8720 1844 8726 1896
rect 9858 1844 9864 1896
rect 9916 1844 9922 1896
rect 10134 1884 10140 1896
rect 10047 1856 10140 1884
rect 10134 1844 10140 1856
rect 10192 1884 10198 1896
rect 10796 1884 10824 1915
rect 10962 1912 10968 1924
rect 11020 1912 11026 1964
rect 11238 1952 11244 1964
rect 11199 1924 11244 1952
rect 11238 1912 11244 1924
rect 11296 1912 11302 1964
rect 10870 1884 10876 1896
rect 10192 1856 10876 1884
rect 10192 1844 10198 1856
rect 10870 1844 10876 1856
rect 10928 1844 10934 1896
rect 11514 1884 11520 1896
rect 10980 1856 11520 1884
rect 9950 1776 9956 1828
rect 10008 1816 10014 1828
rect 10980 1816 11008 1856
rect 11514 1844 11520 1856
rect 11572 1844 11578 1896
rect 11793 1887 11851 1893
rect 11793 1884 11805 1887
rect 11624 1856 11805 1884
rect 10008 1788 11008 1816
rect 10008 1776 10014 1788
rect 11146 1776 11152 1828
rect 11204 1816 11210 1828
rect 11624 1816 11652 1856
rect 11793 1853 11805 1856
rect 11839 1853 11851 1887
rect 11793 1847 11851 1853
rect 11204 1788 11652 1816
rect 11204 1776 11210 1788
rect 4249 1751 4307 1757
rect 4249 1717 4261 1751
rect 4295 1748 4307 1751
rect 4614 1748 4620 1760
rect 4295 1720 4620 1748
rect 4295 1717 4307 1720
rect 4249 1711 4307 1717
rect 4614 1708 4620 1720
rect 4672 1708 4678 1760
rect 5534 1708 5540 1760
rect 5592 1748 5598 1760
rect 9858 1748 9864 1760
rect 5592 1720 9864 1748
rect 5592 1708 5598 1720
rect 9858 1708 9864 1720
rect 9916 1708 9922 1760
rect 11974 1708 11980 1760
rect 12032 1748 12038 1760
rect 13265 1751 13323 1757
rect 13265 1748 13277 1751
rect 12032 1720 13277 1748
rect 12032 1708 12038 1720
rect 13265 1717 13277 1720
rect 13311 1717 13323 1751
rect 13265 1711 13323 1717
rect 1104 1658 13892 1680
rect 1104 1606 4214 1658
rect 4266 1606 4278 1658
rect 4330 1606 4342 1658
rect 4394 1606 4406 1658
rect 4458 1606 4470 1658
rect 4522 1606 12214 1658
rect 12266 1606 12278 1658
rect 12330 1606 12342 1658
rect 12394 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 13892 1658
rect 1104 1584 13892 1606
rect 2777 1547 2835 1553
rect 2777 1513 2789 1547
rect 2823 1544 2835 1547
rect 2866 1544 2872 1556
rect 2823 1516 2872 1544
rect 2823 1513 2835 1516
rect 2777 1507 2835 1513
rect 2866 1504 2872 1516
rect 2924 1504 2930 1556
rect 3326 1504 3332 1556
rect 3384 1544 3390 1556
rect 3881 1547 3939 1553
rect 3881 1544 3893 1547
rect 3384 1516 3893 1544
rect 3384 1504 3390 1516
rect 3881 1513 3893 1516
rect 3927 1513 3939 1547
rect 3881 1507 3939 1513
rect 3970 1504 3976 1556
rect 4028 1544 4034 1556
rect 4028 1516 4752 1544
rect 4028 1504 4034 1516
rect 4246 1476 4252 1488
rect 3528 1448 4252 1476
rect 1578 1300 1584 1352
rect 1636 1340 1642 1352
rect 1765 1343 1823 1349
rect 1765 1340 1777 1343
rect 1636 1312 1777 1340
rect 1636 1300 1642 1312
rect 1765 1309 1777 1312
rect 1811 1309 1823 1343
rect 1765 1303 1823 1309
rect 2593 1343 2651 1349
rect 2593 1309 2605 1343
rect 2639 1340 2651 1343
rect 3142 1340 3148 1352
rect 2639 1312 3148 1340
rect 2639 1309 2651 1312
rect 2593 1303 2651 1309
rect 3142 1300 3148 1312
rect 3200 1300 3206 1352
rect 3528 1349 3556 1448
rect 4246 1436 4252 1448
rect 4304 1476 4310 1488
rect 4614 1476 4620 1488
rect 4304 1448 4620 1476
rect 4304 1436 4310 1448
rect 4614 1436 4620 1448
rect 4672 1436 4678 1488
rect 4724 1476 4752 1516
rect 4982 1504 4988 1556
rect 5040 1544 5046 1556
rect 5169 1547 5227 1553
rect 5169 1544 5181 1547
rect 5040 1516 5181 1544
rect 5040 1504 5046 1516
rect 5169 1513 5181 1516
rect 5215 1513 5227 1547
rect 5350 1544 5356 1556
rect 5311 1516 5356 1544
rect 5169 1507 5227 1513
rect 5350 1504 5356 1516
rect 5408 1504 5414 1556
rect 5442 1504 5448 1556
rect 5500 1544 5506 1556
rect 6089 1547 6147 1553
rect 6089 1544 6101 1547
rect 5500 1516 6101 1544
rect 5500 1504 5506 1516
rect 6089 1513 6101 1516
rect 6135 1513 6147 1547
rect 6638 1544 6644 1556
rect 6599 1516 6644 1544
rect 6089 1507 6147 1513
rect 6638 1504 6644 1516
rect 6696 1504 6702 1556
rect 7374 1504 7380 1556
rect 7432 1544 7438 1556
rect 7469 1547 7527 1553
rect 7469 1544 7481 1547
rect 7432 1516 7481 1544
rect 7432 1504 7438 1516
rect 7469 1513 7481 1516
rect 7515 1513 7527 1547
rect 7469 1507 7527 1513
rect 9398 1504 9404 1556
rect 9456 1544 9462 1556
rect 9585 1547 9643 1553
rect 9585 1544 9597 1547
rect 9456 1516 9597 1544
rect 9456 1504 9462 1516
rect 9585 1513 9597 1516
rect 9631 1513 9643 1547
rect 11330 1544 11336 1556
rect 11291 1516 11336 1544
rect 9585 1507 9643 1513
rect 11330 1504 11336 1516
rect 11388 1504 11394 1556
rect 13446 1544 13452 1556
rect 13407 1516 13452 1544
rect 13446 1504 13452 1516
rect 13504 1504 13510 1556
rect 5534 1476 5540 1488
rect 4724 1448 5540 1476
rect 5534 1436 5540 1448
rect 5592 1436 5598 1488
rect 8662 1436 8668 1488
rect 8720 1476 8726 1488
rect 8941 1479 8999 1485
rect 8941 1476 8953 1479
rect 8720 1448 8953 1476
rect 8720 1436 8726 1448
rect 8941 1445 8953 1448
rect 8987 1445 8999 1479
rect 8941 1439 8999 1445
rect 9214 1436 9220 1488
rect 9272 1476 9278 1488
rect 10134 1476 10140 1488
rect 9272 1448 10140 1476
rect 9272 1436 9278 1448
rect 10134 1436 10140 1448
rect 10192 1436 10198 1488
rect 3878 1368 3884 1420
rect 3936 1408 3942 1420
rect 3936 1380 4476 1408
rect 3936 1368 3942 1380
rect 3421 1343 3479 1349
rect 3421 1309 3433 1343
rect 3467 1309 3479 1343
rect 3421 1303 3479 1309
rect 3513 1343 3571 1349
rect 3513 1309 3525 1343
rect 3559 1309 3571 1343
rect 3513 1303 3571 1309
rect 3436 1272 3464 1303
rect 3970 1300 3976 1352
rect 4028 1349 4034 1352
rect 4028 1343 4071 1349
rect 4059 1309 4071 1343
rect 4028 1303 4071 1309
rect 4028 1300 4034 1303
rect 4154 1300 4160 1352
rect 4212 1340 4218 1352
rect 4448 1349 4476 1380
rect 4890 1368 4896 1420
rect 4948 1408 4954 1420
rect 4948 1380 5580 1408
rect 4948 1368 4954 1380
rect 4433 1343 4491 1349
rect 4212 1312 4257 1340
rect 4212 1300 4218 1312
rect 4433 1309 4445 1343
rect 4479 1309 4491 1343
rect 5442 1340 5448 1352
rect 5403 1312 5448 1340
rect 4433 1303 4491 1309
rect 5442 1300 5448 1312
rect 5500 1300 5506 1352
rect 5552 1349 5580 1380
rect 5626 1368 5632 1420
rect 5684 1408 5690 1420
rect 11238 1408 11244 1420
rect 5684 1380 6224 1408
rect 5684 1368 5690 1380
rect 5537 1343 5595 1349
rect 5537 1309 5549 1343
rect 5583 1309 5595 1343
rect 5537 1303 5595 1309
rect 5810 1300 5816 1352
rect 5868 1340 5874 1352
rect 6196 1349 6224 1380
rect 9646 1380 11244 1408
rect 6181 1343 6239 1349
rect 5868 1312 5913 1340
rect 5868 1300 5874 1312
rect 6181 1309 6193 1343
rect 6227 1309 6239 1343
rect 6181 1303 6239 1309
rect 6270 1300 6276 1352
rect 6328 1340 6334 1352
rect 6365 1343 6423 1349
rect 6365 1340 6377 1343
rect 6328 1312 6377 1340
rect 6328 1300 6334 1312
rect 6365 1309 6377 1312
rect 6411 1309 6423 1343
rect 6546 1340 6552 1352
rect 6507 1312 6552 1340
rect 6365 1303 6423 1309
rect 6546 1300 6552 1312
rect 6604 1300 6610 1352
rect 7285 1343 7343 1349
rect 7285 1309 7297 1343
rect 7331 1309 7343 1343
rect 7285 1303 7343 1309
rect 4172 1272 4200 1300
rect 3436 1244 4200 1272
rect 4246 1232 4252 1284
rect 4304 1272 4310 1284
rect 5828 1272 5856 1300
rect 7300 1272 7328 1303
rect 8754 1300 8760 1352
rect 8812 1340 8818 1352
rect 9401 1343 9459 1349
rect 9401 1340 9413 1343
rect 8812 1312 9413 1340
rect 8812 1300 8818 1312
rect 9401 1309 9413 1312
rect 9447 1340 9459 1343
rect 9646 1340 9674 1380
rect 11164 1349 11192 1380
rect 11238 1368 11244 1380
rect 11296 1368 11302 1420
rect 11514 1368 11520 1420
rect 11572 1408 11578 1420
rect 11701 1411 11759 1417
rect 11701 1408 11713 1411
rect 11572 1380 11713 1408
rect 11572 1368 11578 1380
rect 11701 1377 11713 1380
rect 11747 1377 11759 1411
rect 11974 1408 11980 1420
rect 11935 1380 11980 1408
rect 11701 1371 11759 1377
rect 11974 1368 11980 1380
rect 12032 1368 12038 1420
rect 9447 1312 9674 1340
rect 11149 1343 11207 1349
rect 9447 1309 9459 1312
rect 9401 1303 9459 1309
rect 11149 1309 11161 1343
rect 11195 1309 11207 1343
rect 11149 1303 11207 1309
rect 4304 1244 4349 1272
rect 5828 1244 7328 1272
rect 9125 1275 9183 1281
rect 4304 1232 4310 1244
rect 9125 1241 9137 1275
rect 9171 1272 9183 1275
rect 9214 1272 9220 1284
rect 9171 1244 9220 1272
rect 9171 1241 9183 1244
rect 9125 1235 9183 1241
rect 9214 1232 9220 1244
rect 9272 1232 9278 1284
rect 9309 1275 9367 1281
rect 9309 1241 9321 1275
rect 9355 1241 9367 1275
rect 9309 1235 9367 1241
rect 1578 1204 1584 1216
rect 1539 1176 1584 1204
rect 1578 1164 1584 1176
rect 1636 1164 1642 1216
rect 3513 1207 3571 1213
rect 3513 1173 3525 1207
rect 3559 1204 3571 1207
rect 3786 1204 3792 1216
rect 3559 1176 3792 1204
rect 3559 1173 3571 1176
rect 3513 1167 3571 1173
rect 3786 1164 3792 1176
rect 3844 1164 3850 1216
rect 5258 1164 5264 1216
rect 5316 1204 5322 1216
rect 5629 1207 5687 1213
rect 5629 1204 5641 1207
rect 5316 1176 5641 1204
rect 5316 1164 5322 1176
rect 5629 1173 5641 1176
rect 5675 1173 5687 1207
rect 9324 1204 9352 1235
rect 12618 1232 12624 1284
rect 12676 1232 12682 1284
rect 9674 1204 9680 1216
rect 9324 1176 9680 1204
rect 5629 1167 5687 1173
rect 9674 1164 9680 1176
rect 9732 1164 9738 1216
rect 1104 1114 13892 1136
rect 1104 1062 8214 1114
rect 8266 1062 8278 1114
rect 8330 1062 8342 1114
rect 8394 1062 8406 1114
rect 8458 1062 8470 1114
rect 8522 1062 13892 1114
rect 1104 1040 13892 1062
<< via1 >>
rect 3976 13744 4028 13796
rect 7564 13744 7616 13796
rect 572 13676 624 13728
rect 7196 13676 7248 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 12214 13574 12266 13626
rect 12278 13574 12330 13626
rect 12342 13574 12394 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 1400 13268 1452 13320
rect 2136 13268 2188 13320
rect 3332 13311 3384 13320
rect 2780 13200 2832 13252
rect 2872 13200 2924 13252
rect 3332 13277 3341 13311
rect 3341 13277 3375 13311
rect 3375 13277 3384 13311
rect 3332 13268 3384 13277
rect 3608 13268 3660 13320
rect 5080 13311 5132 13320
rect 5080 13277 5089 13311
rect 5089 13277 5123 13311
rect 5123 13277 5132 13311
rect 5080 13268 5132 13277
rect 5816 13311 5868 13320
rect 5816 13277 5825 13311
rect 5825 13277 5859 13311
rect 5859 13277 5868 13311
rect 5816 13268 5868 13277
rect 6920 13336 6972 13388
rect 7196 13379 7248 13388
rect 7196 13345 7205 13379
rect 7205 13345 7239 13379
rect 7239 13345 7248 13379
rect 7196 13336 7248 13345
rect 8024 13336 8076 13388
rect 9680 13268 9732 13320
rect 10876 13336 10928 13388
rect 10968 13268 11020 13320
rect 12624 13336 12676 13388
rect 12348 13311 12400 13320
rect 12348 13277 12357 13311
rect 12357 13277 12391 13311
rect 12391 13277 12400 13311
rect 12348 13268 12400 13277
rect 4804 13243 4856 13252
rect 4804 13209 4813 13243
rect 4813 13209 4847 13243
rect 4847 13209 4856 13243
rect 4804 13200 4856 13209
rect 6368 13200 6420 13252
rect 9404 13243 9456 13252
rect 9404 13209 9413 13243
rect 9413 13209 9447 13243
rect 9447 13209 9456 13243
rect 9404 13200 9456 13209
rect 9864 13200 9916 13252
rect 10048 13243 10100 13252
rect 10048 13209 10057 13243
rect 10057 13209 10091 13243
rect 10091 13209 10100 13243
rect 10048 13200 10100 13209
rect 10140 13243 10192 13252
rect 10140 13209 10149 13243
rect 10149 13209 10183 13243
rect 10183 13209 10192 13243
rect 10140 13200 10192 13209
rect 12072 13200 12124 13252
rect 12808 13243 12860 13252
rect 12808 13209 12817 13243
rect 12817 13209 12851 13243
rect 12851 13209 12860 13243
rect 12808 13200 12860 13209
rect 12900 13243 12952 13252
rect 12900 13209 12909 13243
rect 12909 13209 12943 13243
rect 12943 13209 12952 13243
rect 12900 13200 12952 13209
rect 7288 13175 7340 13184
rect 7288 13141 7297 13175
rect 7297 13141 7331 13175
rect 7331 13141 7340 13175
rect 7288 13132 7340 13141
rect 10600 13175 10652 13184
rect 10600 13141 10609 13175
rect 10609 13141 10643 13175
rect 10643 13141 10652 13175
rect 10600 13132 10652 13141
rect 11888 13175 11940 13184
rect 11888 13141 11897 13175
rect 11897 13141 11931 13175
rect 11931 13141 11940 13175
rect 11888 13132 11940 13141
rect 8214 13030 8266 13082
rect 8278 13030 8330 13082
rect 8342 13030 8394 13082
rect 8406 13030 8458 13082
rect 8470 13030 8522 13082
rect 1676 12928 1728 12980
rect 6368 12971 6420 12980
rect 2780 12860 2832 12912
rect 5816 12903 5868 12912
rect 5816 12869 5825 12903
rect 5825 12869 5859 12903
rect 5859 12869 5868 12903
rect 5816 12860 5868 12869
rect 6368 12937 6377 12971
rect 6377 12937 6411 12971
rect 6411 12937 6420 12971
rect 6368 12928 6420 12937
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 3332 12792 3384 12844
rect 3608 12792 3660 12844
rect 5080 12792 5132 12844
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 7748 12835 7800 12844
rect 7748 12801 7757 12835
rect 7757 12801 7791 12835
rect 7791 12801 7800 12835
rect 7748 12792 7800 12801
rect 8024 12835 8076 12844
rect 8024 12801 8033 12835
rect 8033 12801 8067 12835
rect 8067 12801 8076 12835
rect 8024 12792 8076 12801
rect 9956 12860 10008 12912
rect 10048 12860 10100 12912
rect 9680 12835 9732 12844
rect 9680 12801 9689 12835
rect 9689 12801 9723 12835
rect 9723 12801 9732 12835
rect 9680 12792 9732 12801
rect 12348 12928 12400 12980
rect 6920 12724 6972 12776
rect 9404 12724 9456 12776
rect 12716 12792 12768 12844
rect 11336 12767 11388 12776
rect 4804 12699 4856 12708
rect 4804 12665 4813 12699
rect 4813 12665 4847 12699
rect 4847 12665 4856 12699
rect 4804 12656 4856 12665
rect 3884 12588 3936 12640
rect 5724 12588 5776 12640
rect 11336 12733 11345 12767
rect 11345 12733 11379 12767
rect 11379 12733 11388 12767
rect 11336 12724 11388 12733
rect 12072 12656 12124 12708
rect 12808 12656 12860 12708
rect 13176 12699 13228 12708
rect 13176 12665 13185 12699
rect 13185 12665 13219 12699
rect 13219 12665 13228 12699
rect 13176 12656 13228 12665
rect 11520 12588 11572 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 12214 12486 12266 12538
rect 12278 12486 12330 12538
rect 12342 12486 12394 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 3332 12427 3384 12436
rect 3332 12393 3341 12427
rect 3341 12393 3375 12427
rect 3375 12393 3384 12427
rect 3332 12384 3384 12393
rect 3608 12384 3660 12436
rect 4160 12248 4212 12300
rect 4344 12291 4396 12300
rect 4344 12257 4353 12291
rect 4353 12257 4387 12291
rect 4387 12257 4396 12291
rect 6920 12384 6972 12436
rect 7748 12359 7800 12368
rect 4344 12248 4396 12257
rect 5724 12291 5776 12300
rect 5724 12257 5733 12291
rect 5733 12257 5767 12291
rect 5767 12257 5776 12291
rect 5724 12248 5776 12257
rect 7748 12325 7757 12359
rect 7757 12325 7791 12359
rect 7791 12325 7800 12359
rect 7748 12316 7800 12325
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 2872 12223 2924 12232
rect 2872 12189 2881 12223
rect 2881 12189 2915 12223
rect 2915 12189 2924 12223
rect 2872 12180 2924 12189
rect 3332 12180 3384 12232
rect 4804 12180 4856 12232
rect 9680 12384 9732 12436
rect 10140 12427 10192 12436
rect 10140 12393 10149 12427
rect 10149 12393 10183 12427
rect 10183 12393 10192 12427
rect 10140 12384 10192 12393
rect 11336 12384 11388 12436
rect 12900 12427 12952 12436
rect 12900 12393 12909 12427
rect 12909 12393 12943 12427
rect 12943 12393 12952 12427
rect 12900 12384 12952 12393
rect 9220 12291 9272 12300
rect 9220 12257 9229 12291
rect 9229 12257 9263 12291
rect 9263 12257 9272 12291
rect 9220 12248 9272 12257
rect 10232 12248 10284 12300
rect 14372 12316 14424 12368
rect 10968 12291 11020 12300
rect 10968 12257 10977 12291
rect 10977 12257 11011 12291
rect 11011 12257 11020 12291
rect 10968 12248 11020 12257
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 9956 12223 10008 12232
rect 9956 12189 9965 12223
rect 9965 12189 9999 12223
rect 9999 12189 10008 12223
rect 9956 12180 10008 12189
rect 11520 12223 11572 12232
rect 3240 12155 3292 12164
rect 3240 12121 3249 12155
rect 3249 12121 3283 12155
rect 3283 12121 3292 12155
rect 3240 12112 3292 12121
rect 5724 12112 5776 12164
rect 9220 12112 9272 12164
rect 11520 12189 11529 12223
rect 11529 12189 11563 12223
rect 11563 12189 11572 12223
rect 11520 12180 11572 12189
rect 12072 12180 12124 12232
rect 12716 12223 12768 12232
rect 12716 12189 12725 12223
rect 12725 12189 12759 12223
rect 12759 12189 12768 12223
rect 12716 12180 12768 12189
rect 13176 12223 13228 12232
rect 13176 12189 13185 12223
rect 13185 12189 13219 12223
rect 13219 12189 13228 12223
rect 13176 12180 13228 12189
rect 4896 12044 4948 12096
rect 6368 12044 6420 12096
rect 8576 12087 8628 12096
rect 8576 12053 8585 12087
rect 8585 12053 8619 12087
rect 8619 12053 8628 12087
rect 8576 12044 8628 12053
rect 9036 12044 9088 12096
rect 9956 12044 10008 12096
rect 11060 12044 11112 12096
rect 13452 12044 13504 12096
rect 8214 11942 8266 11994
rect 8278 11942 8330 11994
rect 8342 11942 8394 11994
rect 8406 11942 8458 11994
rect 8470 11942 8522 11994
rect 1400 11883 1452 11892
rect 1400 11849 1409 11883
rect 1409 11849 1443 11883
rect 1443 11849 1452 11883
rect 1400 11840 1452 11849
rect 3884 11840 3936 11892
rect 4160 11840 4212 11892
rect 5264 11840 5316 11892
rect 3240 11772 3292 11824
rect 9772 11840 9824 11892
rect 10048 11840 10100 11892
rect 2872 11747 2924 11756
rect 2872 11713 2881 11747
rect 2881 11713 2915 11747
rect 2915 11713 2924 11747
rect 8576 11815 8628 11824
rect 8576 11781 8585 11815
rect 8585 11781 8619 11815
rect 8619 11781 8628 11815
rect 8576 11772 8628 11781
rect 2872 11704 2924 11713
rect 5632 11704 5684 11756
rect 1860 11679 1912 11688
rect 1860 11645 1869 11679
rect 1869 11645 1903 11679
rect 1903 11645 1912 11679
rect 1860 11636 1912 11645
rect 2228 11679 2280 11688
rect 1492 11568 1544 11620
rect 2228 11645 2237 11679
rect 2237 11645 2271 11679
rect 2271 11645 2280 11679
rect 2228 11636 2280 11645
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 3424 11679 3476 11688
rect 2780 11636 2832 11645
rect 3424 11645 3433 11679
rect 3433 11645 3467 11679
rect 3467 11645 3476 11679
rect 3424 11636 3476 11645
rect 3332 11611 3384 11620
rect 3332 11577 3341 11611
rect 3341 11577 3375 11611
rect 3375 11577 3384 11611
rect 3332 11568 3384 11577
rect 4344 11636 4396 11688
rect 3976 11500 4028 11552
rect 5172 11679 5224 11688
rect 5172 11645 5181 11679
rect 5181 11645 5215 11679
rect 5215 11645 5224 11679
rect 5172 11636 5224 11645
rect 5264 11679 5316 11688
rect 5264 11645 5273 11679
rect 5273 11645 5307 11679
rect 5307 11645 5316 11679
rect 5264 11636 5316 11645
rect 4988 11568 5040 11620
rect 5356 11611 5408 11620
rect 5356 11577 5365 11611
rect 5365 11577 5399 11611
rect 5399 11577 5408 11611
rect 5356 11568 5408 11577
rect 4896 11500 4948 11552
rect 6460 11704 6512 11756
rect 7104 11747 7156 11756
rect 7104 11713 7113 11747
rect 7113 11713 7147 11747
rect 7147 11713 7156 11747
rect 7104 11704 7156 11713
rect 7472 11747 7524 11756
rect 7472 11713 7481 11747
rect 7481 11713 7515 11747
rect 7515 11713 7524 11747
rect 7472 11704 7524 11713
rect 9956 11772 10008 11824
rect 10324 11772 10376 11824
rect 10140 11704 10192 11756
rect 10416 11704 10468 11756
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 13452 11815 13504 11824
rect 13452 11781 13461 11815
rect 13461 11781 13495 11815
rect 13495 11781 13504 11815
rect 13452 11772 13504 11781
rect 10784 11704 10836 11713
rect 12992 11704 13044 11756
rect 13268 11747 13320 11756
rect 13268 11713 13277 11747
rect 13277 11713 13311 11747
rect 13311 11713 13320 11747
rect 13268 11704 13320 11713
rect 5816 11679 5868 11688
rect 5816 11645 5825 11679
rect 5825 11645 5859 11679
rect 5859 11645 5868 11679
rect 5816 11636 5868 11645
rect 6092 11568 6144 11620
rect 8300 11636 8352 11688
rect 9220 11636 9272 11688
rect 9496 11636 9548 11688
rect 10508 11679 10560 11688
rect 10508 11645 10517 11679
rect 10517 11645 10551 11679
rect 10551 11645 10560 11679
rect 10508 11636 10560 11645
rect 8944 11568 8996 11620
rect 9864 11568 9916 11620
rect 5908 11500 5960 11552
rect 6736 11500 6788 11552
rect 9404 11500 9456 11552
rect 13084 11636 13136 11688
rect 11060 11568 11112 11620
rect 10876 11500 10928 11552
rect 12900 11500 12952 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 12214 11398 12266 11450
rect 12278 11398 12330 11450
rect 12342 11398 12394 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 2780 11296 2832 11348
rect 5632 11296 5684 11348
rect 3240 11228 3292 11280
rect 4988 11228 5040 11280
rect 5264 11271 5316 11280
rect 5264 11237 5273 11271
rect 5273 11237 5307 11271
rect 5307 11237 5316 11271
rect 7104 11296 7156 11348
rect 8300 11339 8352 11348
rect 8300 11305 8309 11339
rect 8309 11305 8343 11339
rect 8343 11305 8352 11339
rect 8300 11296 8352 11305
rect 8944 11339 8996 11348
rect 8944 11305 8953 11339
rect 8953 11305 8987 11339
rect 8987 11305 8996 11339
rect 8944 11296 8996 11305
rect 10140 11339 10192 11348
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 10140 11296 10192 11305
rect 5264 11228 5316 11237
rect 6828 11228 6880 11280
rect 11152 11296 11204 11348
rect 11888 11296 11940 11348
rect 3884 11160 3936 11212
rect 2228 11092 2280 11144
rect 3056 11135 3108 11144
rect 3056 11101 3065 11135
rect 3065 11101 3099 11135
rect 3099 11101 3108 11135
rect 3056 11092 3108 11101
rect 3332 11092 3384 11144
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 4528 11092 4580 11144
rect 4896 11135 4948 11144
rect 4896 11101 4905 11135
rect 4905 11101 4939 11135
rect 4939 11101 4948 11135
rect 4896 11092 4948 11101
rect 5908 11092 5960 11144
rect 6092 11135 6144 11144
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6460 11160 6512 11212
rect 6092 11092 6144 11101
rect 5448 11024 5500 11076
rect 7840 11160 7892 11212
rect 9404 11203 9456 11212
rect 7472 11092 7524 11144
rect 8576 11135 8628 11144
rect 8576 11101 8585 11135
rect 8585 11101 8619 11135
rect 8619 11101 8628 11135
rect 8576 11092 8628 11101
rect 9404 11169 9413 11203
rect 9413 11169 9447 11203
rect 9447 11169 9456 11203
rect 9404 11160 9456 11169
rect 9496 11203 9548 11212
rect 9496 11169 9505 11203
rect 9505 11169 9539 11203
rect 9539 11169 9548 11203
rect 9496 11160 9548 11169
rect 10232 11160 10284 11212
rect 9864 11092 9916 11144
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 11428 11228 11480 11280
rect 12808 11271 12860 11280
rect 12808 11237 12817 11271
rect 12817 11237 12851 11271
rect 12851 11237 12860 11271
rect 12808 11228 12860 11237
rect 10876 11203 10928 11212
rect 10876 11169 10885 11203
rect 10885 11169 10919 11203
rect 10919 11169 10928 11203
rect 10876 11160 10928 11169
rect 11060 11135 11112 11144
rect 2964 10956 3016 11008
rect 6920 11024 6972 11076
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 11060 11092 11112 11101
rect 11152 11092 11204 11144
rect 12348 11092 12400 11144
rect 13452 11092 13504 11144
rect 10968 10956 11020 11008
rect 11060 10956 11112 11008
rect 13360 10999 13412 11008
rect 13360 10965 13369 10999
rect 13369 10965 13403 10999
rect 13403 10965 13412 10999
rect 13360 10956 13412 10965
rect 8214 10854 8266 10906
rect 8278 10854 8330 10906
rect 8342 10854 8394 10906
rect 8406 10854 8458 10906
rect 8470 10854 8522 10906
rect 2228 10752 2280 10804
rect 3424 10752 3476 10804
rect 5172 10752 5224 10804
rect 5816 10752 5868 10804
rect 6184 10752 6236 10804
rect 3332 10727 3384 10736
rect 3332 10693 3341 10727
rect 3341 10693 3375 10727
rect 3375 10693 3384 10727
rect 3332 10684 3384 10693
rect 5356 10684 5408 10736
rect 6368 10727 6420 10736
rect 1676 10659 1728 10668
rect 1676 10625 1685 10659
rect 1685 10625 1719 10659
rect 1719 10625 1728 10659
rect 1676 10616 1728 10625
rect 1492 10591 1544 10600
rect 1492 10557 1501 10591
rect 1501 10557 1535 10591
rect 1535 10557 1544 10591
rect 1492 10548 1544 10557
rect 2872 10616 2924 10668
rect 3056 10616 3108 10668
rect 4528 10659 4580 10668
rect 4528 10625 4537 10659
rect 4537 10625 4571 10659
rect 4571 10625 4580 10659
rect 4528 10616 4580 10625
rect 6368 10693 6377 10727
rect 6377 10693 6411 10727
rect 6411 10693 6420 10727
rect 6368 10684 6420 10693
rect 6644 10684 6696 10736
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 6000 10616 6052 10668
rect 6460 10616 6512 10668
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 7196 10659 7248 10668
rect 7196 10625 7205 10659
rect 7205 10625 7239 10659
rect 7239 10625 7248 10659
rect 7748 10684 7800 10736
rect 7196 10616 7248 10625
rect 7564 10616 7616 10668
rect 5908 10480 5960 10532
rect 6092 10480 6144 10532
rect 7012 10480 7064 10532
rect 7564 10480 7616 10532
rect 7748 10548 7800 10600
rect 8484 10616 8536 10668
rect 10048 10616 10100 10668
rect 10324 10752 10376 10804
rect 11060 10795 11112 10804
rect 10232 10684 10284 10736
rect 10416 10659 10468 10668
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 10416 10616 10468 10625
rect 10508 10616 10560 10668
rect 11060 10761 11069 10795
rect 11069 10761 11103 10795
rect 11103 10761 11112 10795
rect 11060 10752 11112 10761
rect 11520 10795 11572 10804
rect 11520 10761 11529 10795
rect 11529 10761 11563 10795
rect 11563 10761 11572 10795
rect 11520 10752 11572 10761
rect 11980 10795 12032 10804
rect 11980 10761 11989 10795
rect 11989 10761 12023 10795
rect 12023 10761 12032 10795
rect 11980 10752 12032 10761
rect 12900 10727 12952 10736
rect 12900 10693 12909 10727
rect 12909 10693 12943 10727
rect 12943 10693 12952 10727
rect 12900 10684 12952 10693
rect 13360 10684 13412 10736
rect 12348 10659 12400 10668
rect 12348 10625 12357 10659
rect 12357 10625 12391 10659
rect 12391 10625 12400 10659
rect 12348 10616 12400 10625
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 13268 10616 13320 10668
rect 7840 10480 7892 10532
rect 9680 10548 9732 10600
rect 9864 10591 9916 10600
rect 9864 10557 9873 10591
rect 9873 10557 9907 10591
rect 9907 10557 9916 10591
rect 9864 10548 9916 10557
rect 12624 10548 12676 10600
rect 12900 10548 12952 10600
rect 11520 10480 11572 10532
rect 5172 10412 5224 10464
rect 5816 10412 5868 10464
rect 6184 10412 6236 10464
rect 6828 10412 6880 10464
rect 8484 10412 8536 10464
rect 9680 10412 9732 10464
rect 9956 10455 10008 10464
rect 9956 10421 9965 10455
rect 9965 10421 9999 10455
rect 9999 10421 10008 10455
rect 9956 10412 10008 10421
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 10692 10412 10744 10464
rect 11152 10412 11204 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 12214 10310 12266 10362
rect 12278 10310 12330 10362
rect 12342 10310 12394 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 3056 10251 3108 10260
rect 3056 10217 3065 10251
rect 3065 10217 3099 10251
rect 3099 10217 3108 10251
rect 3056 10208 3108 10217
rect 5724 10251 5776 10260
rect 5724 10217 5733 10251
rect 5733 10217 5767 10251
rect 5767 10217 5776 10251
rect 5724 10208 5776 10217
rect 6000 10208 6052 10260
rect 6920 10251 6972 10260
rect 6276 10140 6328 10192
rect 6920 10217 6929 10251
rect 6929 10217 6963 10251
rect 6963 10217 6972 10251
rect 6920 10208 6972 10217
rect 7104 10208 7156 10260
rect 7472 10208 7524 10260
rect 10600 10208 10652 10260
rect 10968 10208 11020 10260
rect 11152 10251 11204 10260
rect 11152 10217 11161 10251
rect 11161 10217 11195 10251
rect 11195 10217 11204 10251
rect 11152 10208 11204 10217
rect 11428 10208 11480 10260
rect 12992 10208 13044 10260
rect 7196 10140 7248 10192
rect 8116 10140 8168 10192
rect 9956 10140 10008 10192
rect 10692 10183 10744 10192
rect 10692 10149 10701 10183
rect 10701 10149 10735 10183
rect 10735 10149 10744 10183
rect 10692 10140 10744 10149
rect 5448 10115 5500 10124
rect 5448 10081 5457 10115
rect 5457 10081 5491 10115
rect 5491 10081 5500 10115
rect 5448 10072 5500 10081
rect 6092 10115 6144 10124
rect 6092 10081 6101 10115
rect 6101 10081 6135 10115
rect 6135 10081 6144 10115
rect 6092 10072 6144 10081
rect 3884 10004 3936 10056
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 5908 10004 5960 10056
rect 6184 10047 6236 10056
rect 2964 9979 3016 9988
rect 2964 9945 2973 9979
rect 2973 9945 3007 9979
rect 3007 9945 3016 9979
rect 2964 9936 3016 9945
rect 6184 10013 6193 10047
rect 6193 10013 6227 10047
rect 6227 10013 6236 10047
rect 6184 10004 6236 10013
rect 7012 10072 7064 10124
rect 7104 10004 7156 10056
rect 7564 10047 7616 10056
rect 6736 9936 6788 9988
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 7840 10004 7892 10056
rect 7656 9936 7708 9988
rect 8668 9936 8720 9988
rect 8852 9936 8904 9988
rect 9496 10047 9548 10056
rect 9496 10013 9505 10047
rect 9505 10013 9539 10047
rect 9539 10013 9548 10047
rect 9496 10004 9548 10013
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 10508 10004 10560 10056
rect 12900 10072 12952 10124
rect 9864 9936 9916 9988
rect 3240 9868 3292 9920
rect 4896 9868 4948 9920
rect 8024 9911 8076 9920
rect 8024 9877 8033 9911
rect 8033 9877 8067 9911
rect 8067 9877 8076 9911
rect 8024 9868 8076 9877
rect 11244 9936 11296 9988
rect 12808 10004 12860 10056
rect 13084 9979 13136 9988
rect 13084 9945 13093 9979
rect 13093 9945 13127 9979
rect 13127 9945 13136 9979
rect 13084 9936 13136 9945
rect 11336 9868 11388 9920
rect 12532 9911 12584 9920
rect 12532 9877 12541 9911
rect 12541 9877 12575 9911
rect 12575 9877 12584 9911
rect 12532 9868 12584 9877
rect 13176 9911 13228 9920
rect 13176 9877 13185 9911
rect 13185 9877 13219 9911
rect 13219 9877 13228 9911
rect 13176 9868 13228 9877
rect 8214 9766 8266 9818
rect 8278 9766 8330 9818
rect 8342 9766 8394 9818
rect 8406 9766 8458 9818
rect 8470 9766 8522 9818
rect 1492 9664 1544 9716
rect 2228 9528 2280 9580
rect 3332 9596 3384 9648
rect 3884 9528 3936 9580
rect 2964 9435 3016 9444
rect 2964 9401 2973 9435
rect 2973 9401 3007 9435
rect 3007 9401 3016 9435
rect 2964 9392 3016 9401
rect 6184 9664 6236 9716
rect 6920 9664 6972 9716
rect 7656 9664 7708 9716
rect 5080 9639 5132 9648
rect 5080 9605 5089 9639
rect 5089 9605 5123 9639
rect 5123 9605 5132 9639
rect 5080 9596 5132 9605
rect 9496 9664 9548 9716
rect 10416 9664 10468 9716
rect 8208 9596 8260 9648
rect 8852 9596 8904 9648
rect 9036 9639 9088 9648
rect 9036 9605 9045 9639
rect 9045 9605 9079 9639
rect 9079 9605 9088 9639
rect 9036 9596 9088 9605
rect 9128 9596 9180 9648
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 7196 9571 7248 9580
rect 6828 9528 6880 9537
rect 7196 9537 7205 9571
rect 7205 9537 7239 9571
rect 7239 9537 7248 9571
rect 7196 9528 7248 9537
rect 7564 9528 7616 9580
rect 8484 9571 8536 9580
rect 8484 9537 8493 9571
rect 8493 9537 8527 9571
rect 8527 9537 8536 9571
rect 8484 9528 8536 9537
rect 5448 9460 5500 9512
rect 4620 9392 4672 9444
rect 8024 9392 8076 9444
rect 8760 9460 8812 9512
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 10232 9528 10284 9580
rect 10508 9460 10560 9512
rect 11060 9596 11112 9648
rect 11428 9596 11480 9648
rect 10876 9571 10928 9580
rect 10876 9537 10885 9571
rect 10885 9537 10919 9571
rect 10919 9537 10928 9571
rect 11520 9571 11572 9580
rect 10876 9528 10928 9537
rect 11152 9460 11204 9512
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 13360 9571 13412 9580
rect 13360 9537 13369 9571
rect 13369 9537 13403 9571
rect 13403 9537 13412 9571
rect 13360 9528 13412 9537
rect 11612 9460 11664 9512
rect 3792 9324 3844 9376
rect 6920 9367 6972 9376
rect 6920 9333 6929 9367
rect 6929 9333 6963 9367
rect 6963 9333 6972 9367
rect 6920 9324 6972 9333
rect 7012 9367 7064 9376
rect 7012 9333 7021 9367
rect 7021 9333 7055 9367
rect 7055 9333 7064 9367
rect 7748 9367 7800 9376
rect 7012 9324 7064 9333
rect 7748 9333 7757 9367
rect 7757 9333 7791 9367
rect 7791 9333 7800 9367
rect 7748 9324 7800 9333
rect 7932 9324 7984 9376
rect 9220 9324 9272 9376
rect 9680 9392 9732 9444
rect 10140 9392 10192 9444
rect 10784 9392 10836 9444
rect 12808 9435 12860 9444
rect 12808 9401 12817 9435
rect 12817 9401 12851 9435
rect 12851 9401 12860 9435
rect 12808 9392 12860 9401
rect 11336 9324 11388 9376
rect 13268 9367 13320 9376
rect 13268 9333 13277 9367
rect 13277 9333 13311 9367
rect 13311 9333 13320 9367
rect 13268 9324 13320 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 12214 9222 12266 9274
rect 12278 9222 12330 9274
rect 12342 9222 12394 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 2228 9163 2280 9172
rect 2228 9129 2237 9163
rect 2237 9129 2271 9163
rect 2271 9129 2280 9163
rect 2228 9120 2280 9129
rect 1492 8984 1544 9036
rect 1768 9027 1820 9036
rect 1768 8993 1777 9027
rect 1777 8993 1811 9027
rect 1811 8993 1820 9027
rect 1768 8984 1820 8993
rect 8116 9120 8168 9172
rect 8300 9120 8352 9172
rect 8944 9120 8996 9172
rect 9128 9163 9180 9172
rect 9128 9129 9137 9163
rect 9137 9129 9171 9163
rect 9171 9129 9180 9163
rect 9128 9120 9180 9129
rect 10140 9120 10192 9172
rect 10232 9120 10284 9172
rect 11152 9120 11204 9172
rect 2964 9052 3016 9104
rect 3332 9095 3384 9104
rect 3332 9061 3341 9095
rect 3341 9061 3375 9095
rect 3375 9061 3384 9095
rect 3332 9052 3384 9061
rect 3884 9095 3936 9104
rect 3884 9061 3893 9095
rect 3893 9061 3927 9095
rect 3927 9061 3936 9095
rect 3884 9052 3936 9061
rect 6920 9052 6972 9104
rect 7288 9095 7340 9104
rect 7288 9061 7297 9095
rect 7297 9061 7331 9095
rect 7331 9061 7340 9095
rect 7288 9052 7340 9061
rect 7564 9052 7616 9104
rect 9680 9052 9732 9104
rect 9772 9052 9824 9104
rect 10324 9052 10376 9104
rect 3792 9027 3844 9036
rect 3792 8993 3801 9027
rect 3801 8993 3835 9027
rect 3835 8993 3844 9027
rect 3792 8984 3844 8993
rect 4620 8984 4672 9036
rect 3240 8916 3292 8968
rect 3608 8959 3660 8968
rect 3608 8925 3617 8959
rect 3617 8925 3651 8959
rect 3651 8925 3660 8959
rect 7196 8984 7248 9036
rect 8760 8984 8812 9036
rect 10048 8984 10100 9036
rect 10784 8984 10836 9036
rect 12808 9052 12860 9104
rect 3608 8916 3660 8925
rect 6736 8959 6788 8968
rect 3148 8891 3200 8900
rect 3148 8857 3157 8891
rect 3157 8857 3191 8891
rect 3191 8857 3200 8891
rect 3148 8848 3200 8857
rect 5356 8848 5408 8900
rect 6736 8925 6745 8959
rect 6745 8925 6779 8959
rect 6779 8925 6788 8959
rect 6736 8916 6788 8925
rect 7472 8959 7524 8968
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 7012 8848 7064 8900
rect 7748 8848 7800 8900
rect 8024 8848 8076 8900
rect 9036 8848 9088 8900
rect 10048 8891 10100 8900
rect 3424 8823 3476 8832
rect 3424 8789 3433 8823
rect 3433 8789 3467 8823
rect 3467 8789 3476 8823
rect 3424 8780 3476 8789
rect 4804 8823 4856 8832
rect 4804 8789 4813 8823
rect 4813 8789 4847 8823
rect 4847 8789 4856 8823
rect 4804 8780 4856 8789
rect 7196 8780 7248 8832
rect 7472 8780 7524 8832
rect 10048 8857 10057 8891
rect 10057 8857 10091 8891
rect 10091 8857 10100 8891
rect 10048 8848 10100 8857
rect 11060 8916 11112 8968
rect 11612 8916 11664 8968
rect 13268 8984 13320 9036
rect 12624 8959 12676 8968
rect 10692 8891 10744 8900
rect 10692 8857 10701 8891
rect 10701 8857 10735 8891
rect 10735 8857 10744 8891
rect 10692 8848 10744 8857
rect 10876 8891 10928 8900
rect 10876 8857 10885 8891
rect 10885 8857 10919 8891
rect 10919 8857 10928 8891
rect 10876 8848 10928 8857
rect 10968 8891 11020 8900
rect 10968 8857 10977 8891
rect 10977 8857 11011 8891
rect 11011 8857 11020 8891
rect 10968 8848 11020 8857
rect 11520 8848 11572 8900
rect 12624 8925 12633 8959
rect 12633 8925 12667 8959
rect 12667 8925 12676 8959
rect 12624 8916 12676 8925
rect 13360 8959 13412 8968
rect 13360 8925 13369 8959
rect 13369 8925 13403 8959
rect 13403 8925 13412 8959
rect 13360 8916 13412 8925
rect 12716 8848 12768 8900
rect 10324 8780 10376 8832
rect 10508 8823 10560 8832
rect 10508 8789 10517 8823
rect 10517 8789 10551 8823
rect 10551 8789 10560 8823
rect 10508 8780 10560 8789
rect 10600 8780 10652 8832
rect 11796 8823 11848 8832
rect 11796 8789 11805 8823
rect 11805 8789 11839 8823
rect 11839 8789 11848 8823
rect 11796 8780 11848 8789
rect 8214 8678 8266 8730
rect 8278 8678 8330 8730
rect 8342 8678 8394 8730
rect 8406 8678 8458 8730
rect 8470 8678 8522 8730
rect 3148 8551 3200 8560
rect 3148 8517 3157 8551
rect 3157 8517 3191 8551
rect 3191 8517 3200 8551
rect 3148 8508 3200 8517
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 3608 8508 3660 8560
rect 7380 8576 7432 8628
rect 7472 8576 7524 8628
rect 7932 8619 7984 8628
rect 7932 8585 7941 8619
rect 7941 8585 7975 8619
rect 7975 8585 7984 8619
rect 7932 8576 7984 8585
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 3332 8440 3384 8492
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 4620 8440 4672 8492
rect 5724 8440 5776 8492
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 5356 8304 5408 8356
rect 7748 8508 7800 8560
rect 8208 8551 8260 8560
rect 8208 8517 8217 8551
rect 8217 8517 8251 8551
rect 8251 8517 8260 8551
rect 8208 8508 8260 8517
rect 9128 8576 9180 8628
rect 8944 8508 8996 8560
rect 10232 8576 10284 8628
rect 7472 8415 7524 8424
rect 7472 8381 7481 8415
rect 7481 8381 7515 8415
rect 7515 8381 7524 8415
rect 7472 8372 7524 8381
rect 7564 8372 7616 8424
rect 7932 8440 7984 8492
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 9864 8508 9916 8560
rect 10416 8551 10468 8560
rect 10416 8517 10425 8551
rect 10425 8517 10459 8551
rect 10459 8517 10468 8551
rect 10416 8508 10468 8517
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 11152 8440 11204 8492
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 11796 8440 11848 8492
rect 12716 8440 12768 8492
rect 9864 8372 9916 8424
rect 10784 8415 10836 8424
rect 10784 8381 10793 8415
rect 10793 8381 10827 8415
rect 10827 8381 10836 8415
rect 10784 8372 10836 8381
rect 6460 8279 6512 8288
rect 6460 8245 6469 8279
rect 6469 8245 6503 8279
rect 6503 8245 6512 8279
rect 6460 8236 6512 8245
rect 7472 8236 7524 8288
rect 7840 8236 7892 8288
rect 8852 8236 8904 8288
rect 9312 8279 9364 8288
rect 9312 8245 9321 8279
rect 9321 8245 9355 8279
rect 9355 8245 9364 8279
rect 9312 8236 9364 8245
rect 9956 8236 10008 8288
rect 13360 8279 13412 8288
rect 13360 8245 13369 8279
rect 13369 8245 13403 8279
rect 13403 8245 13412 8279
rect 13360 8236 13412 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 12214 8134 12266 8186
rect 12278 8134 12330 8186
rect 12342 8134 12394 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 1584 8032 1636 8084
rect 1492 7939 1544 7948
rect 1492 7905 1501 7939
rect 1501 7905 1535 7939
rect 1535 7905 1544 7939
rect 1492 7896 1544 7905
rect 1676 7939 1728 7948
rect 1676 7905 1685 7939
rect 1685 7905 1719 7939
rect 1719 7905 1728 7939
rect 1676 7896 1728 7905
rect 4620 8032 4672 8084
rect 8576 8032 8628 8084
rect 9128 8032 9180 8084
rect 9680 8032 9732 8084
rect 9956 8032 10008 8084
rect 10784 8032 10836 8084
rect 3332 7964 3384 8016
rect 4804 7964 4856 8016
rect 5356 8007 5408 8016
rect 5356 7973 5365 8007
rect 5365 7973 5399 8007
rect 5399 7973 5408 8007
rect 5356 7964 5408 7973
rect 3424 7896 3476 7948
rect 4068 7896 4120 7948
rect 4896 7939 4948 7948
rect 3148 7828 3200 7880
rect 3884 7828 3936 7880
rect 4896 7905 4905 7939
rect 4905 7905 4939 7939
rect 4939 7905 4948 7939
rect 4896 7896 4948 7905
rect 6460 7896 6512 7948
rect 6552 7896 6604 7948
rect 13268 8007 13320 8016
rect 13268 7973 13277 8007
rect 13277 7973 13311 8007
rect 13311 7973 13320 8007
rect 13268 7964 13320 7973
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 8024 7896 8076 7948
rect 8668 7939 8720 7948
rect 8668 7905 8677 7939
rect 8677 7905 8711 7939
rect 8711 7905 8720 7939
rect 8668 7896 8720 7905
rect 8852 7896 8904 7948
rect 9772 7896 9824 7948
rect 7932 7828 7984 7880
rect 8944 7828 8996 7880
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 9312 7828 9364 7837
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 10232 7896 10284 7948
rect 10876 7896 10928 7948
rect 10600 7828 10652 7880
rect 1768 7803 1820 7812
rect 1768 7769 1777 7803
rect 1777 7769 1811 7803
rect 1811 7769 1820 7803
rect 1768 7760 1820 7769
rect 3056 7760 3108 7812
rect 6736 7803 6788 7812
rect 6736 7769 6745 7803
rect 6745 7769 6779 7803
rect 6779 7769 6788 7803
rect 6736 7760 6788 7769
rect 4436 7692 4488 7744
rect 5356 7692 5408 7744
rect 7564 7692 7616 7744
rect 8116 7803 8168 7812
rect 8116 7769 8125 7803
rect 8125 7769 8159 7803
rect 8159 7769 8168 7803
rect 8116 7760 8168 7769
rect 9220 7760 9272 7812
rect 8760 7692 8812 7744
rect 8852 7692 8904 7744
rect 9680 7692 9732 7744
rect 9864 7735 9916 7744
rect 9864 7701 9873 7735
rect 9873 7701 9907 7735
rect 9907 7701 9916 7735
rect 9864 7692 9916 7701
rect 10048 7692 10100 7744
rect 10416 7692 10468 7744
rect 12624 7896 12676 7948
rect 13360 7939 13412 7948
rect 13360 7905 13369 7939
rect 13369 7905 13403 7939
rect 13403 7905 13412 7939
rect 13360 7896 13412 7905
rect 11152 7803 11204 7812
rect 11152 7769 11161 7803
rect 11161 7769 11195 7803
rect 11195 7769 11204 7803
rect 11152 7760 11204 7769
rect 11796 7803 11848 7812
rect 11796 7769 11805 7803
rect 11805 7769 11839 7803
rect 11839 7769 11848 7803
rect 11796 7760 11848 7769
rect 12256 7760 12308 7812
rect 13360 7692 13412 7744
rect 8214 7590 8266 7642
rect 8278 7590 8330 7642
rect 8342 7590 8394 7642
rect 8406 7590 8458 7642
rect 8470 7590 8522 7642
rect 3056 7531 3108 7540
rect 3056 7497 3065 7531
rect 3065 7497 3099 7531
rect 3099 7497 3108 7531
rect 3056 7488 3108 7497
rect 3332 7488 3384 7540
rect 6736 7488 6788 7540
rect 5264 7420 5316 7472
rect 3884 7395 3936 7404
rect 1492 7284 1544 7336
rect 3884 7361 3893 7395
rect 3893 7361 3927 7395
rect 3927 7361 3936 7395
rect 3884 7352 3936 7361
rect 4436 7395 4488 7404
rect 4436 7361 4445 7395
rect 4445 7361 4479 7395
rect 4479 7361 4488 7395
rect 4436 7352 4488 7361
rect 5724 7352 5776 7404
rect 7472 7488 7524 7540
rect 8116 7488 8168 7540
rect 10324 7488 10376 7540
rect 10968 7488 11020 7540
rect 11152 7488 11204 7540
rect 12256 7531 12308 7540
rect 12256 7497 12265 7531
rect 12265 7497 12299 7531
rect 12299 7497 12308 7531
rect 12256 7488 12308 7497
rect 7196 7420 7248 7472
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 7656 7352 7708 7404
rect 9220 7420 9272 7472
rect 9956 7420 10008 7472
rect 8392 7395 8444 7404
rect 8392 7361 8401 7395
rect 8401 7361 8435 7395
rect 8435 7361 8444 7395
rect 8576 7395 8628 7404
rect 8392 7352 8444 7361
rect 8576 7361 8585 7395
rect 8585 7361 8619 7395
rect 8619 7361 8628 7395
rect 8576 7352 8628 7361
rect 8852 7395 8904 7404
rect 8852 7361 8855 7395
rect 8855 7361 8904 7395
rect 8852 7352 8904 7361
rect 9036 7352 9088 7404
rect 9404 7352 9456 7404
rect 9864 7395 9916 7404
rect 9864 7361 9873 7395
rect 9873 7361 9907 7395
rect 9907 7361 9916 7395
rect 9864 7352 9916 7361
rect 10508 7420 10560 7472
rect 10232 7352 10284 7404
rect 10876 7352 10928 7404
rect 11796 7352 11848 7404
rect 12900 7352 12952 7404
rect 13360 7395 13412 7404
rect 13360 7361 13369 7395
rect 13369 7361 13403 7395
rect 13403 7361 13412 7395
rect 13360 7352 13412 7361
rect 3148 7216 3200 7268
rect 2596 7148 2648 7200
rect 5356 7216 5408 7268
rect 7012 7259 7064 7268
rect 7012 7225 7021 7259
rect 7021 7225 7055 7259
rect 7055 7225 7064 7259
rect 7012 7216 7064 7225
rect 8944 7284 8996 7336
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 12808 7327 12860 7336
rect 8760 7216 8812 7268
rect 8852 7216 8904 7268
rect 9772 7216 9824 7268
rect 10876 7216 10928 7268
rect 12808 7293 12817 7327
rect 12817 7293 12851 7327
rect 12851 7293 12860 7327
rect 12808 7284 12860 7293
rect 4620 7148 4672 7200
rect 5080 7148 5132 7200
rect 9036 7148 9088 7200
rect 9496 7148 9548 7200
rect 10784 7148 10836 7200
rect 11336 7148 11388 7200
rect 13176 7191 13228 7200
rect 13176 7157 13185 7191
rect 13185 7157 13219 7191
rect 13219 7157 13228 7191
rect 13176 7148 13228 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 12214 7046 12266 7098
rect 12278 7046 12330 7098
rect 12342 7046 12394 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 3884 6987 3936 6996
rect 3884 6953 3893 6987
rect 3893 6953 3927 6987
rect 3927 6953 3936 6987
rect 3884 6944 3936 6953
rect 5080 6987 5132 6996
rect 5080 6953 5110 6987
rect 5110 6953 5132 6987
rect 5080 6944 5132 6953
rect 7196 6944 7248 6996
rect 7288 6944 7340 6996
rect 8668 6944 8720 6996
rect 9864 6944 9916 6996
rect 10416 6944 10468 6996
rect 12624 6944 12676 6996
rect 6920 6876 6972 6928
rect 7564 6876 7616 6928
rect 7932 6876 7984 6928
rect 8392 6876 8444 6928
rect 10048 6919 10100 6928
rect 2596 6783 2648 6792
rect 2596 6749 2605 6783
rect 2605 6749 2639 6783
rect 2639 6749 2648 6783
rect 2596 6740 2648 6749
rect 3424 6740 3476 6792
rect 3700 6740 3752 6792
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4804 6783 4856 6792
rect 4804 6749 4813 6783
rect 4813 6749 4847 6783
rect 4847 6749 4856 6783
rect 4804 6740 4856 6749
rect 6920 6783 6972 6792
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 5816 6672 5868 6724
rect 2780 6647 2832 6656
rect 2780 6613 2789 6647
rect 2789 6613 2823 6647
rect 2823 6613 2832 6647
rect 2780 6604 2832 6613
rect 2964 6604 3016 6656
rect 7564 6783 7616 6792
rect 7564 6749 7568 6783
rect 7568 6749 7602 6783
rect 7602 6749 7616 6783
rect 7564 6740 7616 6749
rect 7748 6808 7800 6860
rect 8116 6740 8168 6792
rect 8576 6808 8628 6860
rect 8760 6851 8812 6860
rect 8760 6817 8769 6851
rect 8769 6817 8803 6851
rect 8803 6817 8812 6851
rect 9404 6851 9456 6860
rect 8760 6808 8812 6817
rect 8852 6740 8904 6792
rect 9404 6817 9413 6851
rect 9413 6817 9447 6851
rect 9447 6817 9456 6851
rect 9404 6808 9456 6817
rect 10048 6885 10057 6919
rect 10057 6885 10091 6919
rect 10091 6885 10100 6919
rect 10048 6876 10100 6885
rect 10232 6876 10284 6928
rect 9036 6740 9088 6792
rect 9404 6672 9456 6724
rect 9496 6672 9548 6724
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 10784 6783 10836 6792
rect 10784 6749 10793 6783
rect 10793 6749 10827 6783
rect 10827 6749 10836 6783
rect 10784 6740 10836 6749
rect 11336 6740 11388 6792
rect 9220 6604 9272 6656
rect 9680 6604 9732 6656
rect 9956 6604 10008 6656
rect 10232 6604 10284 6656
rect 10784 6604 10836 6656
rect 12808 6808 12860 6860
rect 11612 6740 11664 6792
rect 12348 6740 12400 6792
rect 12624 6740 12676 6792
rect 13176 6783 13228 6792
rect 13176 6749 13185 6783
rect 13185 6749 13219 6783
rect 13219 6749 13228 6783
rect 13176 6740 13228 6749
rect 12256 6604 12308 6656
rect 12716 6647 12768 6656
rect 12716 6613 12725 6647
rect 12725 6613 12759 6647
rect 12759 6613 12768 6647
rect 12716 6604 12768 6613
rect 13268 6647 13320 6656
rect 13268 6613 13277 6647
rect 13277 6613 13311 6647
rect 13311 6613 13320 6647
rect 13268 6604 13320 6613
rect 8214 6502 8266 6554
rect 8278 6502 8330 6554
rect 8342 6502 8394 6554
rect 8406 6502 8458 6554
rect 8470 6502 8522 6554
rect 2780 6400 2832 6452
rect 5816 6443 5868 6452
rect 5816 6409 5825 6443
rect 5825 6409 5859 6443
rect 5859 6409 5868 6443
rect 5816 6400 5868 6409
rect 8116 6443 8168 6452
rect 8116 6409 8125 6443
rect 8125 6409 8159 6443
rect 8159 6409 8168 6443
rect 8116 6400 8168 6409
rect 8576 6400 8628 6452
rect 9496 6400 9548 6452
rect 10048 6400 10100 6452
rect 10232 6400 10284 6452
rect 12348 6400 12400 6452
rect 3884 6307 3936 6316
rect 3884 6273 3893 6307
rect 3893 6273 3927 6307
rect 3927 6273 3936 6307
rect 3884 6264 3936 6273
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 5356 6307 5408 6316
rect 5356 6273 5365 6307
rect 5365 6273 5399 6307
rect 5399 6273 5408 6307
rect 5356 6264 5408 6273
rect 5908 6264 5960 6316
rect 8668 6264 8720 6316
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 9680 6332 9732 6384
rect 10048 6307 10100 6316
rect 10048 6273 10057 6307
rect 10057 6273 10091 6307
rect 10091 6273 10100 6307
rect 10324 6307 10376 6316
rect 10048 6264 10100 6273
rect 10324 6273 10347 6307
rect 10347 6273 10376 6307
rect 10324 6264 10376 6273
rect 12256 6332 12308 6384
rect 12716 6332 12768 6384
rect 10784 6264 10836 6316
rect 1676 6239 1728 6248
rect 1676 6205 1685 6239
rect 1685 6205 1719 6239
rect 1719 6205 1728 6239
rect 1676 6196 1728 6205
rect 3240 6196 3292 6248
rect 3056 6128 3108 6180
rect 3424 6103 3476 6112
rect 3424 6069 3433 6103
rect 3433 6069 3467 6103
rect 3467 6069 3476 6103
rect 3424 6060 3476 6069
rect 3976 6060 4028 6112
rect 4804 6196 4856 6248
rect 7012 6196 7064 6248
rect 7656 6196 7708 6248
rect 9496 6196 9548 6248
rect 9680 6196 9732 6248
rect 8944 6171 8996 6180
rect 8944 6137 8953 6171
rect 8953 6137 8987 6171
rect 8987 6137 8996 6171
rect 8944 6128 8996 6137
rect 9036 6128 9088 6180
rect 5172 6103 5224 6112
rect 5172 6069 5181 6103
rect 5181 6069 5215 6103
rect 5215 6069 5224 6103
rect 5172 6060 5224 6069
rect 8852 6060 8904 6112
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 10048 6060 10100 6069
rect 11152 6103 11204 6112
rect 11152 6069 11161 6103
rect 11161 6069 11195 6103
rect 11195 6069 11204 6103
rect 11152 6060 11204 6069
rect 11704 6239 11756 6248
rect 11704 6205 11713 6239
rect 11713 6205 11747 6239
rect 11747 6205 11756 6239
rect 11704 6196 11756 6205
rect 12624 6060 12676 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 12214 5958 12266 6010
rect 12278 5958 12330 6010
rect 12342 5958 12394 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 2964 5856 3016 5908
rect 3608 5856 3660 5908
rect 7656 5899 7708 5908
rect 7656 5865 7665 5899
rect 7665 5865 7699 5899
rect 7699 5865 7708 5899
rect 7656 5856 7708 5865
rect 8668 5899 8720 5908
rect 8668 5865 8677 5899
rect 8677 5865 8711 5899
rect 8711 5865 8720 5899
rect 8668 5856 8720 5865
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 2044 5695 2096 5704
rect 2044 5661 2053 5695
rect 2053 5661 2087 5695
rect 2087 5661 2096 5695
rect 7196 5720 7248 5772
rect 7840 5720 7892 5772
rect 8576 5720 8628 5772
rect 8852 5720 8904 5772
rect 2044 5652 2096 5661
rect 1676 5516 1728 5568
rect 1952 5516 2004 5568
rect 2964 5652 3016 5704
rect 3056 5695 3108 5704
rect 3056 5661 3065 5695
rect 3065 5661 3099 5695
rect 3099 5661 3108 5695
rect 3056 5652 3108 5661
rect 3332 5627 3384 5636
rect 3332 5593 3341 5627
rect 3341 5593 3375 5627
rect 3375 5593 3384 5627
rect 3332 5584 3384 5593
rect 3516 5627 3568 5636
rect 3516 5593 3525 5627
rect 3525 5593 3559 5627
rect 3559 5593 3568 5627
rect 3516 5584 3568 5593
rect 7472 5652 7524 5704
rect 4160 5627 4212 5636
rect 4160 5593 4169 5627
rect 4169 5593 4203 5627
rect 4203 5593 4212 5627
rect 4160 5584 4212 5593
rect 5172 5584 5224 5636
rect 2964 5516 3016 5568
rect 3884 5516 3936 5568
rect 3976 5516 4028 5568
rect 5080 5516 5132 5568
rect 8300 5652 8352 5704
rect 8760 5652 8812 5704
rect 8944 5695 8996 5704
rect 8944 5661 8953 5695
rect 8953 5661 8987 5695
rect 8987 5661 8996 5695
rect 8944 5652 8996 5661
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 10416 5856 10468 5908
rect 13360 5856 13412 5908
rect 10048 5763 10100 5772
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 10048 5720 10100 5729
rect 8944 5516 8996 5568
rect 9588 5559 9640 5568
rect 9588 5525 9597 5559
rect 9597 5525 9631 5559
rect 9631 5525 9640 5559
rect 9588 5516 9640 5525
rect 11152 5652 11204 5704
rect 11704 5695 11756 5704
rect 11704 5661 11713 5695
rect 11713 5661 11747 5695
rect 11747 5661 11756 5695
rect 11704 5652 11756 5661
rect 11520 5516 11572 5568
rect 11980 5627 12032 5636
rect 11980 5593 11989 5627
rect 11989 5593 12023 5627
rect 12023 5593 12032 5627
rect 11980 5584 12032 5593
rect 12716 5584 12768 5636
rect 8214 5414 8266 5466
rect 8278 5414 8330 5466
rect 8342 5414 8394 5466
rect 8406 5414 8458 5466
rect 8470 5414 8522 5466
rect 1952 5355 2004 5364
rect 1952 5321 1961 5355
rect 1961 5321 1995 5355
rect 1995 5321 2004 5355
rect 1952 5312 2004 5321
rect 3608 5312 3660 5364
rect 4160 5355 4212 5364
rect 4160 5321 4169 5355
rect 4169 5321 4203 5355
rect 4203 5321 4212 5355
rect 4160 5312 4212 5321
rect 2964 5287 3016 5296
rect 2964 5253 2973 5287
rect 2973 5253 3007 5287
rect 3007 5253 3016 5287
rect 2964 5244 3016 5253
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 2044 5219 2096 5228
rect 2044 5185 2054 5219
rect 2054 5185 2088 5219
rect 2088 5185 2096 5219
rect 2044 5176 2096 5185
rect 2780 5108 2832 5160
rect 3056 5219 3108 5228
rect 3056 5185 3065 5219
rect 3065 5185 3099 5219
rect 3099 5185 3108 5219
rect 3056 5176 3108 5185
rect 3608 5219 3660 5228
rect 3608 5185 3612 5219
rect 3612 5185 3646 5219
rect 3646 5185 3660 5219
rect 3608 5176 3660 5185
rect 3424 5108 3476 5160
rect 3884 5176 3936 5228
rect 4436 5219 4488 5228
rect 3332 5040 3384 5092
rect 4436 5185 4445 5219
rect 4445 5185 4479 5219
rect 4479 5185 4488 5219
rect 4436 5176 4488 5185
rect 4068 5151 4120 5160
rect 4068 5117 4077 5151
rect 4077 5117 4111 5151
rect 4111 5117 4120 5151
rect 5632 5312 5684 5364
rect 5448 5244 5500 5296
rect 11980 5312 12032 5364
rect 12716 5355 12768 5364
rect 12716 5321 12725 5355
rect 12725 5321 12759 5355
rect 12759 5321 12768 5355
rect 12716 5312 12768 5321
rect 5172 5219 5224 5228
rect 5172 5185 5180 5219
rect 5180 5185 5214 5219
rect 5214 5185 5224 5219
rect 5172 5176 5224 5185
rect 5540 5219 5592 5228
rect 5540 5185 5549 5219
rect 5549 5185 5583 5219
rect 5583 5185 5592 5219
rect 5540 5176 5592 5185
rect 4068 5108 4120 5117
rect 5172 5040 5224 5092
rect 5356 5151 5408 5160
rect 5356 5117 5365 5151
rect 5365 5117 5399 5151
rect 5399 5117 5408 5151
rect 6828 5176 6880 5228
rect 8300 5219 8352 5228
rect 8300 5185 8309 5219
rect 8309 5185 8343 5219
rect 8343 5185 8352 5219
rect 8300 5176 8352 5185
rect 8760 5219 8812 5228
rect 8760 5185 8769 5219
rect 8769 5185 8803 5219
rect 8803 5185 8812 5219
rect 8760 5176 8812 5185
rect 8944 5219 8996 5228
rect 8944 5185 8953 5219
rect 8953 5185 8987 5219
rect 8987 5185 8996 5219
rect 8944 5176 8996 5185
rect 9588 5244 9640 5296
rect 9404 5176 9456 5228
rect 10416 5244 10468 5296
rect 10784 5287 10836 5296
rect 10784 5253 10793 5287
rect 10793 5253 10827 5287
rect 10827 5253 10836 5287
rect 10784 5244 10836 5253
rect 10876 5244 10928 5296
rect 10140 5176 10192 5228
rect 11612 5176 11664 5228
rect 12624 5176 12676 5228
rect 5356 5108 5408 5117
rect 2412 4972 2464 5024
rect 3240 4972 3292 5024
rect 3608 4972 3660 5024
rect 5448 4972 5500 5024
rect 7472 4972 7524 5024
rect 9864 5108 9916 5160
rect 10692 5108 10744 5160
rect 9220 5040 9272 5092
rect 8392 5015 8444 5024
rect 8392 4981 8401 5015
rect 8401 4981 8435 5015
rect 8435 4981 8444 5015
rect 8392 4972 8444 4981
rect 10048 4972 10100 5024
rect 10416 4972 10468 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 12214 4870 12266 4922
rect 12278 4870 12330 4922
rect 12342 4870 12394 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 2780 4768 2832 4820
rect 3516 4768 3568 4820
rect 4896 4768 4948 4820
rect 5908 4768 5960 4820
rect 6828 4768 6880 4820
rect 8944 4768 8996 4820
rect 9404 4768 9456 4820
rect 10232 4768 10284 4820
rect 1400 4700 1452 4752
rect 2320 4675 2372 4684
rect 2320 4641 2329 4675
rect 2329 4641 2363 4675
rect 2363 4641 2372 4675
rect 2320 4632 2372 4641
rect 3516 4675 3568 4684
rect 3516 4641 3525 4675
rect 3525 4641 3559 4675
rect 3559 4641 3568 4675
rect 3516 4632 3568 4641
rect 4712 4700 4764 4752
rect 5172 4700 5224 4752
rect 6000 4700 6052 4752
rect 8300 4700 8352 4752
rect 10048 4743 10100 4752
rect 10048 4709 10057 4743
rect 10057 4709 10091 4743
rect 10091 4709 10100 4743
rect 10048 4700 10100 4709
rect 1584 4564 1636 4616
rect 1860 4564 1912 4616
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 3976 4632 4028 4684
rect 4344 4632 4396 4684
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 3884 4564 3936 4616
rect 5816 4632 5868 4684
rect 8392 4632 8444 4684
rect 2964 4496 3016 4548
rect 5632 4607 5684 4616
rect 5632 4573 5641 4607
rect 5641 4573 5675 4607
rect 5675 4573 5684 4607
rect 5908 4607 5960 4616
rect 5632 4564 5684 4573
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 6276 4564 6328 4616
rect 5264 4539 5316 4548
rect 2136 4428 2188 4480
rect 3976 4428 4028 4480
rect 4620 4428 4672 4480
rect 5264 4505 5273 4539
rect 5273 4505 5307 4539
rect 5307 4505 5316 4539
rect 5264 4496 5316 4505
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 7196 4607 7248 4616
rect 6552 4564 6604 4573
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7196 4564 7248 4573
rect 8116 4564 8168 4616
rect 9496 4607 9548 4616
rect 5540 4428 5592 4480
rect 5632 4428 5684 4480
rect 6644 4496 6696 4548
rect 7380 4539 7432 4548
rect 7380 4505 7389 4539
rect 7389 4505 7423 4539
rect 7423 4505 7432 4539
rect 7380 4496 7432 4505
rect 8760 4496 8812 4548
rect 9496 4573 9505 4607
rect 9505 4573 9539 4607
rect 9539 4573 9548 4607
rect 9496 4564 9548 4573
rect 9864 4607 9916 4616
rect 9864 4573 9873 4607
rect 9873 4573 9907 4607
rect 9907 4573 9916 4607
rect 9864 4564 9916 4573
rect 10784 4632 10836 4684
rect 10140 4607 10192 4616
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 10692 4607 10744 4616
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 11796 4632 11848 4684
rect 11612 4607 11664 4616
rect 6460 4428 6512 4480
rect 6552 4428 6604 4480
rect 7564 4428 7616 4480
rect 8852 4428 8904 4480
rect 9220 4428 9272 4480
rect 11060 4496 11112 4548
rect 9588 4428 9640 4480
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 11428 4496 11480 4548
rect 8214 4326 8266 4378
rect 8278 4326 8330 4378
rect 8342 4326 8394 4378
rect 8406 4326 8458 4378
rect 8470 4326 8522 4378
rect 3884 4267 3936 4276
rect 3884 4233 3893 4267
rect 3893 4233 3927 4267
rect 3927 4233 3936 4267
rect 3884 4224 3936 4233
rect 3516 4199 3568 4208
rect 3516 4165 3525 4199
rect 3525 4165 3559 4199
rect 3559 4165 3568 4199
rect 3516 4156 3568 4165
rect 3976 4199 4028 4208
rect 3976 4165 3985 4199
rect 3985 4165 4019 4199
rect 4019 4165 4028 4199
rect 3976 4156 4028 4165
rect 4620 4199 4672 4208
rect 4620 4165 4629 4199
rect 4629 4165 4663 4199
rect 4663 4165 4672 4199
rect 4620 4156 4672 4165
rect 5632 4156 5684 4208
rect 1676 4088 1728 4140
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 2320 4131 2372 4140
rect 2320 4097 2329 4131
rect 2329 4097 2363 4131
rect 2363 4097 2372 4131
rect 2320 4088 2372 4097
rect 2596 4131 2648 4140
rect 2596 4097 2605 4131
rect 2605 4097 2639 4131
rect 2639 4097 2648 4131
rect 2596 4088 2648 4097
rect 3056 4131 3108 4140
rect 3056 4097 3065 4131
rect 3065 4097 3099 4131
rect 3099 4097 3108 4131
rect 3056 4088 3108 4097
rect 2044 4063 2096 4072
rect 2044 4029 2053 4063
rect 2053 4029 2087 4063
rect 2087 4029 2096 4063
rect 3792 4088 3844 4140
rect 7380 4224 7432 4276
rect 8116 4224 8168 4276
rect 8852 4156 8904 4208
rect 9496 4224 9548 4276
rect 10140 4224 10192 4276
rect 10508 4224 10560 4276
rect 2044 4020 2096 4029
rect 3976 4020 4028 4072
rect 4344 4063 4396 4072
rect 4344 4029 4353 4063
rect 4353 4029 4387 4063
rect 4387 4029 4396 4063
rect 4344 4020 4396 4029
rect 6460 4131 6512 4140
rect 6460 4097 6469 4131
rect 6469 4097 6503 4131
rect 6503 4097 6512 4131
rect 6460 4088 6512 4097
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6644 4088 6696 4097
rect 6828 4131 6880 4140
rect 6828 4097 6842 4131
rect 6842 4097 6876 4131
rect 6876 4097 6880 4131
rect 7380 4131 7432 4140
rect 6828 4088 6880 4097
rect 7380 4097 7389 4131
rect 7389 4097 7423 4131
rect 7423 4097 7432 4131
rect 7380 4088 7432 4097
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 10324 4131 10376 4140
rect 10324 4097 10334 4131
rect 10334 4097 10368 4131
rect 10368 4097 10376 4131
rect 10692 4224 10744 4276
rect 11796 4199 11848 4208
rect 11796 4165 11805 4199
rect 11805 4165 11839 4199
rect 11839 4165 11848 4199
rect 11796 4156 11848 4165
rect 12808 4156 12860 4208
rect 10324 4088 10376 4097
rect 3792 3884 3844 3936
rect 6736 3952 6788 4004
rect 7472 4020 7524 4072
rect 8116 4063 8168 4072
rect 8116 4029 8125 4063
rect 8125 4029 8159 4063
rect 8159 4029 8168 4063
rect 8116 4020 8168 4029
rect 6184 3884 6236 3936
rect 6644 3884 6696 3936
rect 6920 3884 6972 3936
rect 7656 3884 7708 3936
rect 10232 4063 10284 4072
rect 10232 4029 10241 4063
rect 10241 4029 10275 4063
rect 10275 4029 10284 4063
rect 10968 4131 11020 4140
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 11520 4131 11572 4140
rect 10232 4020 10284 4029
rect 10784 4020 10836 4072
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 10968 3952 11020 4004
rect 11612 3884 11664 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 12214 3782 12266 3834
rect 12278 3782 12330 3834
rect 12342 3782 12394 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 1768 3476 1820 3528
rect 2964 3680 3016 3732
rect 2044 3612 2096 3664
rect 2136 3544 2188 3596
rect 2228 3519 2280 3528
rect 2228 3485 2237 3519
rect 2237 3485 2271 3519
rect 2271 3485 2280 3519
rect 2228 3476 2280 3485
rect 2412 3476 2464 3528
rect 2688 3519 2740 3528
rect 2688 3485 2697 3519
rect 2697 3485 2731 3519
rect 2731 3485 2740 3519
rect 2688 3476 2740 3485
rect 2504 3408 2556 3460
rect 3056 3476 3108 3528
rect 3976 3680 4028 3732
rect 4620 3680 4672 3732
rect 5632 3680 5684 3732
rect 5908 3544 5960 3596
rect 7472 3680 7524 3732
rect 8116 3680 8168 3732
rect 9496 3680 9548 3732
rect 6920 3587 6972 3596
rect 6920 3553 6929 3587
rect 6929 3553 6963 3587
rect 6963 3553 6972 3587
rect 6920 3544 6972 3553
rect 7380 3544 7432 3596
rect 9404 3544 9456 3596
rect 10232 3680 10284 3732
rect 12808 3680 12860 3732
rect 10968 3544 11020 3596
rect 3608 3476 3660 3528
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 9864 3476 9916 3528
rect 9956 3476 10008 3528
rect 12624 3476 12676 3528
rect 3884 3408 3936 3460
rect 4068 3408 4120 3460
rect 4896 3408 4948 3460
rect 5448 3408 5500 3460
rect 6828 3408 6880 3460
rect 7656 3408 7708 3460
rect 9588 3408 9640 3460
rect 10416 3408 10468 3460
rect 11888 3408 11940 3460
rect 2596 3340 2648 3392
rect 4712 3340 4764 3392
rect 5264 3340 5316 3392
rect 6552 3340 6604 3392
rect 11980 3383 12032 3392
rect 11980 3349 11989 3383
rect 11989 3349 12023 3383
rect 12023 3349 12032 3383
rect 11980 3340 12032 3349
rect 12992 3340 13044 3392
rect 8214 3238 8266 3290
rect 8278 3238 8330 3290
rect 8342 3238 8394 3290
rect 8406 3238 8458 3290
rect 8470 3238 8522 3290
rect 2596 3136 2648 3188
rect 4712 3179 4764 3188
rect 4712 3145 4721 3179
rect 4721 3145 4755 3179
rect 4755 3145 4764 3179
rect 4712 3136 4764 3145
rect 5356 3136 5408 3188
rect 6736 3136 6788 3188
rect 10508 3136 10560 3188
rect 1676 3068 1728 3120
rect 1584 3043 1636 3052
rect 1584 3009 1593 3043
rect 1593 3009 1627 3043
rect 1627 3009 1636 3043
rect 1584 3000 1636 3009
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 2504 3000 2556 3052
rect 3056 3043 3108 3052
rect 3056 3009 3065 3043
rect 3065 3009 3099 3043
rect 3099 3009 3108 3043
rect 3056 3000 3108 3009
rect 4068 3000 4120 3052
rect 2044 2932 2096 2984
rect 6552 3068 6604 3120
rect 7288 3111 7340 3120
rect 7288 3077 7297 3111
rect 7297 3077 7331 3111
rect 7331 3077 7340 3111
rect 7288 3068 7340 3077
rect 8668 3068 8720 3120
rect 5080 3043 5132 3052
rect 5080 3009 5089 3043
rect 5089 3009 5123 3043
rect 5123 3009 5132 3043
rect 5080 3000 5132 3009
rect 5816 3043 5868 3052
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 5816 3000 5868 3009
rect 6000 3000 6052 3052
rect 6736 3043 6788 3052
rect 6736 3009 6745 3043
rect 6745 3009 6779 3043
rect 6779 3009 6788 3043
rect 6736 3000 6788 3009
rect 4988 2932 5040 2984
rect 5264 2932 5316 2984
rect 6092 2975 6144 2984
rect 6092 2941 6101 2975
rect 6101 2941 6135 2975
rect 6135 2941 6144 2975
rect 6092 2932 6144 2941
rect 6920 2932 6972 2984
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 7564 3043 7616 3052
rect 7564 3009 7573 3043
rect 7573 3009 7607 3043
rect 7607 3009 7616 3043
rect 9956 3068 10008 3120
rect 11980 3136 12032 3188
rect 12992 3068 13044 3120
rect 7564 3000 7616 3009
rect 9864 3043 9916 3052
rect 9864 3009 9873 3043
rect 9873 3009 9907 3043
rect 9907 3009 9916 3043
rect 9864 3000 9916 3009
rect 9404 2975 9456 2984
rect 9404 2941 9413 2975
rect 9413 2941 9447 2975
rect 9447 2941 9456 2975
rect 9404 2932 9456 2941
rect 10232 3000 10284 3052
rect 10692 3000 10744 3052
rect 10876 3043 10928 3052
rect 10876 3009 10885 3043
rect 10885 3009 10919 3043
rect 10919 3009 10928 3043
rect 10876 3000 10928 3009
rect 10968 3000 11020 3052
rect 11520 3000 11572 3052
rect 11152 2932 11204 2984
rect 12716 2932 12768 2984
rect 5724 2864 5776 2916
rect 7012 2907 7064 2916
rect 7012 2873 7021 2907
rect 7021 2873 7055 2907
rect 7055 2873 7064 2907
rect 7012 2864 7064 2873
rect 7932 2907 7984 2916
rect 7932 2873 7941 2907
rect 7941 2873 7975 2907
rect 7975 2873 7984 2907
rect 7932 2864 7984 2873
rect 9680 2864 9732 2916
rect 10232 2864 10284 2916
rect 10416 2907 10468 2916
rect 10416 2873 10425 2907
rect 10425 2873 10459 2907
rect 10459 2873 10468 2907
rect 10416 2864 10468 2873
rect 1676 2796 1728 2848
rect 3792 2796 3844 2848
rect 3976 2839 4028 2848
rect 3976 2805 3985 2839
rect 3985 2805 4019 2839
rect 4019 2805 4028 2839
rect 3976 2796 4028 2805
rect 6460 2796 6512 2848
rect 13452 2839 13504 2848
rect 13452 2805 13461 2839
rect 13461 2805 13495 2839
rect 13495 2805 13504 2839
rect 13452 2796 13504 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 12214 2694 12266 2746
rect 12278 2694 12330 2746
rect 12342 2694 12394 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 2964 2635 3016 2644
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 1768 2388 1820 2440
rect 2412 2567 2464 2576
rect 2412 2533 2421 2567
rect 2421 2533 2455 2567
rect 2455 2533 2464 2567
rect 2412 2524 2464 2533
rect 2964 2601 2973 2635
rect 2973 2601 3007 2635
rect 3007 2601 3016 2635
rect 2964 2592 3016 2601
rect 3976 2592 4028 2644
rect 4804 2592 4856 2644
rect 5632 2592 5684 2644
rect 7288 2592 7340 2644
rect 7564 2635 7616 2644
rect 3056 2524 3108 2576
rect 3148 2524 3200 2576
rect 4896 2524 4948 2576
rect 5080 2567 5132 2576
rect 5080 2533 5089 2567
rect 5089 2533 5123 2567
rect 5123 2533 5132 2567
rect 5080 2524 5132 2533
rect 7564 2601 7573 2635
rect 7573 2601 7607 2635
rect 7607 2601 7616 2635
rect 7564 2592 7616 2601
rect 8668 2592 8720 2644
rect 9404 2592 9456 2644
rect 11888 2635 11940 2644
rect 11888 2601 11897 2635
rect 11897 2601 11931 2635
rect 11931 2601 11940 2635
rect 11888 2592 11940 2601
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 1584 2320 1636 2372
rect 2504 2388 2556 2440
rect 4068 2456 4120 2508
rect 5448 2499 5500 2508
rect 5448 2465 5457 2499
rect 5457 2465 5491 2499
rect 5491 2465 5500 2499
rect 5448 2456 5500 2465
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 5540 2431 5592 2440
rect 5540 2397 5549 2431
rect 5549 2397 5583 2431
rect 5583 2397 5592 2431
rect 5540 2388 5592 2397
rect 5632 2388 5684 2440
rect 3516 2363 3568 2372
rect 3516 2329 3525 2363
rect 3525 2329 3559 2363
rect 3559 2329 3568 2363
rect 3516 2320 3568 2329
rect 2044 2252 2096 2304
rect 4252 2295 4304 2304
rect 4252 2261 4261 2295
rect 4261 2261 4295 2295
rect 4295 2261 4304 2295
rect 4252 2252 4304 2261
rect 4896 2363 4948 2372
rect 4896 2329 4905 2363
rect 4905 2329 4939 2363
rect 4939 2329 4948 2363
rect 4896 2320 4948 2329
rect 6000 2456 6052 2508
rect 6920 2456 6972 2508
rect 7380 2456 7432 2508
rect 6276 2431 6328 2440
rect 6276 2397 6285 2431
rect 6285 2397 6319 2431
rect 6319 2397 6328 2431
rect 6276 2388 6328 2397
rect 7564 2388 7616 2440
rect 7932 2524 7984 2576
rect 8116 2388 8168 2440
rect 6184 2320 6236 2372
rect 8760 2431 8812 2440
rect 8760 2397 8769 2431
rect 8769 2397 8803 2431
rect 8803 2397 8812 2431
rect 8760 2388 8812 2397
rect 9864 2456 9916 2508
rect 9588 2431 9640 2440
rect 9588 2397 9597 2431
rect 9597 2397 9631 2431
rect 9631 2397 9640 2431
rect 9588 2388 9640 2397
rect 9956 2431 10008 2440
rect 9404 2363 9456 2372
rect 9404 2329 9413 2363
rect 9413 2329 9447 2363
rect 9447 2329 9456 2363
rect 9404 2320 9456 2329
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 11520 2388 11572 2440
rect 12624 2388 12676 2440
rect 12716 2388 12768 2440
rect 13452 2456 13504 2508
rect 9864 2320 9916 2372
rect 10232 2363 10284 2372
rect 10232 2329 10241 2363
rect 10241 2329 10275 2363
rect 10275 2329 10284 2363
rect 10232 2320 10284 2329
rect 13452 2320 13504 2372
rect 11060 2252 11112 2304
rect 11152 2252 11204 2304
rect 12624 2252 12676 2304
rect 8214 2150 8266 2202
rect 8278 2150 8330 2202
rect 8342 2150 8394 2202
rect 8406 2150 8458 2202
rect 8470 2150 8522 2202
rect 1584 2048 1636 2100
rect 2872 1980 2924 2032
rect 3516 2048 3568 2100
rect 8116 2091 8168 2100
rect 3792 1912 3844 1964
rect 1584 1887 1636 1896
rect 1584 1853 1593 1887
rect 1593 1853 1627 1887
rect 1627 1853 1636 1887
rect 1584 1844 1636 1853
rect 3332 1844 3384 1896
rect 4252 1912 4304 1964
rect 5264 1980 5316 2032
rect 5724 2023 5776 2032
rect 5724 1989 5733 2023
rect 5733 1989 5767 2023
rect 5767 1989 5776 2023
rect 5724 1980 5776 1989
rect 6000 1887 6052 1896
rect 4068 1708 4120 1760
rect 6000 1853 6009 1887
rect 6009 1853 6043 1887
rect 6043 1853 6052 1887
rect 7380 1980 7432 2032
rect 8116 2057 8125 2091
rect 8125 2057 8159 2091
rect 8159 2057 8168 2091
rect 8116 2048 8168 2057
rect 9956 2048 10008 2100
rect 10232 2048 10284 2100
rect 11060 2091 11112 2100
rect 11060 2057 11069 2091
rect 11069 2057 11103 2091
rect 11103 2057 11112 2091
rect 11060 2048 11112 2057
rect 9404 1980 9456 2032
rect 11152 1980 11204 2032
rect 11336 1980 11388 2032
rect 10968 1955 11020 1964
rect 6000 1844 6052 1853
rect 6644 1887 6696 1896
rect 6644 1853 6653 1887
rect 6653 1853 6687 1887
rect 6687 1853 6696 1887
rect 6644 1844 6696 1853
rect 8668 1887 8720 1896
rect 8668 1853 8677 1887
rect 8677 1853 8711 1887
rect 8711 1853 8720 1887
rect 8668 1844 8720 1853
rect 9864 1844 9916 1896
rect 10140 1887 10192 1896
rect 10140 1853 10149 1887
rect 10149 1853 10183 1887
rect 10183 1853 10192 1887
rect 10968 1921 10977 1955
rect 10977 1921 11011 1955
rect 11011 1921 11020 1955
rect 10968 1912 11020 1921
rect 11244 1955 11296 1964
rect 11244 1921 11253 1955
rect 11253 1921 11287 1955
rect 11287 1921 11296 1955
rect 11244 1912 11296 1921
rect 10140 1844 10192 1853
rect 10876 1844 10928 1896
rect 11520 1887 11572 1896
rect 9956 1776 10008 1828
rect 11520 1853 11529 1887
rect 11529 1853 11563 1887
rect 11563 1853 11572 1887
rect 11520 1844 11572 1853
rect 11152 1776 11204 1828
rect 4620 1708 4672 1760
rect 5540 1708 5592 1760
rect 9864 1708 9916 1760
rect 11980 1708 12032 1760
rect 4214 1606 4266 1658
rect 4278 1606 4330 1658
rect 4342 1606 4394 1658
rect 4406 1606 4458 1658
rect 4470 1606 4522 1658
rect 12214 1606 12266 1658
rect 12278 1606 12330 1658
rect 12342 1606 12394 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 2872 1504 2924 1556
rect 3332 1504 3384 1556
rect 3976 1504 4028 1556
rect 1584 1300 1636 1352
rect 3148 1300 3200 1352
rect 4252 1436 4304 1488
rect 4620 1436 4672 1488
rect 4988 1504 5040 1556
rect 5356 1547 5408 1556
rect 5356 1513 5365 1547
rect 5365 1513 5399 1547
rect 5399 1513 5408 1547
rect 5356 1504 5408 1513
rect 5448 1504 5500 1556
rect 6644 1547 6696 1556
rect 6644 1513 6653 1547
rect 6653 1513 6687 1547
rect 6687 1513 6696 1547
rect 6644 1504 6696 1513
rect 7380 1504 7432 1556
rect 9404 1504 9456 1556
rect 11336 1547 11388 1556
rect 11336 1513 11345 1547
rect 11345 1513 11379 1547
rect 11379 1513 11388 1547
rect 11336 1504 11388 1513
rect 13452 1547 13504 1556
rect 13452 1513 13461 1547
rect 13461 1513 13495 1547
rect 13495 1513 13504 1547
rect 13452 1504 13504 1513
rect 5540 1436 5592 1488
rect 8668 1436 8720 1488
rect 9220 1436 9272 1488
rect 10140 1436 10192 1488
rect 3884 1368 3936 1420
rect 3976 1343 4028 1352
rect 3976 1309 4025 1343
rect 4025 1309 4028 1343
rect 3976 1300 4028 1309
rect 4160 1343 4212 1352
rect 4160 1309 4169 1343
rect 4169 1309 4203 1343
rect 4203 1309 4212 1343
rect 4896 1368 4948 1420
rect 4160 1300 4212 1309
rect 5448 1343 5500 1352
rect 5448 1309 5457 1343
rect 5457 1309 5491 1343
rect 5491 1309 5500 1343
rect 5448 1300 5500 1309
rect 5632 1368 5684 1420
rect 5816 1343 5868 1352
rect 5816 1309 5825 1343
rect 5825 1309 5859 1343
rect 5859 1309 5868 1343
rect 5816 1300 5868 1309
rect 6276 1300 6328 1352
rect 6552 1343 6604 1352
rect 6552 1309 6561 1343
rect 6561 1309 6595 1343
rect 6595 1309 6604 1343
rect 6552 1300 6604 1309
rect 4252 1275 4304 1284
rect 4252 1241 4261 1275
rect 4261 1241 4295 1275
rect 4295 1241 4304 1275
rect 8760 1300 8812 1352
rect 11244 1368 11296 1420
rect 11520 1368 11572 1420
rect 11980 1411 12032 1420
rect 11980 1377 11989 1411
rect 11989 1377 12023 1411
rect 12023 1377 12032 1411
rect 11980 1368 12032 1377
rect 4252 1232 4304 1241
rect 9220 1232 9272 1284
rect 1584 1207 1636 1216
rect 1584 1173 1593 1207
rect 1593 1173 1627 1207
rect 1627 1173 1636 1207
rect 1584 1164 1636 1173
rect 3792 1164 3844 1216
rect 5264 1164 5316 1216
rect 12624 1232 12676 1284
rect 9680 1164 9732 1216
rect 8214 1062 8266 1114
rect 8278 1062 8330 1114
rect 8342 1062 8394 1114
rect 8406 1062 8458 1114
rect 8470 1062 8522 1114
<< metal2 >>
rect 570 14200 626 15000
rect 1674 14200 1730 15000
rect 2870 14200 2926 15000
rect 3882 14512 3938 14521
rect 3882 14447 3938 14456
rect 584 13734 612 14200
rect 572 13728 624 13734
rect 572 13670 624 13676
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 12850 1440 13262
rect 1688 12986 1716 14200
rect 2884 13376 2912 14200
rect 2884 13348 3004 13376
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 11898 1440 12786
rect 2148 12238 2176 13262
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 2872 13252 2924 13258
rect 2872 13194 2924 13200
rect 2792 12918 2820 13194
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2884 12238 2912 13194
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 1400 11892 1452 11898
rect 1400 11834 1452 11840
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 1860 11688 1912 11694
rect 1858 11656 1860 11665
rect 2228 11688 2280 11694
rect 1912 11656 1914 11665
rect 1492 11620 1544 11626
rect 2228 11630 2280 11636
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 1858 11591 1914 11600
rect 1492 11562 1544 11568
rect 1504 10606 1532 11562
rect 2240 11150 2268 11630
rect 2792 11354 2820 11630
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2240 10810 2268 11086
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 1674 10704 1730 10713
rect 2884 10674 2912 11698
rect 2976 11014 3004 13348
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 3344 12850 3372 13262
rect 3620 12850 3648 13262
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3344 12442 3372 12786
rect 3620 12442 3648 12786
rect 3896 12646 3924 14447
rect 3974 14200 4030 15000
rect 5170 14200 5226 15000
rect 6274 14200 6330 15000
rect 7470 14200 7526 15000
rect 8574 14200 8630 15000
rect 9770 14200 9826 15000
rect 10874 14200 10930 15000
rect 12070 14200 12126 15000
rect 13174 14200 13230 15000
rect 14370 14200 14426 15000
rect 3988 13802 4016 14200
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 3974 13560 4030 13569
rect 4214 13552 4522 13572
rect 3974 13495 4030 13504
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3344 12238 3372 12378
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3988 12186 4016 13495
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 4804 13252 4856 13258
rect 4804 13194 4856 13200
rect 4816 12714 4844 13194
rect 5092 12850 5120 13262
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4066 12608 4122 12617
rect 4066 12543 4122 12552
rect 4080 12434 4108 12543
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4080 12406 4200 12434
rect 4172 12306 4200 12406
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 3240 12164 3292 12170
rect 3988 12158 4200 12186
rect 3240 12106 3292 12112
rect 3252 11830 3280 12106
rect 4172 11898 4200 12158
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 3240 11824 3292 11830
rect 3240 11766 3292 11772
rect 3252 11286 3280 11766
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3332 11620 3384 11626
rect 3332 11562 3384 11568
rect 3240 11280 3292 11286
rect 3240 11222 3292 11228
rect 3344 11150 3372 11562
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 3068 10674 3096 11086
rect 3344 10742 3372 11086
rect 3436 10810 3464 11630
rect 3896 11218 3924 11834
rect 4356 11694 4384 12242
rect 4816 12238 4844 12650
rect 5184 12434 5212 14200
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5828 12918 5856 13262
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5092 12406 5212 12434
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4908 11558 4936 12038
rect 4988 11620 5040 11626
rect 4988 11562 5040 11568
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3988 11150 4016 11494
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4908 11150 4936 11494
rect 5000 11286 5028 11562
rect 4988 11280 5040 11286
rect 4988 11222 5040 11228
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3332 10736 3384 10742
rect 3332 10678 3384 10684
rect 4540 10674 4568 11086
rect 1674 10639 1676 10648
rect 1728 10639 1730 10648
rect 2872 10668 2924 10674
rect 1676 10610 1728 10616
rect 2872 10610 2924 10616
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1504 9722 1532 10542
rect 3068 10266 3096 10610
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 1766 9752 1822 9761
rect 1492 9716 1544 9722
rect 1766 9687 1822 9696
rect 1492 9658 1544 9664
rect 1504 9042 1532 9658
rect 1780 9042 1808 9687
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2240 9178 2268 9522
rect 2976 9450 3004 9930
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2976 9110 3004 9386
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 1492 9036 1544 9042
rect 1492 8978 1544 8984
rect 1768 9036 1820 9042
rect 1768 8978 1820 8984
rect 1504 7993 1532 8978
rect 3252 8974 3280 9862
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 3344 9110 3372 9590
rect 3896 9586 3924 9998
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3804 9042 3832 9318
rect 3896 9110 3924 9522
rect 4620 9444 4672 9450
rect 4620 9386 4672 9392
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 4632 9042 4660 9386
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 1674 8800 1730 8809
rect 1674 8735 1730 8744
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1596 8090 1624 8434
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1490 7984 1546 7993
rect 1688 7954 1716 8735
rect 3160 8566 3188 8842
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3148 8560 3200 8566
rect 3148 8502 3200 8508
rect 1490 7919 1492 7928
rect 1544 7919 1546 7928
rect 1676 7948 1728 7954
rect 1492 7890 1544 7896
rect 1676 7890 1728 7896
rect 1504 7342 1532 7890
rect 3160 7886 3188 8502
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3344 8022 3372 8434
rect 3332 8016 3384 8022
rect 3332 7958 3384 7964
rect 3148 7880 3200 7886
rect 1766 7848 1822 7857
rect 3148 7822 3200 7828
rect 1766 7783 1768 7792
rect 1820 7783 1822 7792
rect 3056 7812 3108 7818
rect 1768 7754 1820 7760
rect 3056 7754 3108 7760
rect 3068 7546 3096 7754
rect 3344 7546 3372 7958
rect 3436 7954 3464 8774
rect 3620 8566 3648 8910
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4172 8378 4200 8434
rect 4080 8350 4200 8378
rect 4080 7954 4108 8350
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4632 8090 4660 8434
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4816 8022 4844 8774
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 4908 7954 4936 9862
rect 5092 9654 5120 12406
rect 5736 12306 5764 12582
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5276 11694 5304 11834
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5184 10810 5212 11630
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5264 11280 5316 11286
rect 5264 11222 5316 11228
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 10062 5212 10406
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3896 7410 3924 7822
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4448 7410 4476 7686
rect 5276 7478 5304 11222
rect 5368 10742 5396 11562
rect 5644 11354 5672 11698
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5356 10736 5408 10742
rect 5356 10678 5408 10684
rect 5460 10130 5488 11018
rect 5736 10266 5764 12106
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 5828 10810 5856 11630
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5920 11150 5948 11494
rect 6104 11150 6132 11562
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5920 10690 5948 11086
rect 5828 10674 5948 10690
rect 5816 10668 5948 10674
rect 5868 10662 5948 10668
rect 6000 10668 6052 10674
rect 5816 10610 5868 10616
rect 6104 10656 6132 11086
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6052 10628 6132 10656
rect 6000 10610 6052 10616
rect 5828 10470 5856 10610
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5460 9518 5488 10066
rect 5920 10062 5948 10474
rect 6012 10266 6040 10610
rect 6196 10554 6224 10746
rect 6104 10538 6224 10554
rect 6092 10532 6224 10538
rect 6144 10526 6224 10532
rect 6092 10474 6144 10480
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6104 10130 6132 10474
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 6196 10062 6224 10406
rect 6288 10198 6316 14200
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7208 13394 7236 13670
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 6368 13252 6420 13258
rect 6368 13194 6420 13200
rect 6380 12986 6408 13194
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6932 12782 6960 13330
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6932 12442 6960 12718
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6368 12096 6420 12102
rect 6368 12038 6420 12044
rect 6380 10742 6408 12038
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6472 11218 6500 11698
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6368 10736 6420 10742
rect 6368 10678 6420 10684
rect 6472 10690 6500 11154
rect 6644 10736 6696 10742
rect 6472 10684 6644 10690
rect 6472 10678 6696 10684
rect 6472 10674 6684 10678
rect 6460 10668 6684 10674
rect 6512 10662 6684 10668
rect 6460 10610 6512 10616
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6196 9722 6224 9998
rect 6748 9994 6776 11494
rect 6828 11280 6880 11286
rect 6828 11222 6880 11228
rect 6840 10470 6868 11222
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6748 9586 6776 9930
rect 6840 9586 6868 10406
rect 6932 10266 6960 11018
rect 7024 10538 7052 12786
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7116 11354 7144 11698
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 7116 10266 7144 10610
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7208 10198 7236 10610
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 6748 8974 6776 9522
rect 6932 9382 6960 9658
rect 7024 9382 7052 10066
rect 7104 10056 7156 10062
rect 7156 10016 7236 10044
rect 7104 9998 7156 10004
rect 7208 9586 7236 10016
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6932 9110 6960 9318
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 7024 8906 7052 9318
rect 7208 9042 7236 9522
rect 7300 9110 7328 13126
rect 7484 12434 7512 14200
rect 7564 13796 7616 13802
rect 7564 13738 7616 13744
rect 7392 12406 7512 12434
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 5368 8362 5396 8842
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5368 8022 5396 8298
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 5368 7750 5396 7958
rect 5736 7886 5764 8434
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6472 7954 6500 8230
rect 6564 7954 6592 8434
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 5736 7410 5764 7822
rect 6736 7812 6788 7818
rect 6736 7754 6788 7760
rect 6748 7546 6776 7754
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 7208 7478 7236 8774
rect 7392 8634 7420 12406
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7484 11762 7512 12174
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7484 11150 7512 11698
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7576 10674 7604 13738
rect 8024 13388 8076 13394
rect 8024 13330 8076 13336
rect 8036 12850 8064 13330
rect 8214 13084 8522 13104
rect 8214 13082 8220 13084
rect 8276 13082 8300 13084
rect 8356 13082 8380 13084
rect 8436 13082 8460 13084
rect 8516 13082 8522 13084
rect 8276 13030 8278 13082
rect 8458 13030 8460 13082
rect 8214 13028 8220 13030
rect 8276 13028 8300 13030
rect 8356 13028 8380 13030
rect 8436 13028 8460 13030
rect 8516 13028 8522 13030
rect 8214 13008 8522 13028
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 7760 12374 7788 12786
rect 8588 12434 8616 14200
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9416 12782 9444 13194
rect 9692 12850 9720 13262
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9692 12442 9720 12786
rect 9680 12436 9732 12442
rect 8588 12406 8708 12434
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8214 11996 8522 12016
rect 8214 11994 8220 11996
rect 8276 11994 8300 11996
rect 8356 11994 8380 11996
rect 8436 11994 8460 11996
rect 8516 11994 8522 11996
rect 8276 11942 8278 11994
rect 8458 11942 8460 11994
rect 8214 11940 8220 11942
rect 8276 11940 8300 11942
rect 8356 11940 8380 11942
rect 8436 11940 8460 11942
rect 8516 11940 8522 11942
rect 8214 11920 8522 11940
rect 8588 11830 8616 12038
rect 8576 11824 8628 11830
rect 8576 11766 8628 11772
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8312 11354 8340 11630
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7760 10606 7788 10678
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7576 10418 7604 10474
rect 7576 10390 7696 10418
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7484 9625 7512 10202
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7470 9616 7526 9625
rect 7576 9586 7604 9998
rect 7668 9994 7696 10390
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7668 9722 7696 9930
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 7470 9551 7526 9560
rect 7564 9580 7616 9586
rect 7484 8974 7512 9551
rect 7564 9522 7616 9528
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7484 8634 7512 8774
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7576 8430 7604 9046
rect 7668 8888 7696 9658
rect 7760 9382 7788 10542
rect 7852 10538 7880 11154
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8214 10908 8522 10928
rect 8214 10906 8220 10908
rect 8276 10906 8300 10908
rect 8356 10906 8380 10908
rect 8436 10906 8460 10908
rect 8516 10906 8522 10908
rect 8276 10854 8278 10906
rect 8458 10854 8460 10906
rect 8214 10852 8220 10854
rect 8276 10852 8300 10854
rect 8356 10852 8380 10854
rect 8436 10852 8460 10854
rect 8516 10852 8522 10854
rect 8214 10832 8522 10852
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7852 10062 7880 10474
rect 8496 10470 8524 10610
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7748 8900 7800 8906
rect 7668 8860 7748 8888
rect 7748 8842 7800 8848
rect 7760 8566 7788 8842
rect 7748 8560 7800 8566
rect 7748 8502 7800 8508
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7484 8294 7512 8366
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7760 8106 7788 8502
rect 7852 8294 7880 9998
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 8036 9450 8064 9862
rect 8024 9444 8076 9450
rect 8024 9386 8076 9392
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7944 8634 7972 9318
rect 8128 9178 8156 10134
rect 8214 9820 8522 9840
rect 8214 9818 8220 9820
rect 8276 9818 8300 9820
rect 8356 9818 8380 9820
rect 8436 9818 8460 9820
rect 8516 9818 8522 9820
rect 8276 9766 8278 9818
rect 8458 9766 8460 9818
rect 8214 9764 8220 9766
rect 8276 9764 8300 9766
rect 8356 9764 8380 9766
rect 8436 9764 8460 9766
rect 8516 9764 8522 9766
rect 8214 9744 8522 9764
rect 8208 9648 8260 9654
rect 8482 9616 8538 9625
rect 8260 9596 8340 9602
rect 8208 9590 8340 9596
rect 8220 9574 8340 9590
rect 8312 9178 8340 9574
rect 8482 9551 8484 9560
rect 8536 9551 8538 9560
rect 8484 9522 8536 9528
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 8036 8634 8064 8842
rect 8214 8732 8522 8752
rect 8214 8730 8220 8732
rect 8276 8730 8300 8732
rect 8356 8730 8380 8732
rect 8436 8730 8460 8732
rect 8516 8730 8522 8732
rect 8276 8678 8278 8730
rect 8458 8678 8460 8730
rect 8214 8676 8220 8678
rect 8276 8676 8300 8678
rect 8356 8676 8380 8678
rect 8436 8676 8460 8678
rect 8516 8676 8522 8678
rect 8214 8656 8522 8676
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7944 8498 7972 8570
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7760 8078 7880 8106
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7196 7472 7248 7478
rect 7196 7414 7248 7420
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2608 6798 2636 7142
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2792 6458 2820 6598
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 1676 6248 1728 6254
rect 1674 6216 1676 6225
rect 1728 6216 1730 6225
rect 1674 6151 1730 6160
rect 1674 6080 1730 6089
rect 1674 6015 1730 6024
rect 1688 5710 1716 6015
rect 2976 5914 3004 6598
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2976 5710 3004 5850
rect 3068 5710 3096 6122
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1412 4758 1440 5170
rect 1596 5137 1624 5170
rect 1582 5128 1638 5137
rect 1582 5063 1638 5072
rect 1400 4752 1452 4758
rect 1400 4694 1452 4700
rect 1596 4622 1624 5063
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1688 4146 1716 5510
rect 1964 5370 1992 5510
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 2056 5234 2084 5646
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2976 5302 3004 5510
rect 2964 5296 3016 5302
rect 3068 5273 3096 5646
rect 2964 5238 3016 5244
rect 3054 5264 3110 5273
rect 2044 5228 2096 5234
rect 3054 5199 3056 5208
rect 2044 5170 2096 5176
rect 3108 5199 3110 5208
rect 3056 5170 3108 5176
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 1860 4616 1912 4622
rect 1780 4576 1860 4604
rect 1780 4185 1808 4576
rect 1860 4558 1912 4564
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 1766 4176 1822 4185
rect 1676 4140 1728 4146
rect 2148 4146 2176 4422
rect 2332 4146 2360 4626
rect 2424 4622 2452 4966
rect 2792 4826 2820 5102
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2412 4616 2464 4622
rect 2464 4576 2544 4604
rect 2412 4558 2464 4564
rect 1766 4111 1822 4120
rect 2136 4140 2188 4146
rect 1676 4082 1728 4088
rect 1582 3224 1638 3233
rect 1582 3159 1638 3168
rect 1596 3058 1624 3159
rect 1688 3126 1716 4082
rect 1780 3534 1808 4111
rect 2136 4082 2188 4088
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2044 4072 2096 4078
rect 2332 4026 2360 4082
rect 2044 4014 2096 4020
rect 2056 3670 2084 4014
rect 2240 3998 2360 4026
rect 2044 3664 2096 3670
rect 2044 3606 2096 3612
rect 2136 3596 2188 3602
rect 2136 3538 2188 3544
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 1676 3120 1728 3126
rect 1676 3062 1728 3068
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 1596 2378 1624 2994
rect 2044 2984 2096 2990
rect 2148 2972 2176 3538
rect 2240 3534 2268 3998
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2424 3058 2452 3470
rect 2516 3466 2544 4576
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2504 3460 2556 3466
rect 2504 3402 2556 3408
rect 2608 3398 2636 4082
rect 2976 3738 3004 4490
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 2608 3194 2636 3334
rect 2700 3233 2728 3470
rect 2686 3224 2742 3233
rect 2596 3188 2648 3194
rect 2686 3159 2742 3168
rect 2596 3130 2648 3136
rect 2502 3088 2558 3097
rect 2412 3052 2464 3058
rect 2502 3023 2504 3032
rect 2412 2994 2464 3000
rect 2556 3023 2558 3032
rect 2504 2994 2556 3000
rect 2096 2944 2176 2972
rect 2044 2926 2096 2932
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1688 2446 1716 2790
rect 2056 2446 2084 2926
rect 2424 2582 2452 2994
rect 2412 2576 2464 2582
rect 2412 2518 2464 2524
rect 2516 2446 2544 2994
rect 2976 2650 3004 3674
rect 3068 3534 3096 4082
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3068 2582 3096 2994
rect 3160 2774 3188 7210
rect 3896 7002 3924 7346
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 3974 7032 4030 7041
rect 3884 6996 3936 7002
rect 4214 7024 4522 7044
rect 3974 6967 4030 6976
rect 3884 6938 3936 6944
rect 3988 6798 4016 6967
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3252 5030 3280 6190
rect 3436 6118 3464 6734
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3344 5098 3372 5578
rect 3436 5166 3464 6054
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3528 4826 3556 5578
rect 3620 5370 3648 5850
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3620 5030 3648 5170
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 3528 4214 3556 4626
rect 3516 4208 3568 4214
rect 3516 4150 3568 4156
rect 3620 3534 3648 4966
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 3160 2746 3280 2774
rect 3056 2576 3108 2582
rect 3056 2518 3108 2524
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 1584 2372 1636 2378
rect 1584 2314 1636 2320
rect 1780 2281 1808 2382
rect 2056 2310 2084 2382
rect 2044 2304 2096 2310
rect 1766 2272 1822 2281
rect 2044 2246 2096 2252
rect 1766 2207 1822 2216
rect 1584 2100 1636 2106
rect 1584 2042 1636 2048
rect 1596 1902 1624 2042
rect 2872 2032 2924 2038
rect 2872 1974 2924 1980
rect 1584 1896 1636 1902
rect 1584 1838 1636 1844
rect 1596 1358 1624 1838
rect 2884 1562 2912 1974
rect 2872 1556 2924 1562
rect 2872 1498 2924 1504
rect 3160 1358 3188 2518
rect 1584 1352 1636 1358
rect 1584 1294 1636 1300
rect 3148 1352 3200 1358
rect 3252 1329 3280 2746
rect 3516 2372 3568 2378
rect 3516 2314 3568 2320
rect 3528 2106 3556 2314
rect 3516 2100 3568 2106
rect 3516 2042 3568 2048
rect 3332 1896 3384 1902
rect 3332 1838 3384 1844
rect 3344 1562 3372 1838
rect 3332 1556 3384 1562
rect 3332 1498 3384 1504
rect 3148 1294 3200 1300
rect 3238 1320 3294 1329
rect 3238 1255 3294 1264
rect 1584 1216 1636 1222
rect 1584 1158 1636 1164
rect 1596 513 1624 1158
rect 3712 800 3740 6734
rect 4632 6322 4660 7142
rect 5092 7002 5120 7142
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 3896 5574 3924 6258
rect 4816 6254 4844 6734
rect 5368 6322 5396 7210
rect 6920 6928 6972 6934
rect 6920 6870 6972 6876
rect 6932 6798 6960 6870
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5828 6458 5856 6666
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 4804 6248 4856 6254
rect 3974 6216 4030 6225
rect 4804 6190 4856 6196
rect 3974 6151 4030 6160
rect 3988 6118 4016 6151
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 3988 5574 4016 6054
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 5184 5642 5212 6054
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 5172 5636 5224 5642
rect 5172 5578 5224 5584
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3896 5234 3924 5510
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3988 4690 4016 5510
rect 4172 5370 4200 5578
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4434 5264 4490 5273
rect 4434 5199 4436 5208
rect 4488 5199 4490 5208
rect 5092 5216 5120 5510
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5172 5228 5224 5234
rect 5092 5188 5172 5216
rect 4436 5170 4488 5176
rect 5172 5170 5224 5176
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 3804 4146 3832 4558
rect 3896 4282 3924 4558
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 3988 4214 4016 4422
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3988 4078 4016 4150
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3804 2854 3832 3878
rect 3988 3738 4016 4014
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 4080 3466 4108 5102
rect 5184 5098 5212 5170
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4356 4078 4384 4626
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4632 4214 4660 4422
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4356 3924 4384 4014
rect 4356 3896 4660 3924
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4632 3738 4660 3896
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4724 3618 4752 4694
rect 4632 3590 4752 3618
rect 3884 3460 3936 3466
rect 3884 3402 3936 3408
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3804 1970 3832 2382
rect 3792 1964 3844 1970
rect 3792 1906 3844 1912
rect 3804 1222 3832 1906
rect 3896 1426 3924 3402
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4080 2961 4108 2994
rect 4066 2952 4122 2961
rect 4066 2887 4122 2896
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 3988 2650 4016 2790
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 4080 2514 4108 2887
rect 4632 2774 4660 3590
rect 4908 3466 4936 4762
rect 5184 4758 5212 5034
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 5368 4570 5396 5102
rect 5460 5030 5488 5238
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5276 4554 5396 4570
rect 5264 4548 5396 4554
rect 5316 4542 5396 4548
rect 5264 4490 5316 4496
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4724 3194 4752 3334
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4632 2746 4844 2774
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4816 2650 4844 2746
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 4908 2582 4936 3402
rect 5276 3398 5304 4490
rect 5460 3466 5488 4966
rect 5552 4486 5580 5170
rect 5644 4622 5672 5306
rect 5920 4826 5948 6258
rect 7024 6254 7052 7210
rect 7208 7002 7236 7414
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7300 7002 7328 7346
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6840 4826 6868 5170
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5552 3720 5580 4422
rect 5644 4214 5672 4422
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 5632 3732 5684 3738
rect 5552 3692 5632 3720
rect 5632 3674 5684 3680
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5356 3188 5408 3194
rect 5460 3176 5488 3402
rect 5408 3148 5580 3176
rect 5356 3130 5408 3136
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 4896 2576 4948 2582
rect 4894 2544 4896 2553
rect 4948 2544 4950 2553
rect 4068 2508 4120 2514
rect 4894 2479 4950 2488
rect 4068 2450 4120 2456
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4252 2304 4304 2310
rect 4252 2246 4304 2252
rect 4264 1970 4292 2246
rect 4252 1964 4304 1970
rect 4252 1906 4304 1912
rect 4264 1850 4292 1906
rect 4080 1822 4292 1850
rect 4080 1766 4108 1822
rect 4632 1766 4660 2382
rect 4896 2372 4948 2378
rect 4896 2314 4948 2320
rect 4068 1760 4120 1766
rect 4068 1702 4120 1708
rect 4620 1760 4672 1766
rect 4620 1702 4672 1708
rect 3976 1556 4028 1562
rect 3976 1498 4028 1504
rect 3884 1420 3936 1426
rect 3884 1362 3936 1368
rect 3988 1358 4016 1498
rect 4080 1442 4108 1702
rect 4214 1660 4522 1680
rect 4214 1658 4220 1660
rect 4276 1658 4300 1660
rect 4356 1658 4380 1660
rect 4436 1658 4460 1660
rect 4516 1658 4522 1660
rect 4276 1606 4278 1658
rect 4458 1606 4460 1658
rect 4214 1604 4220 1606
rect 4276 1604 4300 1606
rect 4356 1604 4380 1606
rect 4436 1604 4460 1606
rect 4516 1604 4522 1606
rect 4214 1584 4522 1604
rect 4632 1494 4660 1702
rect 4252 1488 4304 1494
rect 4080 1414 4200 1442
rect 4252 1430 4304 1436
rect 4620 1488 4672 1494
rect 4620 1430 4672 1436
rect 4172 1358 4200 1414
rect 3976 1352 4028 1358
rect 3976 1294 4028 1300
rect 4160 1352 4212 1358
rect 4160 1294 4212 1300
rect 4264 1290 4292 1430
rect 4908 1426 4936 2314
rect 5000 1562 5028 2926
rect 5092 2582 5120 2994
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 5276 2446 5304 2926
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5264 2440 5316 2446
rect 5316 2400 5396 2428
rect 5264 2382 5316 2388
rect 5264 2032 5316 2038
rect 5264 1974 5316 1980
rect 4988 1556 5040 1562
rect 4988 1498 5040 1504
rect 4896 1420 4948 1426
rect 4896 1362 4948 1368
rect 4252 1284 4304 1290
rect 4252 1226 4304 1232
rect 5276 1222 5304 1974
rect 5368 1562 5396 2400
rect 5460 1562 5488 2450
rect 5552 2446 5580 3148
rect 5828 3058 5856 4626
rect 5920 4622 5948 4762
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5644 2446 5672 2586
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5552 1766 5580 2382
rect 5540 1760 5592 1766
rect 5540 1702 5592 1708
rect 5356 1556 5408 1562
rect 5356 1498 5408 1504
rect 5448 1556 5500 1562
rect 5448 1498 5500 1504
rect 5460 1358 5488 1498
rect 5552 1494 5580 1702
rect 5540 1488 5592 1494
rect 5540 1430 5592 1436
rect 5644 1426 5672 2382
rect 5736 2038 5764 2858
rect 5814 2544 5870 2553
rect 5814 2479 5870 2488
rect 5724 2032 5776 2038
rect 5724 1974 5776 1980
rect 5632 1420 5684 1426
rect 5632 1362 5684 1368
rect 5828 1358 5856 2479
rect 5920 1884 5948 3538
rect 6012 3534 6040 4694
rect 7208 4622 7236 5714
rect 7484 5710 7512 7482
rect 7576 6934 7604 7686
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7576 6798 7604 6870
rect 7668 6848 7696 7346
rect 7748 6860 7800 6866
rect 7668 6820 7748 6848
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7668 6254 7696 6820
rect 7748 6802 7800 6808
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7668 5914 7696 6190
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7852 5778 7880 8078
rect 8036 7954 8064 8570
rect 8208 8560 8260 8566
rect 8206 8528 8208 8537
rect 8260 8528 8262 8537
rect 8588 8514 8616 11086
rect 8680 9994 8708 12406
rect 9680 12378 9732 12384
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9232 12170 9260 12242
rect 9220 12164 9272 12170
rect 9220 12106 9272 12112
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8956 11354 8984 11562
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8668 9988 8720 9994
rect 8668 9930 8720 9936
rect 8852 9988 8904 9994
rect 8852 9930 8904 9936
rect 8864 9654 8892 9930
rect 9048 9654 9076 12038
rect 9232 11694 9260 12106
rect 9784 11898 9812 14200
rect 10230 13424 10286 13433
rect 10888 13394 10916 14200
rect 10230 13359 10286 13368
rect 10876 13388 10928 13394
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 10140 13252 10192 13258
rect 10140 13194 10192 13200
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9416 11218 9444 11494
rect 9508 11218 9536 11630
rect 9876 11626 9904 13194
rect 10060 12918 10088 13194
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 10048 12912 10100 12918
rect 10048 12854 10100 12860
rect 9968 12238 9996 12854
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9968 11830 9996 12038
rect 10060 11898 10088 12854
rect 10152 12442 10180 13194
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10244 12306 10272 13359
rect 10876 13330 10928 13336
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 10152 11354 10180 11698
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9876 10606 9904 11086
rect 10048 10668 10100 10674
rect 10152 10656 10180 11290
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10244 10742 10272 11154
rect 10336 11150 10364 11766
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 10100 10628 10180 10656
rect 10048 10610 10100 10616
rect 9680 10600 9732 10606
rect 9864 10600 9916 10606
rect 9732 10560 9812 10588
rect 9680 10542 9732 10548
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9692 10062 9720 10406
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9508 9722 9536 9998
rect 9678 9752 9734 9761
rect 9496 9716 9548 9722
rect 9678 9687 9734 9696
rect 9496 9658 9548 9664
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 9036 9648 9088 9654
rect 9128 9648 9180 9654
rect 9036 9590 9088 9596
rect 9126 9616 9128 9625
rect 9180 9616 9182 9625
rect 9312 9580 9364 9586
rect 9126 9551 9182 9560
rect 9232 9540 9312 9568
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8772 9042 8800 9454
rect 9232 9382 9260 9540
rect 9312 9522 9364 9528
rect 9692 9450 9720 9687
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8588 8486 8708 8514
rect 8206 8463 8262 8472
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7944 6934 7972 7822
rect 7932 6928 7984 6934
rect 7932 6870 7984 6876
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7944 5658 7972 6870
rect 8036 6780 8064 7890
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8128 7546 8156 7754
rect 8214 7644 8522 7664
rect 8214 7642 8220 7644
rect 8276 7642 8300 7644
rect 8356 7642 8380 7644
rect 8436 7642 8460 7644
rect 8516 7642 8522 7644
rect 8276 7590 8278 7642
rect 8458 7590 8460 7642
rect 8214 7588 8220 7590
rect 8276 7588 8300 7590
rect 8356 7588 8380 7590
rect 8436 7588 8460 7590
rect 8516 7588 8522 7590
rect 8214 7568 8522 7588
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8588 7410 8616 8026
rect 8680 7954 8708 8486
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 8404 6934 8432 7346
rect 8680 7002 8708 7890
rect 8772 7750 8800 8978
rect 8956 8566 8984 9114
rect 9036 8900 9088 8906
rect 9140 8888 9168 9114
rect 9692 9110 9720 9386
rect 9784 9110 9812 10560
rect 9864 10542 9916 10548
rect 9876 9994 9904 10542
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9968 10198 9996 10406
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9864 9988 9916 9994
rect 9864 9930 9916 9936
rect 9876 9674 9904 9930
rect 9876 9646 9996 9674
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9088 8860 9168 8888
rect 9036 8842 9088 8848
rect 9140 8634 9168 8860
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 8944 8560 8996 8566
rect 8944 8502 8996 8508
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8864 7954 8892 8230
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8956 7886 8984 8502
rect 9140 8090 9168 8570
rect 9496 8492 9548 8498
rect 9784 8480 9812 9046
rect 9968 8786 9996 9646
rect 10060 9042 10088 10406
rect 10244 9586 10272 10678
rect 10336 9761 10364 10746
rect 10428 10674 10456 11698
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10520 10674 10548 11630
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10322 9752 10378 9761
rect 10428 9722 10456 10610
rect 10520 10146 10548 10610
rect 10612 10266 10640 13126
rect 10980 12306 11008 13262
rect 12084 13258 12112 14200
rect 12214 13628 12522 13648
rect 12214 13626 12220 13628
rect 12276 13626 12300 13628
rect 12356 13626 12380 13628
rect 12436 13626 12460 13628
rect 12516 13626 12522 13628
rect 12276 13574 12278 13626
rect 12458 13574 12460 13626
rect 12214 13572 12220 13574
rect 12276 13572 12300 13574
rect 12356 13572 12380 13574
rect 12436 13572 12460 13574
rect 12516 13572 12522 13574
rect 12214 13552 12522 13572
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11348 12442 11376 12718
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 11532 12238 11560 12582
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10704 10198 10732 10406
rect 10692 10192 10744 10198
rect 10520 10118 10640 10146
rect 10692 10134 10744 10140
rect 10508 10056 10560 10062
rect 10506 10024 10508 10033
rect 10560 10024 10562 10033
rect 10506 9959 10562 9968
rect 10322 9687 10378 9696
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 10152 9178 10180 9386
rect 10244 9178 10272 9522
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 10060 8906 10088 8978
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 9968 8758 10088 8786
rect 9864 8560 9916 8566
rect 9548 8452 9812 8480
rect 9862 8528 9864 8537
rect 9916 8528 9918 8537
rect 9862 8463 9918 8472
rect 9496 8434 9548 8440
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9324 7886 9352 8230
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 8944 7880 8996 7886
rect 8850 7848 8906 7857
rect 8944 7822 8996 7828
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 8850 7783 8906 7792
rect 9220 7812 9272 7818
rect 8864 7750 8892 7783
rect 9220 7754 9272 7760
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8772 7274 8800 7686
rect 9232 7478 9260 7754
rect 9692 7750 9720 8026
rect 9784 7954 9812 8452
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9876 7886 9904 8366
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9968 8090 9996 8230
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9864 7880 9916 7886
rect 9916 7828 9996 7834
rect 9864 7822 9996 7828
rect 9876 7806 9996 7822
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9220 7472 9272 7478
rect 9220 7414 9272 7420
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 8864 7274 8892 7346
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8852 7268 8904 7274
rect 8852 7210 8904 7216
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 8772 6866 8800 7210
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8116 6792 8168 6798
rect 8036 6752 8116 6780
rect 8116 6734 8168 6740
rect 8128 6458 8156 6734
rect 8214 6556 8522 6576
rect 8214 6554 8220 6556
rect 8276 6554 8300 6556
rect 8356 6554 8380 6556
rect 8436 6554 8460 6556
rect 8516 6554 8522 6556
rect 8276 6502 8278 6554
rect 8458 6502 8460 6554
rect 8214 6500 8220 6502
rect 8276 6500 8300 6502
rect 8356 6500 8380 6502
rect 8436 6500 8460 6502
rect 8516 6500 8522 6502
rect 8214 6480 8522 6500
rect 8588 6458 8616 6802
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8588 5778 8616 6394
rect 8864 6322 8892 6734
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8680 5914 8708 6258
rect 8956 6186 8984 7278
rect 9048 7206 9076 7346
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9048 6798 9076 7142
rect 9416 6866 9444 7346
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 9048 6322 9076 6734
rect 9508 6730 9536 7142
rect 9404 6724 9456 6730
rect 9404 6666 9456 6672
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 9036 6180 9088 6186
rect 9036 6122 9088 6128
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8864 5778 8892 6054
rect 9048 5794 9076 6122
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8956 5766 9076 5794
rect 8300 5704 8352 5710
rect 7944 5652 8300 5658
rect 7944 5646 8352 5652
rect 7944 5630 8340 5646
rect 8128 5216 8156 5630
rect 8214 5468 8522 5488
rect 8214 5466 8220 5468
rect 8276 5466 8300 5468
rect 8356 5466 8380 5468
rect 8436 5466 8460 5468
rect 8516 5466 8522 5468
rect 8276 5414 8278 5466
rect 8458 5414 8460 5466
rect 8214 5412 8220 5414
rect 8276 5412 8300 5414
rect 8356 5412 8380 5414
rect 8436 5412 8460 5414
rect 8516 5412 8522 5414
rect 8214 5392 8522 5412
rect 8300 5228 8352 5234
rect 8128 5188 8300 5216
rect 8300 5170 8352 5176
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 6276 4616 6328 4622
rect 6552 4616 6604 4622
rect 6328 4576 6552 4604
rect 6276 4558 6328 4564
rect 6552 4558 6604 4564
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 6564 4486 6592 4558
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 7380 4548 7432 4554
rect 7380 4490 7432 4496
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 6472 4146 6500 4422
rect 6656 4146 6684 4490
rect 7392 4282 7420 4490
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6090 3088 6146 3097
rect 6000 3052 6052 3058
rect 6090 3023 6146 3032
rect 6000 2994 6052 3000
rect 6012 2514 6040 2994
rect 6104 2990 6132 3023
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6196 2378 6224 3878
rect 6472 2854 6500 4082
rect 6656 3942 6684 4082
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6564 3126 6592 3334
rect 6748 3194 6776 3946
rect 6840 3466 6868 4082
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6932 3602 6960 3878
rect 7392 3602 7420 4082
rect 7484 4078 7512 4966
rect 8312 4758 8340 5170
rect 8392 5024 8444 5030
rect 8588 5012 8616 5714
rect 8956 5710 8984 5766
rect 9232 5710 9260 6598
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 8772 5234 8800 5646
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8956 5234 8984 5510
rect 9416 5234 9444 6666
rect 9508 6458 9536 6666
rect 9692 6662 9720 7686
rect 9876 7410 9904 7686
rect 9968 7478 9996 7806
rect 10060 7750 10088 8758
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9956 7336 10008 7342
rect 10008 7296 10088 7324
rect 9956 7278 10008 7284
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9680 6384 9732 6390
rect 9784 6372 9812 7210
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9732 6344 9812 6372
rect 9680 6326 9732 6332
rect 9496 6248 9548 6254
rect 9680 6248 9732 6254
rect 9496 6190 9548 6196
rect 9678 6216 9680 6225
rect 9732 6216 9734 6225
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 8444 4984 8616 5012
rect 8392 4966 8444 4972
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8404 4690 8432 4966
rect 8956 4826 8984 5170
rect 9508 5114 9536 6190
rect 9678 6151 9734 6160
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9600 5302 9628 5510
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9876 5166 9904 6938
rect 10060 6934 10088 7296
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9864 5160 9916 5166
rect 9220 5092 9272 5098
rect 9508 5086 9628 5114
rect 9864 5102 9916 5108
rect 9220 5034 9272 5040
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7576 4146 7604 4422
rect 8128 4282 8156 4558
rect 8760 4548 8812 4554
rect 8760 4490 8812 4496
rect 8214 4380 8522 4400
rect 8214 4378 8220 4380
rect 8276 4378 8300 4380
rect 8356 4378 8380 4380
rect 8436 4378 8460 4380
rect 8516 4378 8522 4380
rect 8276 4326 8278 4378
rect 8458 4326 8460 4378
rect 8214 4324 8220 4326
rect 8276 4324 8300 4326
rect 8356 4324 8380 4326
rect 8436 4324 8460 4326
rect 8516 4324 8522 4326
rect 8214 4304 8522 4324
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 7484 3738 7512 4014
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7668 3466 7696 3878
rect 8128 3738 8156 4014
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 8214 3292 8522 3312
rect 8214 3290 8220 3292
rect 8276 3290 8300 3292
rect 8356 3290 8380 3292
rect 8436 3290 8460 3292
rect 8516 3290 8522 3292
rect 8276 3238 8278 3290
rect 8458 3238 8460 3290
rect 8214 3236 8220 3238
rect 8276 3236 8300 3238
rect 8356 3236 8380 3238
rect 8436 3236 8460 3238
rect 8516 3236 8522 3238
rect 8214 3216 8522 3236
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 6184 2372 6236 2378
rect 6184 2314 6236 2320
rect 6000 1896 6052 1902
rect 5920 1856 6000 1884
rect 6000 1838 6052 1844
rect 6288 1358 6316 2382
rect 6564 1358 6592 3062
rect 6748 3058 6776 3130
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 8668 3120 8720 3126
rect 8668 3062 8720 3068
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 7010 2952 7066 2961
rect 6932 2514 6960 2926
rect 7010 2887 7012 2896
rect 7064 2887 7066 2896
rect 7012 2858 7064 2864
rect 7300 2650 7328 3062
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7392 2514 7420 2994
rect 7576 2650 7604 2994
rect 7932 2916 7984 2922
rect 7932 2858 7984 2864
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 7576 2446 7604 2586
rect 7944 2582 7972 2858
rect 8680 2650 8708 3062
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 7932 2576 7984 2582
rect 7932 2518 7984 2524
rect 8772 2446 8800 4490
rect 9232 4486 9260 5034
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 8864 4214 8892 4422
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 9232 3534 9260 4422
rect 9416 3602 9444 4762
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9508 4282 9536 4558
rect 9600 4486 9628 5086
rect 9876 4622 9904 5102
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9588 4480 9640 4486
rect 9968 4468 9996 6598
rect 10060 6458 10088 6870
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10060 6225 10088 6258
rect 10046 6216 10102 6225
rect 10046 6151 10102 6160
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10060 5778 10088 6054
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 10152 5234 10180 9114
rect 10244 8634 10272 9114
rect 10324 9104 10376 9110
rect 10324 9046 10376 9052
rect 10336 8838 10364 9046
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10428 8566 10456 9658
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10520 8838 10548 9454
rect 10612 8838 10640 10118
rect 10704 8906 10732 10134
rect 10796 9450 10824 11698
rect 11072 11626 11100 12038
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10888 11218 10916 11494
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 11072 11150 11100 11562
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11164 11150 11192 11290
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 10980 10554 11008 10950
rect 11072 10810 11100 10950
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10980 10526 11284 10554
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11164 10266 11192 10406
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 10980 10146 11008 10202
rect 10980 10118 11100 10146
rect 11072 10044 11100 10118
rect 11256 10112 11284 10526
rect 11440 10266 11468 11222
rect 11532 10810 11560 12174
rect 11900 11354 11928 13126
rect 12360 12986 12388 13262
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 12072 12708 12124 12714
rect 12072 12650 12124 12656
rect 12084 12238 12112 12650
rect 12214 12540 12522 12560
rect 12214 12538 12220 12540
rect 12276 12538 12300 12540
rect 12356 12538 12380 12540
rect 12436 12538 12460 12540
rect 12516 12538 12522 12540
rect 12276 12486 12278 12538
rect 12458 12486 12460 12538
rect 12214 12484 12220 12486
rect 12276 12484 12300 12486
rect 12356 12484 12380 12486
rect 12436 12484 12460 12486
rect 12516 12484 12522 12486
rect 12214 12464 12522 12484
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12214 11452 12522 11472
rect 12214 11450 12220 11452
rect 12276 11450 12300 11452
rect 12356 11450 12380 11452
rect 12436 11450 12460 11452
rect 12516 11450 12522 11452
rect 12276 11398 12278 11450
rect 12458 11398 12460 11450
rect 12214 11396 12220 11398
rect 12276 11396 12300 11398
rect 12356 11396 12380 11398
rect 12436 11396 12460 11398
rect 12516 11396 12522 11398
rect 12214 11376 12522 11396
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11978 11248 12034 11257
rect 11978 11183 12034 11192
rect 11992 10810 12020 11183
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 12360 10674 12388 11086
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12636 10606 12664 13330
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12728 12238 12756 12786
rect 12820 12714 12848 13194
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12912 12442 12940 13194
rect 13188 12866 13216 14200
rect 13096 12838 13216 12866
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12820 10674 12848 11222
rect 12912 10742 12940 11494
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 13004 10674 13032 11698
rect 13096 11694 13124 12838
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 13188 12238 13216 12650
rect 14384 12374 14412 14200
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13464 11830 13492 12038
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 13280 10674 13308 11698
rect 13464 11150 13492 11766
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13372 10742 13400 10950
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 11520 10532 11572 10538
rect 11520 10474 11572 10480
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 10980 10016 11100 10044
rect 11164 10084 11284 10112
rect 10874 9752 10930 9761
rect 10874 9687 10930 9696
rect 10888 9586 10916 9687
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10416 8560 10468 8566
rect 10230 8528 10286 8537
rect 10416 8502 10468 8508
rect 10230 8463 10232 8472
rect 10284 8463 10286 8472
rect 10232 8434 10284 8440
rect 10244 7954 10272 8434
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10244 6934 10272 7346
rect 10232 6928 10284 6934
rect 10232 6870 10284 6876
rect 10336 6798 10364 7482
rect 10428 7002 10456 7686
rect 10520 7478 10548 8774
rect 10796 8514 10824 8978
rect 10980 8906 11008 10016
rect 11164 9976 11192 10084
rect 11072 9948 11192 9976
rect 11244 9988 11296 9994
rect 11072 9654 11100 9948
rect 11244 9930 11296 9936
rect 11256 9674 11284 9930
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 11164 9646 11284 9674
rect 11348 9674 11376 9862
rect 11348 9654 11468 9674
rect 11348 9648 11480 9654
rect 11348 9646 11428 9648
rect 11072 8974 11100 9590
rect 11164 9518 11192 9646
rect 11428 9590 11480 9596
rect 11532 9586 11560 10474
rect 12214 10364 12522 10384
rect 12214 10362 12220 10364
rect 12276 10362 12300 10364
rect 12356 10362 12380 10364
rect 12436 10362 12460 10364
rect 12516 10362 12522 10364
rect 12276 10310 12278 10362
rect 12458 10310 12460 10362
rect 12214 10308 12220 10310
rect 12276 10308 12300 10310
rect 12356 10308 12380 10310
rect 12436 10308 12460 10310
rect 12516 10308 12522 10310
rect 12214 10288 12522 10308
rect 12820 10062 12848 10610
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12912 10130 12940 10542
rect 13004 10266 13032 10610
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12544 9586 12572 9862
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 12532 9580 12584 9586
rect 12584 9540 12756 9568
rect 12532 9522 12584 9528
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 11164 9178 11192 9454
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10876 8900 10928 8906
rect 10876 8842 10928 8848
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10704 8486 10824 8514
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10244 6458 10272 6598
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10060 4758 10088 4966
rect 10244 4826 10272 6394
rect 10336 6322 10364 6734
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10336 5930 10364 6258
rect 10336 5914 10456 5930
rect 10336 5908 10468 5914
rect 10336 5902 10416 5908
rect 10416 5850 10468 5856
rect 10416 5296 10468 5302
rect 10416 5238 10468 5244
rect 10428 5030 10456 5238
rect 10416 5024 10468 5030
rect 10336 4984 10416 5012
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 9588 4422 9640 4428
rect 9876 4440 9996 4468
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9508 3738 9536 4218
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9600 3466 9628 4422
rect 9876 3534 9904 4440
rect 10152 4282 10180 4558
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10336 4146 10364 4984
rect 10416 4966 10468 4972
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 10244 3738 10272 4014
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9968 3126 9996 3470
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9416 2650 9444 2926
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 7564 2440 7616 2446
rect 8116 2440 8168 2446
rect 7564 2382 7616 2388
rect 8114 2408 8116 2417
rect 8760 2440 8812 2446
rect 8168 2408 8170 2417
rect 9588 2440 9640 2446
rect 8760 2382 8812 2388
rect 9402 2408 9458 2417
rect 8114 2343 8170 2352
rect 8128 2106 8156 2343
rect 8214 2204 8522 2224
rect 8214 2202 8220 2204
rect 8276 2202 8300 2204
rect 8356 2202 8380 2204
rect 8436 2202 8460 2204
rect 8516 2202 8522 2204
rect 8276 2150 8278 2202
rect 8458 2150 8460 2202
rect 8214 2148 8220 2150
rect 8276 2148 8300 2150
rect 8356 2148 8380 2150
rect 8436 2148 8460 2150
rect 8516 2148 8522 2150
rect 8214 2128 8522 2148
rect 8116 2100 8168 2106
rect 8116 2042 8168 2048
rect 7380 2032 7432 2038
rect 7380 1974 7432 1980
rect 6644 1896 6696 1902
rect 6644 1838 6696 1844
rect 6656 1562 6684 1838
rect 7392 1562 7420 1974
rect 8668 1896 8720 1902
rect 8668 1838 8720 1844
rect 6644 1556 6696 1562
rect 6644 1498 6696 1504
rect 7380 1556 7432 1562
rect 7380 1498 7432 1504
rect 8680 1494 8708 1838
rect 8668 1488 8720 1494
rect 8668 1430 8720 1436
rect 8772 1358 8800 2382
rect 9692 2428 9720 2858
rect 9876 2514 9904 2994
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 9640 2400 9720 2428
rect 9588 2382 9640 2388
rect 9402 2343 9404 2352
rect 9456 2343 9458 2352
rect 9404 2314 9456 2320
rect 9404 2032 9456 2038
rect 9404 1974 9456 1980
rect 9416 1562 9444 1974
rect 9404 1556 9456 1562
rect 9404 1498 9456 1504
rect 9220 1488 9272 1494
rect 9220 1430 9272 1436
rect 5448 1352 5500 1358
rect 5448 1294 5500 1300
rect 5816 1352 5868 1358
rect 5816 1294 5868 1300
rect 6276 1352 6328 1358
rect 6276 1294 6328 1300
rect 6552 1352 6604 1358
rect 6552 1294 6604 1300
rect 8760 1352 8812 1358
rect 8760 1294 8812 1300
rect 9232 1290 9260 1430
rect 9220 1284 9272 1290
rect 9220 1226 9272 1232
rect 9692 1222 9720 2400
rect 9876 2378 9904 2450
rect 9968 2446 9996 3062
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10244 2922 10272 2994
rect 10428 2922 10456 3402
rect 10520 3194 10548 4218
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 10232 2916 10284 2922
rect 10232 2858 10284 2864
rect 10416 2916 10468 2922
rect 10416 2858 10468 2864
rect 10612 2774 10640 7822
rect 10704 6644 10732 8486
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10796 8090 10824 8366
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10888 7954 10916 8842
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 10980 7546 11008 8842
rect 11164 8498 11192 9114
rect 11348 8498 11376 9318
rect 11532 8906 11560 9522
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11624 8974 11652 9454
rect 12214 9276 12522 9296
rect 12214 9274 12220 9276
rect 12276 9274 12300 9276
rect 12356 9274 12380 9276
rect 12436 9274 12460 9276
rect 12516 9274 12522 9276
rect 12276 9222 12278 9274
rect 12458 9222 12460 9274
rect 12214 9220 12220 9222
rect 12276 9220 12300 9222
rect 12356 9220 12380 9222
rect 12436 9220 12460 9222
rect 12516 9220 12522 9222
rect 12214 9200 12522 9220
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 11164 7546 11192 7754
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 10980 7426 11008 7482
rect 10888 7410 11008 7426
rect 10876 7404 11008 7410
rect 10928 7398 11008 7404
rect 10876 7346 10928 7352
rect 10876 7268 10928 7274
rect 10876 7210 10928 7216
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10796 6798 10824 7142
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10784 6656 10836 6662
rect 10704 6616 10784 6644
rect 10784 6598 10836 6604
rect 10784 6316 10836 6322
rect 10888 6304 10916 7210
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11348 6798 11376 7142
rect 11624 6798 11652 8910
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11808 8498 11836 8774
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11808 7818 11836 8434
rect 12214 8188 12522 8208
rect 12214 8186 12220 8188
rect 12276 8186 12300 8188
rect 12356 8186 12380 8188
rect 12436 8186 12460 8188
rect 12516 8186 12522 8188
rect 12276 8134 12278 8186
rect 12458 8134 12460 8186
rect 12214 8132 12220 8134
rect 12276 8132 12300 8134
rect 12356 8132 12380 8134
rect 12436 8132 12460 8134
rect 12516 8132 12522 8134
rect 12214 8112 12522 8132
rect 12636 7954 12664 8910
rect 12728 8906 12756 9540
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12820 9110 12848 9386
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 12912 8956 12940 10066
rect 13082 10024 13138 10033
rect 13082 9959 13084 9968
rect 13136 9959 13138 9968
rect 13084 9930 13136 9936
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 12820 8928 12940 8956
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 12728 8498 12756 8842
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 11808 7410 11836 7754
rect 12268 7546 12296 7754
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 12214 7100 12522 7120
rect 12214 7098 12220 7100
rect 12276 7098 12300 7100
rect 12356 7098 12380 7100
rect 12436 7098 12460 7100
rect 12516 7098 12522 7100
rect 12276 7046 12278 7098
rect 12458 7046 12460 7098
rect 12214 7044 12220 7046
rect 12276 7044 12300 7046
rect 12356 7044 12380 7046
rect 12436 7044 12460 7046
rect 12516 7044 12522 7046
rect 12214 7024 12522 7044
rect 12636 7002 12664 7890
rect 12820 7342 12848 8928
rect 13188 8809 13216 9862
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13280 9042 13308 9318
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13372 8974 13400 9522
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13174 8800 13230 8809
rect 13372 8786 13400 8910
rect 13174 8735 13230 8744
rect 13280 8758 13400 8786
rect 13280 8022 13308 8758
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13268 8016 13320 8022
rect 13268 7958 13320 7964
rect 13372 7954 13400 8230
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13372 7410 13400 7686
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12820 6866 12848 7278
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12268 6390 12296 6598
rect 12360 6458 12388 6734
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 10836 6276 10916 6304
rect 10784 6258 10836 6264
rect 10796 5302 10824 6258
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11164 5710 11192 6054
rect 11716 5710 11744 6190
rect 12636 6118 12664 6734
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12728 6390 12756 6598
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12214 6012 12522 6032
rect 12214 6010 12220 6012
rect 12276 6010 12300 6012
rect 12356 6010 12380 6012
rect 12436 6010 12460 6012
rect 12516 6010 12522 6012
rect 12276 5958 12278 6010
rect 12458 5958 12460 6010
rect 12214 5956 12220 5958
rect 12276 5956 12300 5958
rect 12356 5956 12380 5958
rect 12436 5956 12460 5958
rect 12516 5956 12522 5958
rect 12214 5936 12522 5956
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11980 5636 12032 5642
rect 11980 5578 12032 5584
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 10784 5296 10836 5302
rect 10784 5238 10836 5244
rect 10876 5296 10928 5302
rect 10928 5244 11008 5250
rect 10876 5238 11008 5244
rect 10888 5222 11008 5238
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10704 4622 10732 5102
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10704 4282 10732 4558
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10796 4078 10824 4626
rect 10980 4146 11008 5222
rect 11072 4554 11468 4570
rect 11060 4548 11480 4554
rect 11112 4542 11428 4548
rect 11060 4490 11112 4496
rect 11428 4490 11480 4496
rect 11532 4146 11560 5510
rect 11992 5370 12020 5578
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 12636 5234 12664 6054
rect 12716 5636 12768 5642
rect 12716 5578 12768 5584
rect 12728 5370 12756 5578
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 11624 4622 11652 5170
rect 12214 4924 12522 4944
rect 12214 4922 12220 4924
rect 12276 4922 12300 4924
rect 12356 4922 12380 4924
rect 12436 4922 12460 4924
rect 12516 4922 12522 4924
rect 12276 4870 12278 4922
rect 12458 4870 12460 4922
rect 12214 4868 12220 4870
rect 12276 4868 12300 4870
rect 12356 4868 12380 4870
rect 12436 4868 12460 4870
rect 12516 4868 12522 4870
rect 12214 4848 12522 4868
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10980 4010 11008 4082
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10980 3602 11008 3946
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10704 3148 11008 3176
rect 10704 3058 10732 3148
rect 10980 3058 11008 3148
rect 11532 3058 11560 4082
rect 11624 3942 11652 4558
rect 11808 4214 11836 4626
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 12214 3836 12522 3856
rect 12214 3834 12220 3836
rect 12276 3834 12300 3836
rect 12356 3834 12380 3836
rect 12436 3834 12460 3836
rect 12516 3834 12522 3836
rect 12276 3782 12278 3834
rect 12458 3782 12460 3834
rect 12214 3780 12220 3782
rect 12276 3780 12300 3782
rect 12356 3780 12380 3782
rect 12436 3780 12460 3782
rect 12516 3780 12522 3782
rect 12214 3760 12522 3780
rect 12636 3534 12664 5170
rect 12808 4208 12860 4214
rect 12808 4150 12860 4156
rect 12820 3738 12848 4150
rect 12912 3777 12940 7346
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13188 6798 13216 7142
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13280 6225 13308 6598
rect 13266 6216 13322 6225
rect 13266 6151 13322 6160
rect 13372 5914 13400 7346
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 12898 3768 12954 3777
rect 12808 3732 12860 3738
rect 12898 3703 12954 3712
rect 12808 3674 12860 3680
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 11888 3460 11940 3466
rect 11888 3402 11940 3408
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 10612 2746 10824 2774
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 9864 2372 9916 2378
rect 9864 2314 9916 2320
rect 9876 1902 9904 2314
rect 9968 2106 9996 2382
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 10244 2106 10272 2314
rect 9956 2100 10008 2106
rect 9956 2042 10008 2048
rect 10232 2100 10284 2106
rect 10232 2042 10284 2048
rect 9864 1896 9916 1902
rect 9864 1838 9916 1844
rect 9876 1766 9904 1838
rect 9968 1834 9996 2042
rect 10140 1896 10192 1902
rect 10140 1838 10192 1844
rect 9956 1828 10008 1834
rect 9956 1770 10008 1776
rect 9864 1760 9916 1766
rect 9864 1702 9916 1708
rect 10152 1494 10180 1838
rect 10140 1488 10192 1494
rect 10140 1430 10192 1436
rect 10796 1329 10824 2746
rect 10888 1902 10916 2994
rect 10980 1970 11008 2994
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 11164 2310 11192 2926
rect 11532 2774 11560 2994
rect 11532 2746 11652 2774
rect 11520 2440 11572 2446
rect 11256 2400 11520 2428
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 11072 2106 11100 2246
rect 11060 2100 11112 2106
rect 11060 2042 11112 2048
rect 11164 2038 11192 2246
rect 11152 2032 11204 2038
rect 11152 1974 11204 1980
rect 11256 1970 11284 2400
rect 11520 2382 11572 2388
rect 11624 2292 11652 2746
rect 11900 2650 11928 3402
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11992 3194 12020 3334
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12214 2748 12522 2768
rect 12214 2746 12220 2748
rect 12276 2746 12300 2748
rect 12356 2746 12380 2748
rect 12436 2746 12460 2748
rect 12516 2746 12522 2748
rect 12276 2694 12278 2746
rect 12458 2694 12460 2746
rect 12214 2692 12220 2694
rect 12276 2692 12300 2694
rect 12356 2692 12380 2694
rect 12436 2692 12460 2694
rect 12516 2692 12522 2694
rect 12214 2672 12522 2692
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 12636 2446 12664 3470
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 13004 3126 13032 3334
rect 12992 3120 13044 3126
rect 12992 3062 13044 3068
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12728 2446 12756 2926
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 13464 2514 13492 2790
rect 13452 2508 13504 2514
rect 13452 2450 13504 2456
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 13452 2372 13504 2378
rect 13452 2314 13504 2320
rect 11532 2264 11652 2292
rect 12624 2304 12676 2310
rect 11336 2032 11388 2038
rect 11336 1974 11388 1980
rect 10968 1964 11020 1970
rect 10968 1906 11020 1912
rect 11244 1964 11296 1970
rect 11244 1906 11296 1912
rect 10876 1896 10928 1902
rect 10876 1838 10928 1844
rect 11152 1828 11204 1834
rect 11152 1770 11204 1776
rect 10782 1320 10838 1329
rect 10782 1255 10838 1264
rect 3792 1216 3844 1222
rect 3792 1158 3844 1164
rect 5264 1216 5316 1222
rect 5264 1158 5316 1164
rect 9680 1216 9732 1222
rect 9680 1158 9732 1164
rect 8214 1116 8522 1136
rect 8214 1114 8220 1116
rect 8276 1114 8300 1116
rect 8356 1114 8380 1116
rect 8436 1114 8460 1116
rect 8516 1114 8522 1116
rect 8276 1062 8278 1114
rect 8458 1062 8460 1114
rect 8214 1060 8220 1062
rect 8276 1060 8300 1062
rect 8356 1060 8380 1062
rect 8436 1060 8460 1062
rect 8516 1060 8522 1062
rect 8214 1040 8522 1060
rect 11164 800 11192 1770
rect 11256 1426 11284 1906
rect 11348 1562 11376 1974
rect 11532 1902 11560 2264
rect 12624 2246 12676 2252
rect 11520 1896 11572 1902
rect 11520 1838 11572 1844
rect 11336 1556 11388 1562
rect 11336 1498 11388 1504
rect 11532 1426 11560 1838
rect 11980 1760 12032 1766
rect 11980 1702 12032 1708
rect 11992 1426 12020 1702
rect 12214 1660 12522 1680
rect 12214 1658 12220 1660
rect 12276 1658 12300 1660
rect 12356 1658 12380 1660
rect 12436 1658 12460 1660
rect 12516 1658 12522 1660
rect 12276 1606 12278 1658
rect 12458 1606 12460 1658
rect 12214 1604 12220 1606
rect 12276 1604 12300 1606
rect 12356 1604 12380 1606
rect 12436 1604 12460 1606
rect 12516 1604 12522 1606
rect 12214 1584 12522 1604
rect 11244 1420 11296 1426
rect 11244 1362 11296 1368
rect 11520 1420 11572 1426
rect 11520 1362 11572 1368
rect 11980 1420 12032 1426
rect 11980 1362 12032 1368
rect 12636 1290 12664 2246
rect 13464 1562 13492 2314
rect 13452 1556 13504 1562
rect 13452 1498 13504 1504
rect 12624 1284 12676 1290
rect 12624 1226 12676 1232
rect 1582 504 1638 513
rect 1582 439 1638 448
rect 3698 0 3754 800
rect 11150 0 11206 800
<< via2 >>
rect 3882 14456 3938 14512
rect 1858 11636 1860 11656
rect 1860 11636 1912 11656
rect 1912 11636 1914 11656
rect 1858 11600 1914 11636
rect 1674 10668 1730 10704
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 3974 13504 4030 13560
rect 4066 12552 4122 12608
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 1674 10648 1676 10668
rect 1676 10648 1728 10668
rect 1728 10648 1730 10668
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 1766 9696 1822 9752
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 1674 8744 1730 8800
rect 1490 7948 1546 7984
rect 1490 7928 1492 7948
rect 1492 7928 1544 7948
rect 1544 7928 1546 7948
rect 1766 7812 1822 7848
rect 1766 7792 1768 7812
rect 1768 7792 1820 7812
rect 1820 7792 1822 7812
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 8220 13082 8276 13084
rect 8300 13082 8356 13084
rect 8380 13082 8436 13084
rect 8460 13082 8516 13084
rect 8220 13030 8266 13082
rect 8266 13030 8276 13082
rect 8300 13030 8330 13082
rect 8330 13030 8342 13082
rect 8342 13030 8356 13082
rect 8380 13030 8394 13082
rect 8394 13030 8406 13082
rect 8406 13030 8436 13082
rect 8460 13030 8470 13082
rect 8470 13030 8516 13082
rect 8220 13028 8276 13030
rect 8300 13028 8356 13030
rect 8380 13028 8436 13030
rect 8460 13028 8516 13030
rect 8220 11994 8276 11996
rect 8300 11994 8356 11996
rect 8380 11994 8436 11996
rect 8460 11994 8516 11996
rect 8220 11942 8266 11994
rect 8266 11942 8276 11994
rect 8300 11942 8330 11994
rect 8330 11942 8342 11994
rect 8342 11942 8356 11994
rect 8380 11942 8394 11994
rect 8394 11942 8406 11994
rect 8406 11942 8436 11994
rect 8460 11942 8470 11994
rect 8470 11942 8516 11994
rect 8220 11940 8276 11942
rect 8300 11940 8356 11942
rect 8380 11940 8436 11942
rect 8460 11940 8516 11942
rect 7470 9560 7526 9616
rect 8220 10906 8276 10908
rect 8300 10906 8356 10908
rect 8380 10906 8436 10908
rect 8460 10906 8516 10908
rect 8220 10854 8266 10906
rect 8266 10854 8276 10906
rect 8300 10854 8330 10906
rect 8330 10854 8342 10906
rect 8342 10854 8356 10906
rect 8380 10854 8394 10906
rect 8394 10854 8406 10906
rect 8406 10854 8436 10906
rect 8460 10854 8470 10906
rect 8470 10854 8516 10906
rect 8220 10852 8276 10854
rect 8300 10852 8356 10854
rect 8380 10852 8436 10854
rect 8460 10852 8516 10854
rect 8220 9818 8276 9820
rect 8300 9818 8356 9820
rect 8380 9818 8436 9820
rect 8460 9818 8516 9820
rect 8220 9766 8266 9818
rect 8266 9766 8276 9818
rect 8300 9766 8330 9818
rect 8330 9766 8342 9818
rect 8342 9766 8356 9818
rect 8380 9766 8394 9818
rect 8394 9766 8406 9818
rect 8406 9766 8436 9818
rect 8460 9766 8470 9818
rect 8470 9766 8516 9818
rect 8220 9764 8276 9766
rect 8300 9764 8356 9766
rect 8380 9764 8436 9766
rect 8460 9764 8516 9766
rect 8482 9580 8538 9616
rect 8482 9560 8484 9580
rect 8484 9560 8536 9580
rect 8536 9560 8538 9580
rect 8220 8730 8276 8732
rect 8300 8730 8356 8732
rect 8380 8730 8436 8732
rect 8460 8730 8516 8732
rect 8220 8678 8266 8730
rect 8266 8678 8276 8730
rect 8300 8678 8330 8730
rect 8330 8678 8342 8730
rect 8342 8678 8356 8730
rect 8380 8678 8394 8730
rect 8394 8678 8406 8730
rect 8406 8678 8436 8730
rect 8460 8678 8470 8730
rect 8470 8678 8516 8730
rect 8220 8676 8276 8678
rect 8300 8676 8356 8678
rect 8380 8676 8436 8678
rect 8460 8676 8516 8678
rect 1674 6196 1676 6216
rect 1676 6196 1728 6216
rect 1728 6196 1730 6216
rect 1674 6160 1730 6196
rect 1674 6024 1730 6080
rect 1582 5072 1638 5128
rect 3054 5228 3110 5264
rect 3054 5208 3056 5228
rect 3056 5208 3108 5228
rect 3108 5208 3110 5228
rect 1766 4120 1822 4176
rect 1582 3168 1638 3224
rect 2686 3168 2742 3224
rect 2502 3052 2558 3088
rect 2502 3032 2504 3052
rect 2504 3032 2556 3052
rect 2556 3032 2558 3052
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3974 6976 4030 7032
rect 1766 2216 1822 2272
rect 3238 1264 3294 1320
rect 3974 6160 4030 6216
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4434 5228 4490 5264
rect 4434 5208 4436 5228
rect 4436 5208 4488 5228
rect 4488 5208 4490 5228
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4066 2896 4122 2952
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4894 2524 4896 2544
rect 4896 2524 4948 2544
rect 4948 2524 4950 2544
rect 4894 2488 4950 2524
rect 4220 1658 4276 1660
rect 4300 1658 4356 1660
rect 4380 1658 4436 1660
rect 4460 1658 4516 1660
rect 4220 1606 4266 1658
rect 4266 1606 4276 1658
rect 4300 1606 4330 1658
rect 4330 1606 4342 1658
rect 4342 1606 4356 1658
rect 4380 1606 4394 1658
rect 4394 1606 4406 1658
rect 4406 1606 4436 1658
rect 4460 1606 4470 1658
rect 4470 1606 4516 1658
rect 4220 1604 4276 1606
rect 4300 1604 4356 1606
rect 4380 1604 4436 1606
rect 4460 1604 4516 1606
rect 5814 2488 5870 2544
rect 8206 8508 8208 8528
rect 8208 8508 8260 8528
rect 8260 8508 8262 8528
rect 8206 8472 8262 8508
rect 10230 13368 10286 13424
rect 9678 9696 9734 9752
rect 9126 9596 9128 9616
rect 9128 9596 9180 9616
rect 9180 9596 9182 9616
rect 9126 9560 9182 9596
rect 8220 7642 8276 7644
rect 8300 7642 8356 7644
rect 8380 7642 8436 7644
rect 8460 7642 8516 7644
rect 8220 7590 8266 7642
rect 8266 7590 8276 7642
rect 8300 7590 8330 7642
rect 8330 7590 8342 7642
rect 8342 7590 8356 7642
rect 8380 7590 8394 7642
rect 8394 7590 8406 7642
rect 8406 7590 8436 7642
rect 8460 7590 8470 7642
rect 8470 7590 8516 7642
rect 8220 7588 8276 7590
rect 8300 7588 8356 7590
rect 8380 7588 8436 7590
rect 8460 7588 8516 7590
rect 10322 9696 10378 9752
rect 12220 13626 12276 13628
rect 12300 13626 12356 13628
rect 12380 13626 12436 13628
rect 12460 13626 12516 13628
rect 12220 13574 12266 13626
rect 12266 13574 12276 13626
rect 12300 13574 12330 13626
rect 12330 13574 12342 13626
rect 12342 13574 12356 13626
rect 12380 13574 12394 13626
rect 12394 13574 12406 13626
rect 12406 13574 12436 13626
rect 12460 13574 12470 13626
rect 12470 13574 12516 13626
rect 12220 13572 12276 13574
rect 12300 13572 12356 13574
rect 12380 13572 12436 13574
rect 12460 13572 12516 13574
rect 10506 10004 10508 10024
rect 10508 10004 10560 10024
rect 10560 10004 10562 10024
rect 10506 9968 10562 10004
rect 9862 8508 9864 8528
rect 9864 8508 9916 8528
rect 9916 8508 9918 8528
rect 9862 8472 9918 8508
rect 8850 7792 8906 7848
rect 8220 6554 8276 6556
rect 8300 6554 8356 6556
rect 8380 6554 8436 6556
rect 8460 6554 8516 6556
rect 8220 6502 8266 6554
rect 8266 6502 8276 6554
rect 8300 6502 8330 6554
rect 8330 6502 8342 6554
rect 8342 6502 8356 6554
rect 8380 6502 8394 6554
rect 8394 6502 8406 6554
rect 8406 6502 8436 6554
rect 8460 6502 8470 6554
rect 8470 6502 8516 6554
rect 8220 6500 8276 6502
rect 8300 6500 8356 6502
rect 8380 6500 8436 6502
rect 8460 6500 8516 6502
rect 8220 5466 8276 5468
rect 8300 5466 8356 5468
rect 8380 5466 8436 5468
rect 8460 5466 8516 5468
rect 8220 5414 8266 5466
rect 8266 5414 8276 5466
rect 8300 5414 8330 5466
rect 8330 5414 8342 5466
rect 8342 5414 8356 5466
rect 8380 5414 8394 5466
rect 8394 5414 8406 5466
rect 8406 5414 8436 5466
rect 8460 5414 8470 5466
rect 8470 5414 8516 5466
rect 8220 5412 8276 5414
rect 8300 5412 8356 5414
rect 8380 5412 8436 5414
rect 8460 5412 8516 5414
rect 6090 3032 6146 3088
rect 9678 6196 9680 6216
rect 9680 6196 9732 6216
rect 9732 6196 9734 6216
rect 9678 6160 9734 6196
rect 8220 4378 8276 4380
rect 8300 4378 8356 4380
rect 8380 4378 8436 4380
rect 8460 4378 8516 4380
rect 8220 4326 8266 4378
rect 8266 4326 8276 4378
rect 8300 4326 8330 4378
rect 8330 4326 8342 4378
rect 8342 4326 8356 4378
rect 8380 4326 8394 4378
rect 8394 4326 8406 4378
rect 8406 4326 8436 4378
rect 8460 4326 8470 4378
rect 8470 4326 8516 4378
rect 8220 4324 8276 4326
rect 8300 4324 8356 4326
rect 8380 4324 8436 4326
rect 8460 4324 8516 4326
rect 8220 3290 8276 3292
rect 8300 3290 8356 3292
rect 8380 3290 8436 3292
rect 8460 3290 8516 3292
rect 8220 3238 8266 3290
rect 8266 3238 8276 3290
rect 8300 3238 8330 3290
rect 8330 3238 8342 3290
rect 8342 3238 8356 3290
rect 8380 3238 8394 3290
rect 8394 3238 8406 3290
rect 8406 3238 8436 3290
rect 8460 3238 8470 3290
rect 8470 3238 8516 3290
rect 8220 3236 8276 3238
rect 8300 3236 8356 3238
rect 8380 3236 8436 3238
rect 8460 3236 8516 3238
rect 7010 2916 7066 2952
rect 7010 2896 7012 2916
rect 7012 2896 7064 2916
rect 7064 2896 7066 2916
rect 10046 6160 10102 6216
rect 12220 12538 12276 12540
rect 12300 12538 12356 12540
rect 12380 12538 12436 12540
rect 12460 12538 12516 12540
rect 12220 12486 12266 12538
rect 12266 12486 12276 12538
rect 12300 12486 12330 12538
rect 12330 12486 12342 12538
rect 12342 12486 12356 12538
rect 12380 12486 12394 12538
rect 12394 12486 12406 12538
rect 12406 12486 12436 12538
rect 12460 12486 12470 12538
rect 12470 12486 12516 12538
rect 12220 12484 12276 12486
rect 12300 12484 12356 12486
rect 12380 12484 12436 12486
rect 12460 12484 12516 12486
rect 12220 11450 12276 11452
rect 12300 11450 12356 11452
rect 12380 11450 12436 11452
rect 12460 11450 12516 11452
rect 12220 11398 12266 11450
rect 12266 11398 12276 11450
rect 12300 11398 12330 11450
rect 12330 11398 12342 11450
rect 12342 11398 12356 11450
rect 12380 11398 12394 11450
rect 12394 11398 12406 11450
rect 12406 11398 12436 11450
rect 12460 11398 12470 11450
rect 12470 11398 12516 11450
rect 12220 11396 12276 11398
rect 12300 11396 12356 11398
rect 12380 11396 12436 11398
rect 12460 11396 12516 11398
rect 11978 11192 12034 11248
rect 10874 9696 10930 9752
rect 10230 8492 10286 8528
rect 10230 8472 10232 8492
rect 10232 8472 10284 8492
rect 10284 8472 10286 8492
rect 12220 10362 12276 10364
rect 12300 10362 12356 10364
rect 12380 10362 12436 10364
rect 12460 10362 12516 10364
rect 12220 10310 12266 10362
rect 12266 10310 12276 10362
rect 12300 10310 12330 10362
rect 12330 10310 12342 10362
rect 12342 10310 12356 10362
rect 12380 10310 12394 10362
rect 12394 10310 12406 10362
rect 12406 10310 12436 10362
rect 12460 10310 12470 10362
rect 12470 10310 12516 10362
rect 12220 10308 12276 10310
rect 12300 10308 12356 10310
rect 12380 10308 12436 10310
rect 12460 10308 12516 10310
rect 8114 2388 8116 2408
rect 8116 2388 8168 2408
rect 8168 2388 8170 2408
rect 8114 2352 8170 2388
rect 8220 2202 8276 2204
rect 8300 2202 8356 2204
rect 8380 2202 8436 2204
rect 8460 2202 8516 2204
rect 8220 2150 8266 2202
rect 8266 2150 8276 2202
rect 8300 2150 8330 2202
rect 8330 2150 8342 2202
rect 8342 2150 8356 2202
rect 8380 2150 8394 2202
rect 8394 2150 8406 2202
rect 8406 2150 8436 2202
rect 8460 2150 8470 2202
rect 8470 2150 8516 2202
rect 8220 2148 8276 2150
rect 8300 2148 8356 2150
rect 8380 2148 8436 2150
rect 8460 2148 8516 2150
rect 9402 2372 9458 2408
rect 9402 2352 9404 2372
rect 9404 2352 9456 2372
rect 9456 2352 9458 2372
rect 12220 9274 12276 9276
rect 12300 9274 12356 9276
rect 12380 9274 12436 9276
rect 12460 9274 12516 9276
rect 12220 9222 12266 9274
rect 12266 9222 12276 9274
rect 12300 9222 12330 9274
rect 12330 9222 12342 9274
rect 12342 9222 12356 9274
rect 12380 9222 12394 9274
rect 12394 9222 12406 9274
rect 12406 9222 12436 9274
rect 12460 9222 12470 9274
rect 12470 9222 12516 9274
rect 12220 9220 12276 9222
rect 12300 9220 12356 9222
rect 12380 9220 12436 9222
rect 12460 9220 12516 9222
rect 12220 8186 12276 8188
rect 12300 8186 12356 8188
rect 12380 8186 12436 8188
rect 12460 8186 12516 8188
rect 12220 8134 12266 8186
rect 12266 8134 12276 8186
rect 12300 8134 12330 8186
rect 12330 8134 12342 8186
rect 12342 8134 12356 8186
rect 12380 8134 12394 8186
rect 12394 8134 12406 8186
rect 12406 8134 12436 8186
rect 12460 8134 12470 8186
rect 12470 8134 12516 8186
rect 12220 8132 12276 8134
rect 12300 8132 12356 8134
rect 12380 8132 12436 8134
rect 12460 8132 12516 8134
rect 13082 9988 13138 10024
rect 13082 9968 13084 9988
rect 13084 9968 13136 9988
rect 13136 9968 13138 9988
rect 12220 7098 12276 7100
rect 12300 7098 12356 7100
rect 12380 7098 12436 7100
rect 12460 7098 12516 7100
rect 12220 7046 12266 7098
rect 12266 7046 12276 7098
rect 12300 7046 12330 7098
rect 12330 7046 12342 7098
rect 12342 7046 12356 7098
rect 12380 7046 12394 7098
rect 12394 7046 12406 7098
rect 12406 7046 12436 7098
rect 12460 7046 12470 7098
rect 12470 7046 12516 7098
rect 12220 7044 12276 7046
rect 12300 7044 12356 7046
rect 12380 7044 12436 7046
rect 12460 7044 12516 7046
rect 13174 8744 13230 8800
rect 12220 6010 12276 6012
rect 12300 6010 12356 6012
rect 12380 6010 12436 6012
rect 12460 6010 12516 6012
rect 12220 5958 12266 6010
rect 12266 5958 12276 6010
rect 12300 5958 12330 6010
rect 12330 5958 12342 6010
rect 12342 5958 12356 6010
rect 12380 5958 12394 6010
rect 12394 5958 12406 6010
rect 12406 5958 12436 6010
rect 12460 5958 12470 6010
rect 12470 5958 12516 6010
rect 12220 5956 12276 5958
rect 12300 5956 12356 5958
rect 12380 5956 12436 5958
rect 12460 5956 12516 5958
rect 12220 4922 12276 4924
rect 12300 4922 12356 4924
rect 12380 4922 12436 4924
rect 12460 4922 12516 4924
rect 12220 4870 12266 4922
rect 12266 4870 12276 4922
rect 12300 4870 12330 4922
rect 12330 4870 12342 4922
rect 12342 4870 12356 4922
rect 12380 4870 12394 4922
rect 12394 4870 12406 4922
rect 12406 4870 12436 4922
rect 12460 4870 12470 4922
rect 12470 4870 12516 4922
rect 12220 4868 12276 4870
rect 12300 4868 12356 4870
rect 12380 4868 12436 4870
rect 12460 4868 12516 4870
rect 12220 3834 12276 3836
rect 12300 3834 12356 3836
rect 12380 3834 12436 3836
rect 12460 3834 12516 3836
rect 12220 3782 12266 3834
rect 12266 3782 12276 3834
rect 12300 3782 12330 3834
rect 12330 3782 12342 3834
rect 12342 3782 12356 3834
rect 12380 3782 12394 3834
rect 12394 3782 12406 3834
rect 12406 3782 12436 3834
rect 12460 3782 12470 3834
rect 12470 3782 12516 3834
rect 12220 3780 12276 3782
rect 12300 3780 12356 3782
rect 12380 3780 12436 3782
rect 12460 3780 12516 3782
rect 13266 6160 13322 6216
rect 12898 3712 12954 3768
rect 12220 2746 12276 2748
rect 12300 2746 12356 2748
rect 12380 2746 12436 2748
rect 12460 2746 12516 2748
rect 12220 2694 12266 2746
rect 12266 2694 12276 2746
rect 12300 2694 12330 2746
rect 12330 2694 12342 2746
rect 12342 2694 12356 2746
rect 12380 2694 12394 2746
rect 12394 2694 12406 2746
rect 12406 2694 12436 2746
rect 12460 2694 12470 2746
rect 12470 2694 12516 2746
rect 12220 2692 12276 2694
rect 12300 2692 12356 2694
rect 12380 2692 12436 2694
rect 12460 2692 12516 2694
rect 10782 1264 10838 1320
rect 8220 1114 8276 1116
rect 8300 1114 8356 1116
rect 8380 1114 8436 1116
rect 8460 1114 8516 1116
rect 8220 1062 8266 1114
rect 8266 1062 8276 1114
rect 8300 1062 8330 1114
rect 8330 1062 8342 1114
rect 8342 1062 8356 1114
rect 8380 1062 8394 1114
rect 8394 1062 8406 1114
rect 8406 1062 8436 1114
rect 8460 1062 8470 1114
rect 8470 1062 8516 1114
rect 8220 1060 8276 1062
rect 8300 1060 8356 1062
rect 8380 1060 8436 1062
rect 8460 1060 8516 1062
rect 12220 1658 12276 1660
rect 12300 1658 12356 1660
rect 12380 1658 12436 1660
rect 12460 1658 12516 1660
rect 12220 1606 12266 1658
rect 12266 1606 12276 1658
rect 12300 1606 12330 1658
rect 12330 1606 12342 1658
rect 12342 1606 12356 1658
rect 12380 1606 12394 1658
rect 12394 1606 12406 1658
rect 12406 1606 12436 1658
rect 12460 1606 12470 1658
rect 12470 1606 12516 1658
rect 12220 1604 12276 1606
rect 12300 1604 12356 1606
rect 12380 1604 12436 1606
rect 12460 1604 12516 1606
rect 1582 448 1638 504
<< metal3 >>
rect 0 14514 800 14544
rect 3877 14514 3943 14517
rect 0 14512 3943 14514
rect 0 14456 3882 14512
rect 3938 14456 3943 14512
rect 0 14454 3943 14456
rect 0 14424 800 14454
rect 3877 14451 3943 14454
rect 14200 13698 15000 13728
rect 12758 13638 15000 13698
rect 4208 13632 4528 13633
rect 0 13562 800 13592
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 12208 13632 12528 13633
rect 12208 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12528 13632
rect 12208 13567 12528 13568
rect 3969 13562 4035 13565
rect 0 13560 4035 13562
rect 0 13504 3974 13560
rect 4030 13504 4035 13560
rect 0 13502 4035 13504
rect 0 13472 800 13502
rect 3969 13499 4035 13502
rect 10225 13426 10291 13429
rect 12758 13426 12818 13638
rect 14200 13608 15000 13638
rect 10225 13424 12818 13426
rect 10225 13368 10230 13424
rect 10286 13368 12818 13424
rect 10225 13366 12818 13368
rect 10225 13363 10291 13366
rect 8208 13088 8528 13089
rect 8208 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8528 13088
rect 8208 13023 8528 13024
rect 0 12610 800 12640
rect 4061 12610 4127 12613
rect 0 12608 4127 12610
rect 0 12552 4066 12608
rect 4122 12552 4127 12608
rect 0 12550 4127 12552
rect 0 12520 800 12550
rect 4061 12547 4127 12550
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 12208 12544 12528 12545
rect 12208 12480 12216 12544
rect 12280 12480 12296 12544
rect 12360 12480 12376 12544
rect 12440 12480 12456 12544
rect 12520 12480 12528 12544
rect 12208 12479 12528 12480
rect 8208 12000 8528 12001
rect 8208 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8528 12000
rect 8208 11935 8528 11936
rect 0 11658 800 11688
rect 1853 11658 1919 11661
rect 0 11656 1919 11658
rect 0 11600 1858 11656
rect 1914 11600 1919 11656
rect 0 11598 1919 11600
rect 0 11568 800 11598
rect 1853 11595 1919 11598
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 12208 11456 12528 11457
rect 12208 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12528 11456
rect 12208 11391 12528 11392
rect 11973 11250 12039 11253
rect 14200 11250 15000 11280
rect 11973 11248 15000 11250
rect 11973 11192 11978 11248
rect 12034 11192 15000 11248
rect 11973 11190 15000 11192
rect 11973 11187 12039 11190
rect 14200 11160 15000 11190
rect 8208 10912 8528 10913
rect 8208 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8528 10912
rect 8208 10847 8528 10848
rect 0 10706 800 10736
rect 1669 10706 1735 10709
rect 0 10704 1735 10706
rect 0 10648 1674 10704
rect 1730 10648 1735 10704
rect 0 10646 1735 10648
rect 0 10616 800 10646
rect 1669 10643 1735 10646
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 12208 10368 12528 10369
rect 12208 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12528 10368
rect 12208 10303 12528 10304
rect 10501 10026 10567 10029
rect 13077 10026 13143 10029
rect 10501 10024 13143 10026
rect 10501 9968 10506 10024
rect 10562 9968 13082 10024
rect 13138 9968 13143 10024
rect 10501 9966 13143 9968
rect 10501 9963 10567 9966
rect 13077 9963 13143 9966
rect 8208 9824 8528 9825
rect 0 9754 800 9784
rect 8208 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8528 9824
rect 8208 9759 8528 9760
rect 1761 9754 1827 9757
rect 0 9752 1827 9754
rect 0 9696 1766 9752
rect 1822 9696 1827 9752
rect 0 9694 1827 9696
rect 0 9664 800 9694
rect 1761 9691 1827 9694
rect 9673 9754 9739 9757
rect 10317 9754 10383 9757
rect 10869 9754 10935 9757
rect 9673 9752 10935 9754
rect 9673 9696 9678 9752
rect 9734 9696 10322 9752
rect 10378 9696 10874 9752
rect 10930 9696 10935 9752
rect 9673 9694 10935 9696
rect 9673 9691 9739 9694
rect 10317 9691 10383 9694
rect 10869 9691 10935 9694
rect 7465 9618 7531 9621
rect 8477 9618 8543 9621
rect 9121 9618 9187 9621
rect 7465 9616 9187 9618
rect 7465 9560 7470 9616
rect 7526 9560 8482 9616
rect 8538 9560 9126 9616
rect 9182 9560 9187 9616
rect 7465 9558 9187 9560
rect 7465 9555 7531 9558
rect 8477 9555 8543 9558
rect 9121 9555 9187 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 12208 9280 12528 9281
rect 12208 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12528 9280
rect 12208 9215 12528 9216
rect 0 8802 800 8832
rect 1669 8802 1735 8805
rect 0 8800 1735 8802
rect 0 8744 1674 8800
rect 1730 8744 1735 8800
rect 0 8742 1735 8744
rect 0 8712 800 8742
rect 1669 8739 1735 8742
rect 13169 8802 13235 8805
rect 14200 8802 15000 8832
rect 13169 8800 15000 8802
rect 13169 8744 13174 8800
rect 13230 8744 15000 8800
rect 13169 8742 15000 8744
rect 13169 8739 13235 8742
rect 8208 8736 8528 8737
rect 8208 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8528 8736
rect 14200 8712 15000 8742
rect 8208 8671 8528 8672
rect 8201 8530 8267 8533
rect 9857 8530 9923 8533
rect 10225 8530 10291 8533
rect 8201 8528 10291 8530
rect 8201 8472 8206 8528
rect 8262 8472 9862 8528
rect 9918 8472 10230 8528
rect 10286 8472 10291 8528
rect 8201 8470 10291 8472
rect 8201 8467 8267 8470
rect 9857 8467 9923 8470
rect 10225 8467 10291 8470
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 12208 8192 12528 8193
rect 12208 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12528 8192
rect 12208 8127 12528 8128
rect 0 7986 800 8016
rect 1485 7986 1551 7989
rect 0 7984 1551 7986
rect 0 7928 1490 7984
rect 1546 7928 1551 7984
rect 0 7926 1551 7928
rect 0 7896 800 7926
rect 1485 7923 1551 7926
rect 1761 7850 1827 7853
rect 8845 7850 8911 7853
rect 1761 7848 8911 7850
rect 1761 7792 1766 7848
rect 1822 7792 8850 7848
rect 8906 7792 8911 7848
rect 1761 7790 8911 7792
rect 1761 7787 1827 7790
rect 8845 7787 8911 7790
rect 8208 7648 8528 7649
rect 8208 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8528 7648
rect 8208 7583 8528 7584
rect 4208 7104 4528 7105
rect 0 7034 800 7064
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 12208 7104 12528 7105
rect 12208 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12528 7104
rect 12208 7039 12528 7040
rect 3969 7034 4035 7037
rect 0 7032 4035 7034
rect 0 6976 3974 7032
rect 4030 6976 4035 7032
rect 0 6974 4035 6976
rect 0 6944 800 6974
rect 3969 6971 4035 6974
rect 8208 6560 8528 6561
rect 8208 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8528 6560
rect 8208 6495 8528 6496
rect 1669 6218 1735 6221
rect 3969 6218 4035 6221
rect 1669 6216 4035 6218
rect 1669 6160 1674 6216
rect 1730 6160 3974 6216
rect 4030 6160 4035 6216
rect 1669 6158 4035 6160
rect 1669 6155 1735 6158
rect 3969 6155 4035 6158
rect 9673 6218 9739 6221
rect 10041 6218 10107 6221
rect 9673 6216 10107 6218
rect 9673 6160 9678 6216
rect 9734 6160 10046 6216
rect 10102 6160 10107 6216
rect 9673 6158 10107 6160
rect 9673 6155 9739 6158
rect 10041 6155 10107 6158
rect 13261 6218 13327 6221
rect 14200 6218 15000 6248
rect 13261 6216 15000 6218
rect 13261 6160 13266 6216
rect 13322 6160 15000 6216
rect 13261 6158 15000 6160
rect 13261 6155 13327 6158
rect 14200 6128 15000 6158
rect 0 6082 800 6112
rect 1669 6082 1735 6085
rect 0 6080 1735 6082
rect 0 6024 1674 6080
rect 1730 6024 1735 6080
rect 0 6022 1735 6024
rect 0 5992 800 6022
rect 1669 6019 1735 6022
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 12208 6016 12528 6017
rect 12208 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12528 6016
rect 12208 5951 12528 5952
rect 8208 5472 8528 5473
rect 8208 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8528 5472
rect 8208 5407 8528 5408
rect 3049 5266 3115 5269
rect 4429 5266 4495 5269
rect 3049 5264 4495 5266
rect 3049 5208 3054 5264
rect 3110 5208 4434 5264
rect 4490 5208 4495 5264
rect 3049 5206 4495 5208
rect 3049 5203 3115 5206
rect 4429 5203 4495 5206
rect 0 5130 800 5160
rect 1577 5130 1643 5133
rect 0 5128 1643 5130
rect 0 5072 1582 5128
rect 1638 5072 1643 5128
rect 0 5070 1643 5072
rect 0 5040 800 5070
rect 1577 5067 1643 5070
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 12208 4928 12528 4929
rect 12208 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12528 4928
rect 12208 4863 12528 4864
rect 8208 4384 8528 4385
rect 8208 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8528 4384
rect 8208 4319 8528 4320
rect 0 4178 800 4208
rect 1761 4178 1827 4181
rect 0 4176 1827 4178
rect 0 4120 1766 4176
rect 1822 4120 1827 4176
rect 0 4118 1827 4120
rect 0 4088 800 4118
rect 1761 4115 1827 4118
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 12208 3840 12528 3841
rect 12208 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12528 3840
rect 12208 3775 12528 3776
rect 12893 3770 12959 3773
rect 14200 3770 15000 3800
rect 12893 3768 15000 3770
rect 12893 3712 12898 3768
rect 12954 3712 15000 3768
rect 12893 3710 15000 3712
rect 12893 3707 12959 3710
rect 14200 3680 15000 3710
rect 8208 3296 8528 3297
rect 0 3226 800 3256
rect 8208 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8528 3296
rect 8208 3231 8528 3232
rect 1577 3226 1643 3229
rect 2681 3226 2747 3229
rect 0 3224 2747 3226
rect 0 3168 1582 3224
rect 1638 3168 2686 3224
rect 2742 3168 2747 3224
rect 0 3166 2747 3168
rect 0 3136 800 3166
rect 1577 3163 1643 3166
rect 2681 3163 2747 3166
rect 2497 3090 2563 3093
rect 6085 3090 6151 3093
rect 2497 3088 6151 3090
rect 2497 3032 2502 3088
rect 2558 3032 6090 3088
rect 6146 3032 6151 3088
rect 2497 3030 6151 3032
rect 2497 3027 2563 3030
rect 6085 3027 6151 3030
rect 4061 2954 4127 2957
rect 7005 2954 7071 2957
rect 4061 2952 7071 2954
rect 4061 2896 4066 2952
rect 4122 2896 7010 2952
rect 7066 2896 7071 2952
rect 4061 2894 7071 2896
rect 4061 2891 4127 2894
rect 7005 2891 7071 2894
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 12208 2752 12528 2753
rect 12208 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12528 2752
rect 12208 2687 12528 2688
rect 4889 2546 4955 2549
rect 5809 2546 5875 2549
rect 4889 2544 5875 2546
rect 4889 2488 4894 2544
rect 4950 2488 5814 2544
rect 5870 2488 5875 2544
rect 4889 2486 5875 2488
rect 4889 2483 4955 2486
rect 5809 2483 5875 2486
rect 8109 2410 8175 2413
rect 9397 2410 9463 2413
rect 8109 2408 9463 2410
rect 8109 2352 8114 2408
rect 8170 2352 9402 2408
rect 9458 2352 9463 2408
rect 8109 2350 9463 2352
rect 8109 2347 8175 2350
rect 9397 2347 9463 2350
rect 0 2274 800 2304
rect 1761 2274 1827 2277
rect 0 2272 1827 2274
rect 0 2216 1766 2272
rect 1822 2216 1827 2272
rect 0 2214 1827 2216
rect 0 2184 800 2214
rect 1761 2211 1827 2214
rect 8208 2208 8528 2209
rect 8208 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8528 2208
rect 8208 2143 8528 2144
rect 4208 1664 4528 1665
rect 4208 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4528 1664
rect 4208 1599 4528 1600
rect 12208 1664 12528 1665
rect 12208 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12528 1664
rect 12208 1599 12528 1600
rect 0 1322 800 1352
rect 3233 1322 3299 1325
rect 0 1320 3299 1322
rect 0 1264 3238 1320
rect 3294 1264 3299 1320
rect 0 1262 3299 1264
rect 0 1232 800 1262
rect 3233 1259 3299 1262
rect 10777 1322 10843 1325
rect 14200 1322 15000 1352
rect 10777 1320 15000 1322
rect 10777 1264 10782 1320
rect 10838 1264 15000 1320
rect 10777 1262 15000 1264
rect 10777 1259 10843 1262
rect 14200 1232 15000 1262
rect 8208 1120 8528 1121
rect 8208 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8528 1120
rect 8208 1055 8528 1056
rect 0 506 800 536
rect 1577 506 1643 509
rect 0 504 1643 506
rect 0 448 1582 504
rect 1638 448 1643 504
rect 0 446 1643 448
rect 0 416 800 446
rect 1577 443 1643 446
<< via3 >>
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 12216 13628 12280 13632
rect 12216 13572 12220 13628
rect 12220 13572 12276 13628
rect 12276 13572 12280 13628
rect 12216 13568 12280 13572
rect 12296 13628 12360 13632
rect 12296 13572 12300 13628
rect 12300 13572 12356 13628
rect 12356 13572 12360 13628
rect 12296 13568 12360 13572
rect 12376 13628 12440 13632
rect 12376 13572 12380 13628
rect 12380 13572 12436 13628
rect 12436 13572 12440 13628
rect 12376 13568 12440 13572
rect 12456 13628 12520 13632
rect 12456 13572 12460 13628
rect 12460 13572 12516 13628
rect 12516 13572 12520 13628
rect 12456 13568 12520 13572
rect 8216 13084 8280 13088
rect 8216 13028 8220 13084
rect 8220 13028 8276 13084
rect 8276 13028 8280 13084
rect 8216 13024 8280 13028
rect 8296 13084 8360 13088
rect 8296 13028 8300 13084
rect 8300 13028 8356 13084
rect 8356 13028 8360 13084
rect 8296 13024 8360 13028
rect 8376 13084 8440 13088
rect 8376 13028 8380 13084
rect 8380 13028 8436 13084
rect 8436 13028 8440 13084
rect 8376 13024 8440 13028
rect 8456 13084 8520 13088
rect 8456 13028 8460 13084
rect 8460 13028 8516 13084
rect 8516 13028 8520 13084
rect 8456 13024 8520 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 12216 12540 12280 12544
rect 12216 12484 12220 12540
rect 12220 12484 12276 12540
rect 12276 12484 12280 12540
rect 12216 12480 12280 12484
rect 12296 12540 12360 12544
rect 12296 12484 12300 12540
rect 12300 12484 12356 12540
rect 12356 12484 12360 12540
rect 12296 12480 12360 12484
rect 12376 12540 12440 12544
rect 12376 12484 12380 12540
rect 12380 12484 12436 12540
rect 12436 12484 12440 12540
rect 12376 12480 12440 12484
rect 12456 12540 12520 12544
rect 12456 12484 12460 12540
rect 12460 12484 12516 12540
rect 12516 12484 12520 12540
rect 12456 12480 12520 12484
rect 8216 11996 8280 12000
rect 8216 11940 8220 11996
rect 8220 11940 8276 11996
rect 8276 11940 8280 11996
rect 8216 11936 8280 11940
rect 8296 11996 8360 12000
rect 8296 11940 8300 11996
rect 8300 11940 8356 11996
rect 8356 11940 8360 11996
rect 8296 11936 8360 11940
rect 8376 11996 8440 12000
rect 8376 11940 8380 11996
rect 8380 11940 8436 11996
rect 8436 11940 8440 11996
rect 8376 11936 8440 11940
rect 8456 11996 8520 12000
rect 8456 11940 8460 11996
rect 8460 11940 8516 11996
rect 8516 11940 8520 11996
rect 8456 11936 8520 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 12216 11452 12280 11456
rect 12216 11396 12220 11452
rect 12220 11396 12276 11452
rect 12276 11396 12280 11452
rect 12216 11392 12280 11396
rect 12296 11452 12360 11456
rect 12296 11396 12300 11452
rect 12300 11396 12356 11452
rect 12356 11396 12360 11452
rect 12296 11392 12360 11396
rect 12376 11452 12440 11456
rect 12376 11396 12380 11452
rect 12380 11396 12436 11452
rect 12436 11396 12440 11452
rect 12376 11392 12440 11396
rect 12456 11452 12520 11456
rect 12456 11396 12460 11452
rect 12460 11396 12516 11452
rect 12516 11396 12520 11452
rect 12456 11392 12520 11396
rect 8216 10908 8280 10912
rect 8216 10852 8220 10908
rect 8220 10852 8276 10908
rect 8276 10852 8280 10908
rect 8216 10848 8280 10852
rect 8296 10908 8360 10912
rect 8296 10852 8300 10908
rect 8300 10852 8356 10908
rect 8356 10852 8360 10908
rect 8296 10848 8360 10852
rect 8376 10908 8440 10912
rect 8376 10852 8380 10908
rect 8380 10852 8436 10908
rect 8436 10852 8440 10908
rect 8376 10848 8440 10852
rect 8456 10908 8520 10912
rect 8456 10852 8460 10908
rect 8460 10852 8516 10908
rect 8516 10852 8520 10908
rect 8456 10848 8520 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 12216 10364 12280 10368
rect 12216 10308 12220 10364
rect 12220 10308 12276 10364
rect 12276 10308 12280 10364
rect 12216 10304 12280 10308
rect 12296 10364 12360 10368
rect 12296 10308 12300 10364
rect 12300 10308 12356 10364
rect 12356 10308 12360 10364
rect 12296 10304 12360 10308
rect 12376 10364 12440 10368
rect 12376 10308 12380 10364
rect 12380 10308 12436 10364
rect 12436 10308 12440 10364
rect 12376 10304 12440 10308
rect 12456 10364 12520 10368
rect 12456 10308 12460 10364
rect 12460 10308 12516 10364
rect 12516 10308 12520 10364
rect 12456 10304 12520 10308
rect 8216 9820 8280 9824
rect 8216 9764 8220 9820
rect 8220 9764 8276 9820
rect 8276 9764 8280 9820
rect 8216 9760 8280 9764
rect 8296 9820 8360 9824
rect 8296 9764 8300 9820
rect 8300 9764 8356 9820
rect 8356 9764 8360 9820
rect 8296 9760 8360 9764
rect 8376 9820 8440 9824
rect 8376 9764 8380 9820
rect 8380 9764 8436 9820
rect 8436 9764 8440 9820
rect 8376 9760 8440 9764
rect 8456 9820 8520 9824
rect 8456 9764 8460 9820
rect 8460 9764 8516 9820
rect 8516 9764 8520 9820
rect 8456 9760 8520 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 12216 9276 12280 9280
rect 12216 9220 12220 9276
rect 12220 9220 12276 9276
rect 12276 9220 12280 9276
rect 12216 9216 12280 9220
rect 12296 9276 12360 9280
rect 12296 9220 12300 9276
rect 12300 9220 12356 9276
rect 12356 9220 12360 9276
rect 12296 9216 12360 9220
rect 12376 9276 12440 9280
rect 12376 9220 12380 9276
rect 12380 9220 12436 9276
rect 12436 9220 12440 9276
rect 12376 9216 12440 9220
rect 12456 9276 12520 9280
rect 12456 9220 12460 9276
rect 12460 9220 12516 9276
rect 12516 9220 12520 9276
rect 12456 9216 12520 9220
rect 8216 8732 8280 8736
rect 8216 8676 8220 8732
rect 8220 8676 8276 8732
rect 8276 8676 8280 8732
rect 8216 8672 8280 8676
rect 8296 8732 8360 8736
rect 8296 8676 8300 8732
rect 8300 8676 8356 8732
rect 8356 8676 8360 8732
rect 8296 8672 8360 8676
rect 8376 8732 8440 8736
rect 8376 8676 8380 8732
rect 8380 8676 8436 8732
rect 8436 8676 8440 8732
rect 8376 8672 8440 8676
rect 8456 8732 8520 8736
rect 8456 8676 8460 8732
rect 8460 8676 8516 8732
rect 8516 8676 8520 8732
rect 8456 8672 8520 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 12216 8188 12280 8192
rect 12216 8132 12220 8188
rect 12220 8132 12276 8188
rect 12276 8132 12280 8188
rect 12216 8128 12280 8132
rect 12296 8188 12360 8192
rect 12296 8132 12300 8188
rect 12300 8132 12356 8188
rect 12356 8132 12360 8188
rect 12296 8128 12360 8132
rect 12376 8188 12440 8192
rect 12376 8132 12380 8188
rect 12380 8132 12436 8188
rect 12436 8132 12440 8188
rect 12376 8128 12440 8132
rect 12456 8188 12520 8192
rect 12456 8132 12460 8188
rect 12460 8132 12516 8188
rect 12516 8132 12520 8188
rect 12456 8128 12520 8132
rect 8216 7644 8280 7648
rect 8216 7588 8220 7644
rect 8220 7588 8276 7644
rect 8276 7588 8280 7644
rect 8216 7584 8280 7588
rect 8296 7644 8360 7648
rect 8296 7588 8300 7644
rect 8300 7588 8356 7644
rect 8356 7588 8360 7644
rect 8296 7584 8360 7588
rect 8376 7644 8440 7648
rect 8376 7588 8380 7644
rect 8380 7588 8436 7644
rect 8436 7588 8440 7644
rect 8376 7584 8440 7588
rect 8456 7644 8520 7648
rect 8456 7588 8460 7644
rect 8460 7588 8516 7644
rect 8516 7588 8520 7644
rect 8456 7584 8520 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 12216 7100 12280 7104
rect 12216 7044 12220 7100
rect 12220 7044 12276 7100
rect 12276 7044 12280 7100
rect 12216 7040 12280 7044
rect 12296 7100 12360 7104
rect 12296 7044 12300 7100
rect 12300 7044 12356 7100
rect 12356 7044 12360 7100
rect 12296 7040 12360 7044
rect 12376 7100 12440 7104
rect 12376 7044 12380 7100
rect 12380 7044 12436 7100
rect 12436 7044 12440 7100
rect 12376 7040 12440 7044
rect 12456 7100 12520 7104
rect 12456 7044 12460 7100
rect 12460 7044 12516 7100
rect 12516 7044 12520 7100
rect 12456 7040 12520 7044
rect 8216 6556 8280 6560
rect 8216 6500 8220 6556
rect 8220 6500 8276 6556
rect 8276 6500 8280 6556
rect 8216 6496 8280 6500
rect 8296 6556 8360 6560
rect 8296 6500 8300 6556
rect 8300 6500 8356 6556
rect 8356 6500 8360 6556
rect 8296 6496 8360 6500
rect 8376 6556 8440 6560
rect 8376 6500 8380 6556
rect 8380 6500 8436 6556
rect 8436 6500 8440 6556
rect 8376 6496 8440 6500
rect 8456 6556 8520 6560
rect 8456 6500 8460 6556
rect 8460 6500 8516 6556
rect 8516 6500 8520 6556
rect 8456 6496 8520 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 12216 6012 12280 6016
rect 12216 5956 12220 6012
rect 12220 5956 12276 6012
rect 12276 5956 12280 6012
rect 12216 5952 12280 5956
rect 12296 6012 12360 6016
rect 12296 5956 12300 6012
rect 12300 5956 12356 6012
rect 12356 5956 12360 6012
rect 12296 5952 12360 5956
rect 12376 6012 12440 6016
rect 12376 5956 12380 6012
rect 12380 5956 12436 6012
rect 12436 5956 12440 6012
rect 12376 5952 12440 5956
rect 12456 6012 12520 6016
rect 12456 5956 12460 6012
rect 12460 5956 12516 6012
rect 12516 5956 12520 6012
rect 12456 5952 12520 5956
rect 8216 5468 8280 5472
rect 8216 5412 8220 5468
rect 8220 5412 8276 5468
rect 8276 5412 8280 5468
rect 8216 5408 8280 5412
rect 8296 5468 8360 5472
rect 8296 5412 8300 5468
rect 8300 5412 8356 5468
rect 8356 5412 8360 5468
rect 8296 5408 8360 5412
rect 8376 5468 8440 5472
rect 8376 5412 8380 5468
rect 8380 5412 8436 5468
rect 8436 5412 8440 5468
rect 8376 5408 8440 5412
rect 8456 5468 8520 5472
rect 8456 5412 8460 5468
rect 8460 5412 8516 5468
rect 8516 5412 8520 5468
rect 8456 5408 8520 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 12216 4924 12280 4928
rect 12216 4868 12220 4924
rect 12220 4868 12276 4924
rect 12276 4868 12280 4924
rect 12216 4864 12280 4868
rect 12296 4924 12360 4928
rect 12296 4868 12300 4924
rect 12300 4868 12356 4924
rect 12356 4868 12360 4924
rect 12296 4864 12360 4868
rect 12376 4924 12440 4928
rect 12376 4868 12380 4924
rect 12380 4868 12436 4924
rect 12436 4868 12440 4924
rect 12376 4864 12440 4868
rect 12456 4924 12520 4928
rect 12456 4868 12460 4924
rect 12460 4868 12516 4924
rect 12516 4868 12520 4924
rect 12456 4864 12520 4868
rect 8216 4380 8280 4384
rect 8216 4324 8220 4380
rect 8220 4324 8276 4380
rect 8276 4324 8280 4380
rect 8216 4320 8280 4324
rect 8296 4380 8360 4384
rect 8296 4324 8300 4380
rect 8300 4324 8356 4380
rect 8356 4324 8360 4380
rect 8296 4320 8360 4324
rect 8376 4380 8440 4384
rect 8376 4324 8380 4380
rect 8380 4324 8436 4380
rect 8436 4324 8440 4380
rect 8376 4320 8440 4324
rect 8456 4380 8520 4384
rect 8456 4324 8460 4380
rect 8460 4324 8516 4380
rect 8516 4324 8520 4380
rect 8456 4320 8520 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 12216 3836 12280 3840
rect 12216 3780 12220 3836
rect 12220 3780 12276 3836
rect 12276 3780 12280 3836
rect 12216 3776 12280 3780
rect 12296 3836 12360 3840
rect 12296 3780 12300 3836
rect 12300 3780 12356 3836
rect 12356 3780 12360 3836
rect 12296 3776 12360 3780
rect 12376 3836 12440 3840
rect 12376 3780 12380 3836
rect 12380 3780 12436 3836
rect 12436 3780 12440 3836
rect 12376 3776 12440 3780
rect 12456 3836 12520 3840
rect 12456 3780 12460 3836
rect 12460 3780 12516 3836
rect 12516 3780 12520 3836
rect 12456 3776 12520 3780
rect 8216 3292 8280 3296
rect 8216 3236 8220 3292
rect 8220 3236 8276 3292
rect 8276 3236 8280 3292
rect 8216 3232 8280 3236
rect 8296 3292 8360 3296
rect 8296 3236 8300 3292
rect 8300 3236 8356 3292
rect 8356 3236 8360 3292
rect 8296 3232 8360 3236
rect 8376 3292 8440 3296
rect 8376 3236 8380 3292
rect 8380 3236 8436 3292
rect 8436 3236 8440 3292
rect 8376 3232 8440 3236
rect 8456 3292 8520 3296
rect 8456 3236 8460 3292
rect 8460 3236 8516 3292
rect 8516 3236 8520 3292
rect 8456 3232 8520 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 12216 2748 12280 2752
rect 12216 2692 12220 2748
rect 12220 2692 12276 2748
rect 12276 2692 12280 2748
rect 12216 2688 12280 2692
rect 12296 2748 12360 2752
rect 12296 2692 12300 2748
rect 12300 2692 12356 2748
rect 12356 2692 12360 2748
rect 12296 2688 12360 2692
rect 12376 2748 12440 2752
rect 12376 2692 12380 2748
rect 12380 2692 12436 2748
rect 12436 2692 12440 2748
rect 12376 2688 12440 2692
rect 12456 2748 12520 2752
rect 12456 2692 12460 2748
rect 12460 2692 12516 2748
rect 12516 2692 12520 2748
rect 12456 2688 12520 2692
rect 8216 2204 8280 2208
rect 8216 2148 8220 2204
rect 8220 2148 8276 2204
rect 8276 2148 8280 2204
rect 8216 2144 8280 2148
rect 8296 2204 8360 2208
rect 8296 2148 8300 2204
rect 8300 2148 8356 2204
rect 8356 2148 8360 2204
rect 8296 2144 8360 2148
rect 8376 2204 8440 2208
rect 8376 2148 8380 2204
rect 8380 2148 8436 2204
rect 8436 2148 8440 2204
rect 8376 2144 8440 2148
rect 8456 2204 8520 2208
rect 8456 2148 8460 2204
rect 8460 2148 8516 2204
rect 8516 2148 8520 2204
rect 8456 2144 8520 2148
rect 4216 1660 4280 1664
rect 4216 1604 4220 1660
rect 4220 1604 4276 1660
rect 4276 1604 4280 1660
rect 4216 1600 4280 1604
rect 4296 1660 4360 1664
rect 4296 1604 4300 1660
rect 4300 1604 4356 1660
rect 4356 1604 4360 1660
rect 4296 1600 4360 1604
rect 4376 1660 4440 1664
rect 4376 1604 4380 1660
rect 4380 1604 4436 1660
rect 4436 1604 4440 1660
rect 4376 1600 4440 1604
rect 4456 1660 4520 1664
rect 4456 1604 4460 1660
rect 4460 1604 4516 1660
rect 4516 1604 4520 1660
rect 4456 1600 4520 1604
rect 12216 1660 12280 1664
rect 12216 1604 12220 1660
rect 12220 1604 12276 1660
rect 12276 1604 12280 1660
rect 12216 1600 12280 1604
rect 12296 1660 12360 1664
rect 12296 1604 12300 1660
rect 12300 1604 12356 1660
rect 12356 1604 12360 1660
rect 12296 1600 12360 1604
rect 12376 1660 12440 1664
rect 12376 1604 12380 1660
rect 12380 1604 12436 1660
rect 12436 1604 12440 1660
rect 12376 1600 12440 1604
rect 12456 1660 12520 1664
rect 12456 1604 12460 1660
rect 12460 1604 12516 1660
rect 12516 1604 12520 1660
rect 12456 1600 12520 1604
rect 8216 1116 8280 1120
rect 8216 1060 8220 1116
rect 8220 1060 8276 1116
rect 8276 1060 8280 1116
rect 8216 1056 8280 1060
rect 8296 1116 8360 1120
rect 8296 1060 8300 1116
rect 8300 1060 8356 1116
rect 8356 1060 8360 1116
rect 8296 1056 8360 1060
rect 8376 1116 8440 1120
rect 8376 1060 8380 1116
rect 8380 1060 8436 1116
rect 8436 1060 8440 1116
rect 8376 1056 8440 1060
rect 8456 1116 8520 1120
rect 8456 1060 8460 1116
rect 8460 1060 8516 1116
rect 8516 1060 8520 1116
rect 8456 1056 8520 1060
<< metal4 >>
rect 4208 13632 4528 13648
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12488 4296 12544
rect 4360 12488 4376 12544
rect 4440 12488 4456 12544
rect 4520 12480 4528 12544
rect 4208 12252 4250 12480
rect 4486 12252 4528 12480
rect 4208 11456 4528 12252
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4488 4528 4864
rect 4208 4252 4250 4488
rect 4486 4252 4528 4488
rect 4208 3840 4528 4252
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 1664 4528 2688
rect 4208 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4528 1664
rect 4208 1040 4528 1600
rect 8208 13088 8528 13648
rect 8208 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8528 13088
rect 8208 12000 8528 13024
rect 8208 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8528 12000
rect 8208 10912 8528 11936
rect 8208 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8528 10912
rect 8208 9824 8528 10848
rect 8208 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8528 9824
rect 8208 8736 8528 9760
rect 8208 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8528 8736
rect 8208 8488 8528 8672
rect 8208 8252 8250 8488
rect 8486 8252 8528 8488
rect 8208 7648 8528 8252
rect 8208 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8528 7648
rect 8208 6560 8528 7584
rect 8208 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8528 6560
rect 8208 5472 8528 6496
rect 8208 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8528 5472
rect 8208 4384 8528 5408
rect 8208 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8528 4384
rect 8208 3296 8528 4320
rect 8208 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8528 3296
rect 8208 2208 8528 3232
rect 8208 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8528 2208
rect 8208 1120 8528 2144
rect 8208 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8528 1120
rect 8208 1040 8528 1056
rect 12208 13632 12528 13648
rect 12208 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12528 13632
rect 12208 12544 12528 13568
rect 12208 12480 12216 12544
rect 12280 12488 12296 12544
rect 12360 12488 12376 12544
rect 12440 12488 12456 12544
rect 12520 12480 12528 12544
rect 12208 12252 12250 12480
rect 12486 12252 12528 12480
rect 12208 11456 12528 12252
rect 12208 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12528 11456
rect 12208 10368 12528 11392
rect 12208 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12528 10368
rect 12208 9280 12528 10304
rect 12208 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12528 9280
rect 12208 8192 12528 9216
rect 12208 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12528 8192
rect 12208 7104 12528 8128
rect 12208 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12528 7104
rect 12208 6016 12528 7040
rect 12208 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12528 6016
rect 12208 4928 12528 5952
rect 12208 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12528 4928
rect 12208 4488 12528 4864
rect 12208 4252 12250 4488
rect 12486 4252 12528 4488
rect 12208 3840 12528 4252
rect 12208 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12528 3840
rect 12208 2752 12528 3776
rect 12208 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12528 2752
rect 12208 1664 12528 2688
rect 12208 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12528 1664
rect 12208 1040 12528 1600
<< via4 >>
rect 4250 12480 4280 12488
rect 4280 12480 4296 12488
rect 4296 12480 4360 12488
rect 4360 12480 4376 12488
rect 4376 12480 4440 12488
rect 4440 12480 4456 12488
rect 4456 12480 4486 12488
rect 4250 12252 4486 12480
rect 4250 4252 4486 4488
rect 8250 8252 8486 8488
rect 12250 12480 12280 12488
rect 12280 12480 12296 12488
rect 12296 12480 12360 12488
rect 12360 12480 12376 12488
rect 12376 12480 12440 12488
rect 12440 12480 12456 12488
rect 12456 12480 12486 12488
rect 12250 12252 12486 12480
rect 12250 4252 12486 4488
<< metal5 >>
rect 1104 12488 13892 12530
rect 1104 12252 4250 12488
rect 4486 12252 12250 12488
rect 12486 12252 13892 12488
rect 1104 12210 13892 12252
rect 1104 8488 13892 8530
rect 1104 8252 8250 8488
rect 8486 8252 13892 8488
rect 1104 8210 13892 8252
rect 1104 4488 13892 4530
rect 1104 4252 4250 4488
rect 4486 4252 12250 4488
rect 12486 4252 13892 4488
rect 1104 4210 13892 4252
use sky130_fd_sc_hd__fill_1  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 1380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 2852 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1638025753
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 1380 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 1840 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _328_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 1840 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 2576 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _376_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 1564 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 4508 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 3680 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 4140 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 5612 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _184_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 4508 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _361_
timestamp 1638025753
transform -1 0 6072 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52
timestamp 1638025753
transform 1 0 5888 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62
timestamp 1638025753
transform 1 0 6808 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1638025753
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1638025753
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1638025753
transform 1 0 6072 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 6256 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _320_
timestamp 1638025753
transform -1 0 5888 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 6348 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _360_
timestamp 1638025753
transform 1 0 6348 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_1_78
timestamp 1638025753
transform 1 0 8280 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66
timestamp 1638025753
transform 1 0 7176 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_70 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 7544 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1638025753
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1638025753
transform 1 0 8648 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _321_
timestamp 1638025753
transform 1 0 7268 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _189_
timestamp 1638025753
transform -1 0 9384 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _371_
timestamp 1638025753
transform 1 0 8372 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_0_105
timestamp 1638025753
transform 1 0 10764 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_93
timestamp 1638025753
transform 1 0 9660 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _309_
timestamp 1638025753
transform -1 0 11316 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _310_
timestamp 1638025753
transform 1 0 9384 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _325_
timestamp 1638025753
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _188_
timestamp 1638025753
transform -1 0 11040 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1638025753
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1638025753
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1638025753
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1638025753
transform 1 0 11500 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _356_
timestamp 1638025753
transform 1 0 11500 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _357_
timestamp 1638025753
transform 1 0 11684 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1638025753
transform -1 0 13892 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1638025753
transform -1 0 13892 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_134
timestamp 1638025753
transform 1 0 13432 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_18
timestamp 1638025753
transform 1 0 2760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1638025753
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1638025753
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _209_
timestamp 1638025753
transform -1 0 2760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_2  _200_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 2852 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 1656 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1638025753
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1638025753
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 5520 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_2  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 4600 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _275_
timestamp 1638025753
transform 1 0 5520 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2ai_2  _206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_78
timestamp 1638025753
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1638025753
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _306_
timestamp 1638025753
transform -1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _185_
timestamp 1638025753
transform -1 0 9660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_2  _194_
timestamp 1638025753
transform 1 0 7452 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1638025753
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _372_
timestamp 1638025753
transform 1 0 9936 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_2_120
timestamp 1638025753
transform 1 0 12144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _308_
timestamp 1638025753
transform -1 0 12144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _324_
timestamp 1638025753
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_2  _178_
timestamp 1638025753
transform 1 0 12604 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1638025753
transform -1 0 13892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_134
timestamp 1638025753
transform 1 0 13432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1638025753
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1638025753
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 1932 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1638025753
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_2  _225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 1932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_37
timestamp 1638025753
transform 1 0 4508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_33
timestamp 1638025753
transform 1 0 4140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_24
timestamp 1638025753
transform 1 0 3312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1638025753
transform -1 0 4876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1638025753
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 4876 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1638025753
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_48
timestamp 1638025753
transform 1 0 5520 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1638025753
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _193_
timestamp 1638025753
transform 1 0 6440 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _208_
timestamp 1638025753
transform 1 0 5612 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _195_
timestamp 1638025753
transform -1 0 7636 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_71
timestamp 1638025753
transform 1 0 7636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _375_
timestamp 1638025753
transform -1 0 9752 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_3_94
timestamp 1638025753
transform 1 0 9752 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _187_
timestamp 1638025753
transform 1 0 9844 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and4_2  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 11316 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1638025753
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1638025753
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1638025753
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _358_
timestamp 1638025753
transform 1 0 11684 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1638025753
transform -1 0 13892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1638025753
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1638025753
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_2  _211_
timestamp 1638025753
transform -1 0 2944 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _183_
timestamp 1638025753
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_2  _204_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 2300 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1638025753
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _377_
timestamp 1638025753
transform -1 0 5704 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_4_58
timestamp 1638025753
transform 1 0 6440 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _374_
timestamp 1638025753
transform 1 0 6624 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__and4_2  _272_
timestamp 1638025753
transform 1 0 5704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1638025753
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1638025753
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _233_
timestamp 1638025753
transform 1 0 9660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_2  _373_
timestamp 1638025753
transform 1 0 10212 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_4_120
timestamp 1638025753
transform 1 0 12144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_129
timestamp 1638025753
transform 1 0 12972 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _316_
timestamp 1638025753
transform 1 0 12420 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _323_
timestamp 1638025753
transform 1 0 12696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_135
timestamp 1638025753
transform 1 0 13524 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1638025753
transform -1 0 13892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_19
timestamp 1638025753
transform 1 0 2852 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1638025753
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1638025753
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _205_
timestamp 1638025753
transform 1 0 2576 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _190_
timestamp 1638025753
transform 1 0 2944 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _217_
timestamp 1638025753
transform 1 0 1748 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_5_32
timestamp 1638025753
transform 1 0 4048 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _359_
timestamp 1638025753
transform 1 0 4324 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_2  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 3404 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1638025753
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1638025753
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _186_
timestamp 1638025753
transform 1 0 6440 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_69
timestamp 1638025753
transform 1 0 7452 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1638025753
transform -1 0 7452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _307_
timestamp 1638025753
transform 1 0 7544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _364_
timestamp 1638025753
transform 1 0 7820 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_5_103
timestamp 1638025753
transform 1 0 10580 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _237_
timestamp 1638025753
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _234_
timestamp 1638025753
transform -1 0 10580 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1638025753
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _365_
timestamp 1638025753
transform 1 0 11500 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1638025753
transform -1 0 13892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_134
timestamp 1638025753
transform 1 0 13432 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_2  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 1840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _202_
timestamp 1638025753
transform 1 0 1380 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_2  _201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 2392 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1638025753
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1638025753
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1638025753
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _212_
timestamp 1638025753
transform -1 0 3312 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_2  _198_
timestamp 1638025753
transform 1 0 2760 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1638025753
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_17
timestamp 1638025753
transform 1 0 2668 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1638025753
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_39
timestamp 1638025753
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_38
timestamp 1638025753
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1638025753
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _270_
timestamp 1638025753
transform -1 0 4692 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_2  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 4876 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _180_
timestamp 1638025753
transform -1 0 4048 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_2  _213_
timestamp 1638025753
transform -1 0 4600 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _271_
timestamp 1638025753
transform 1 0 4968 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_62
timestamp 1638025753
transform 1 0 6808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_53
timestamp 1638025753
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1638025753
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _269_
timestamp 1638025753
transform 1 0 5796 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1638025753
transform -1 0 6532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _319_
timestamp 1638025753
transform 1 0 6532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _322_
timestamp 1638025753
transform -1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _362_
timestamp 1638025753
transform -1 0 8280 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1638025753
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_71
timestamp 1638025753
transform 1 0 7636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1638025753
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_81
timestamp 1638025753
transform 1 0 8556 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1638025753
transform 1 0 8280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _317_
timestamp 1638025753
transform -1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _219_
timestamp 1638025753
transform 1 0 7176 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _250_
timestamp 1638025753
transform 1 0 8740 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _224_
timestamp 1638025753
transform -1 0 10580 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_2  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 9568 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1638025753
transform -1 0 9568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_90
timestamp 1638025753
transform 1 0 9384 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_96
timestamp 1638025753
transform 1 0 9936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_88
timestamp 1638025753
transform 1 0 9200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o22ai_2  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 11500 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_2  _238_
timestamp 1638025753
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_100
timestamp 1638025753
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_103
timestamp 1638025753
transform 1 0 10580 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_122
timestamp 1638025753
transform 1 0 12328 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1638025753
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_127
timestamp 1638025753
transform 1 0 12788 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_116
timestamp 1638025753
transform 1 0 11776 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1638025753
transform -1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _311_
timestamp 1638025753
transform 1 0 12512 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_2  _264_
timestamp 1638025753
transform -1 0 12328 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_135
timestamp 1638025753
transform 1 0 13524 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1638025753
transform -1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1638025753
transform -1 0 13892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_134
timestamp 1638025753
transform 1 0 13432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1638025753
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1638025753
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_2  _216_
timestamp 1638025753
transform -1 0 2024 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o221ai_2  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 2024 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1638025753
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1638025753
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1638025753
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _214_
timestamp 1638025753
transform -1 0 3588 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _363_
timestamp 1638025753
transform 1 0 3864 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_8_51
timestamp 1638025753
transform 1 0 5796 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_63
timestamp 1638025753
transform 1 0 6900 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_69
timestamp 1638025753
transform 1 0 7452 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1638025753
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1638025753
transform -1 0 8096 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1638025753
transform 1 0 7544 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 8924 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_2  _247_
timestamp 1638025753
transform -1 0 8832 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _366_
timestamp 1638025753
transform 1 0 9752 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _370_
timestamp 1638025753
transform 1 0 11684 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1638025753
transform -1 0 13892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1638025753
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1638025753
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _378_
timestamp 1638025753
transform 1 0 1656 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1638025753
transform 1 0 3588 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 3956 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1638025753
transform -1 0 3956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_52
timestamp 1638025753
transform 1 0 5888 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1638025753
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_47
timestamp 1638025753
transform 1 0 5428 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _312_
timestamp 1638025753
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _313_
timestamp 1638025753
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _318_
timestamp 1638025753
transform -1 0 5428 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _369_
timestamp 1638025753
transform 1 0 6348 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_9_78
timestamp 1638025753
transform 1 0 8280 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_87
timestamp 1638025753
transform 1 0 9108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _256_
timestamp 1638025753
transform -1 0 9108 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1638025753
transform 1 0 8372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _262_
timestamp 1638025753
transform -1 0 9844 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _315_
timestamp 1638025753
transform -1 0 11408 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _258_
timestamp 1638025753
transform 1 0 10672 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _263_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 9844 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1638025753
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1638025753
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _367_
timestamp 1638025753
transform 1 0 11684 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1638025753
transform -1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_15
timestamp 1638025753
transform 1 0 2484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1638025753
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_19
timestamp 1638025753
transform 1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1638025753
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _327_
timestamp 1638025753
transform 1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1638025753
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1638025753
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_34
timestamp 1638025753
transform 1 0 4232 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _181_
timestamp 1638025753
transform 1 0 3772 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1638025753
transform -1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _368_
timestamp 1638025753
transform 1 0 4784 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1638025753
transform -1 0 6992 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1638025753
transform -1 0 7268 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1638025753
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_2  _254_
timestamp 1638025753
transform -1 0 8096 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_2  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_2  _243_
timestamp 1638025753
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_104
timestamp 1638025753
transform 1 0 10672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_94
timestamp 1638025753
transform 1 0 9752 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_2  _240_
timestamp 1638025753
transform -1 0 10672 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_2  _260_
timestamp 1638025753
transform 1 0 10764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_113
timestamp 1638025753
transform 1 0 11500 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _314_
timestamp 1638025753
transform 1 0 12512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _333_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 12788 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_2  _261_
timestamp 1638025753
transform -1 0 12512 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1638025753
transform -1 0 13892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1638025753
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp11
timestamp 1638025753
transform -1 0 2576 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 2944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 3220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_23
timestamp 1638025753
transform 1 0 3220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_38
timestamp 1638025753
transform 1 0 4600 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_32
timestamp 1638025753
transform 1 0 4048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00
timestamp 1638025753
transform 1 0 4232 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _182_
timestamp 1638025753
transform 1 0 3588 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 1638025753
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1638025753
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_50
timestamp 1638025753
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 6716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _255_
timestamp 1638025753
transform 1 0 6716 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_11_77
timestamp 1638025753
transform 1 0 8188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _251_
timestamp 1638025753
transform 1 0 9108 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _242_
timestamp 1638025753
transform 1 0 8372 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _257_
timestamp 1638025753
transform 1 0 7360 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_101
timestamp 1638025753
transform 1 0 10396 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _259_
timestamp 1638025753
transform 1 0 10488 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_2  _241_
timestamp 1638025753
transform 1 0 9568 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_130
timestamp 1638025753
transform 1 0 13064 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1638025753
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1638025753
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_116
timestamp 1638025753
transform 1 0 11776 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1638025753
transform 1 0 11960 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1638025753
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _326_
timestamp 1638025753
transform -1 0 13432 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _331_
timestamp 1638025753
transform 1 0 12236 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1638025753
transform -1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_134
timestamp 1638025753
transform 1 0 13432 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_19
timestamp 1638025753
transform 1 0 2852 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1638025753
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 2208 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen1
timestamp 1638025753
transform -1 0 3588 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1638025753
transform -1 0 2208 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1638025753
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1638025753
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_39
timestamp 1638025753
transform 1 0 4692 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen0
timestamp 1638025753
transform 1 0 4876 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.reseten0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 3772 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0
timestamp 1638025753
transform -1 0 4692 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_12_48
timestamp 1638025753
transform 1 0 5520 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen1
timestamp 1638025753
transform -1 0 7360 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 6716 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_12_80
timestamp 1638025753
transform 1 0 8464 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1638025753
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_68
timestamp 1638025753
transform 1 0 7360 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1638025753
transform -1 0 8832 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1638025753
transform 1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1638025753
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _252_
timestamp 1638025753
transform 1 0 7544 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_12_105
timestamp 1638025753
transform 1 0 10764 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_99
timestamp 1638025753
transform 1 0 10212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen1
timestamp 1638025753
transform -1 0 11776 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _170_
timestamp 1638025753
transform 1 0 10488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _239_
timestamp 1638025753
transform -1 0 10212 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1638025753
transform -1 0 11132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen1
timestamp 1638025753
transform 1 0 12788 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb1
timestamp 1638025753
transform -1 0 12788 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1638025753
transform -1 0 13892 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_134
timestamp 1638025753
transform 1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1638025753
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_13
timestamp 1638025753
transform 1 0 2300 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1638025753
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1638025753
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1638025753
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp 1638025753
transform 1 0 2392 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 3036 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1638025753
transform -1 0 2300 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[0\].id.delayenb0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 1564 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_14_43
timestamp 1638025753
transform 1 0 5060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1638025753
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 4784 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_34
timestamp 1638025753
transform 1 0 4232 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1638025753
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen1
timestamp 1638025753
transform -1 0 4416 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0
timestamp 1638025753
transform -1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[0\].id.delayenb1
timestamp 1638025753
transform -1 0 4232 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_8  ringosc.iss.delayenb0
timestamp 1638025753
transform 1 0 4416 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_14_63
timestamp 1638025753
transform 1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1638025753
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_60
timestamp 1638025753
transform 1 0 6624 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1638025753
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1638025753
transform 1 0 6808 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_2  _289_
timestamp 1638025753
transform 1 0 6164 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1638025753
transform -1 0 6624 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _290_
timestamp 1638025753
transform 1 0 7268 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _291_
timestamp 1638025753
transform 1 0 7636 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _229_
timestamp 1638025753
transform 1 0 8280 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _280_
timestamp 1638025753
transform -1 0 8372 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1638025753
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _223_
timestamp 1638025753
transform 1 0 9108 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1638025753
transform 1 0 8740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1638025753
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_86
timestamp 1638025753
transform 1 0 9016 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1638025753
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1638025753
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen0
timestamp 1638025753
transform -1 0 11408 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1638025753
transform -1 0 10764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1638025753
transform 1 0 10120 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_2  _304_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 9200 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _221_
timestamp 1638025753
transform -1 0 10120 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _227_
timestamp 1638025753
transform 1 0 10948 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _232_
timestamp 1638025753
transform -1 0 10488 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 10948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1638025753
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_112
timestamp 1638025753
transform 1 0 11408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1638025753
transform -1 0 13432 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp 1638025753
transform 1 0 11960 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1638025753
transform 1 0 11592 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[10\].id.delayenb1
timestamp 1638025753
transform 1 0 12604 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp 1638025753
transform 1 0 11500 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1638025753
transform -1 0 13892 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1638025753
transform -1 0 13892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_134
timestamp 1638025753
transform 1 0 13432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1638025753
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1638025753
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[1\].id.delayenb0
timestamp 1638025753
transform 1 0 1656 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_15_39
timestamp 1638025753
transform 1 0 4692 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_24
timestamp 1638025753
transform 1 0 3312 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1638025753
transform 1 0 4416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _330_
timestamp 1638025753
transform -1 0 5612 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[1\].id.delayenb1
timestamp 1638025753
transform -1 0 4416 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1638025753
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1638025753
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1638025753
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_2  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 6348 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_15_67
timestamp 1638025753
transform 1 0 7268 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_76
timestamp 1638025753
transform 1 0 8096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__o31a_2  _303_
timestamp 1638025753
transform 1 0 8924 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _278_
timestamp 1638025753
transform -1 0 8096 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _297_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 8280 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1638025753
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_93
timestamp 1638025753
transform 1 0 9660 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1638025753
transform 1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _231_
timestamp 1638025753
transform 1 0 10396 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1638025753
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[10\].id.delayenb0
timestamp 1638025753
transform 1 0 11500 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1638025753
transform -1 0 13432 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1638025753
transform -1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_134
timestamp 1638025753
transform 1 0 13432 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_15
timestamp 1638025753
transform 1 0 2484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1638025753
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1638025753
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1638025753
transform 1 0 2852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1638025753
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1638025753
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1638025753
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_32
timestamp 1638025753
transform 1 0 4048 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _354_
timestamp 1638025753
transform 1 0 4784 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1638025753
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_59
timestamp 1638025753
transform 1 0 6532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_2  _285_
timestamp 1638025753
transform 1 0 6808 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__o41a_2  _286_
timestamp 1638025753
transform 1 0 5612 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  FILLER_16_72
timestamp 1638025753
transform 1 0 7728 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1638025753
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1638025753
transform 1 0 8004 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_2  _298_
timestamp 1638025753
transform 1 0 8924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_98
timestamp 1638025753
transform 1 0 10120 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_94
timestamp 1638025753
transform 1 0 9752 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_2  _300_
timestamp 1638025753
transform 1 0 10212 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or3_2  _294_
timestamp 1638025753
transform 1 0 11132 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_121
timestamp 1638025753
transform 1 0 12236 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_115
timestamp 1638025753
transform 1 0 11684 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1638025753
transform 1 0 12328 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _335_
timestamp 1638025753
transform 1 0 12696 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_135
timestamp 1638025753
transform 1 0 13524 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1638025753
transform -1 0 13892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_12
timestamp 1638025753
transform 1 0 2208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1638025753
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _348_
timestamp 1638025753
transform -1 0 2208 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[2\].id.delayenb1
timestamp 1638025753
transform 1 0 2576 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_17_30
timestamp 1638025753
transform 1 0 3864 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1638025753
transform 1 0 3588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb1
timestamp 1638025753
transform -1 0 5520 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1638025753
transform -1 0 4508 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1638025753
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o31a_2  _281_
timestamp 1638025753
transform 1 0 6808 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _282_
timestamp 1638025753
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _279_
timestamp 1638025753
transform -1 0 6808 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_17_84
timestamp 1638025753
transform 1 0 8832 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _332_
timestamp 1638025753
transform -1 0 8372 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _288_
timestamp 1638025753
transform 1 0 8372 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_17_100
timestamp 1638025753
transform 1 0 10304 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o41a_2  _296_
timestamp 1638025753
transform 1 0 9384 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__o311a_2  _293_
timestamp 1638025753
transform -1 0 11224 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1638025753
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1638025753
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 1638025753
transform 1 0 12328 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen1
timestamp 1638025753
transform 1 0 12972 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _337_
timestamp 1638025753
transform 1 0 11500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1638025753
transform -1 0 13892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1638025753
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1638025753
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[2\].id.delayenb0
timestamp 1638025753
transform 1 0 1564 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1638025753
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1638025753
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1638025753
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[5\].id.delayenb0
timestamp 1638025753
transform 1 0 3956 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1638025753
transform 1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_49
timestamp 1638025753
transform 1 0 5612 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _334_
timestamp 1638025753
transform -1 0 7268 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_2  _283_
timestamp 1638025753
transform 1 0 5704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_75
timestamp 1638025753
transform 1 0 8004 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1638025753
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_67
timestamp 1638025753
transform 1 0 7268 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1638025753
transform -1 0 8372 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _301_
timestamp 1638025753
transform 1 0 8372 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _343_
timestamp 1638025753
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_94
timestamp 1638025753
transform 1 0 9752 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_2  _295_
timestamp 1638025753
transform 1 0 10028 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 10856 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_112
timestamp 1638025753
transform 1 0 11408 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1638025753
transform -1 0 13432 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[9\].id.delayenb0
timestamp 1638025753
transform 1 0 11500 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1638025753
transform -1 0 13892 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 1638025753
transform 1 0 13432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1638025753
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1638025753
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1638025753
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp 1638025753
transform 1 0 2208 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen1
timestamp 1638025753
transform 1 0 2852 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _346_
timestamp 1638025753
transform 1 0 1380 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[3\].id.delayenb1
timestamp 1638025753
transform 1 0 2116 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  FILLER_20_38
timestamp 1638025753
transform 1 0 4600 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_26
timestamp 1638025753
transform 1 0 3496 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1638025753
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1638025753
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1638025753
transform 1 0 4600 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1638025753
transform 1 0 3128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1638025753
transform 1 0 4876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _342_
timestamp 1638025753
transform -1 0 4600 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _344_
timestamp 1638025753
transform 1 0 3772 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1638025753
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1638025753
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_45
timestamp 1638025753
transform 1 0 5244 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1638025753
transform 1 0 5888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen1
timestamp 1638025753
transform -1 0 5888 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1638025753
transform 1 0 6992 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _340_
timestamp 1638025753
transform -1 0 6256 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_2  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 6992 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[6\].id.delayenb0
timestamp 1638025753
transform 1 0 6256 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_19_87
timestamp 1638025753
transform 1 0 9108 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_68
timestamp 1638025753
transform 1 0 7360 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1638025753
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1638025753
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp 1638025753
transform 1 0 7912 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen1
timestamp 1638025753
transform -1 0 9108 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _339_
timestamp 1638025753
transform -1 0 9936 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[6\].id.delayenb1
timestamp 1638025753
transform -1 0 8464 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1638025753
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_100
timestamp 1638025753
transform 1 0 10304 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_99
timestamp 1638025753
transform 1 0 10212 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1638025753
transform -1 0 10212 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _329_
timestamp 1638025753
transform -1 0 11224 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1638025753
transform 1 0 10396 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _349_
timestamp 1638025753
transform 1 0 9200 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1638025753
transform -1 0 10304 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _292_
timestamp 1638025753
transform 1 0 11500 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1638025753
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1638025753
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_110
timestamp 1638025753
transform 1 0 11224 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_118
timestamp 1638025753
transform 1 0 11960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1638025753
transform 1 0 12788 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1638025753
transform -1 0 12512 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1638025753
transform 1 0 13064 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1638025753
transform 1 0 12512 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[8\].id.delayenb1
timestamp 1638025753
transform 1 0 11500 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[9\].id.delayenb1
timestamp 1638025753
transform 1 0 12512 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_19_135
timestamp 1638025753
transform 1 0 13524 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1638025753
transform -1 0 13892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1638025753
transform -1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_134
timestamp 1638025753
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_21
timestamp 1638025753
transform 1 0 3036 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1638025753
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[3\].id.delayenb0
timestamp 1638025753
transform 1 0 1380 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1638025753
transform 1 0 3128 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[4\].id.delayenb0
timestamp 1638025753
transform 1 0 3496 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1638025753
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1638025753
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1638025753
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _336_
timestamp 1638025753
transform -1 0 7452 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[4\].id.delayenb1
timestamp 1638025753
transform 1 0 5152 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1638025753
transform 1 0 7452 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1638025753
transform 1 0 7636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[7\].id.delayenb0
timestamp 1638025753
transform 1 0 8004 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_21_104
timestamp 1638025753
transform 1 0 10672 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen1
timestamp 1638025753
transform 1 0 10764 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[7\].id.delayenb1
timestamp 1638025753
transform 1 0 9660 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1638025753
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1638025753
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[8\].id.delayenb0
timestamp 1638025753
transform 1 0 11868 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_21_135
timestamp 1638025753
transform 1 0 13524 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1638025753
transform -1 0 13892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1638025753
transform 1 0 1748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1638025753
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1638025753
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp 1638025753
transform 1 0 1840 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen1
timestamp 1638025753
transform 1 0 2484 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1638025753
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_29
timestamp 1638025753
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_42
timestamp 1638025753
transform 1 0 4968 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1638025753
transform 1 0 3128 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1638025753
transform 1 0 4324 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1638025753
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1638025753
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_57
timestamp 1638025753
transform 1 0 6348 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_54
timestamp 1638025753
transform 1 0 6072 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen1
timestamp 1638025753
transform 1 0 5152 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _338_
timestamp 1638025753
transform -1 0 7728 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1638025753
transform 1 0 5796 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_72
timestamp 1638025753
transform 1 0 7728 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1638025753
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1638025753
transform 1 0 8924 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_22_108
timestamp 1638025753
transform 1 0 11040 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen1
timestamp 1638025753
transform 1 0 9568 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _345_
timestamp 1638025753
transform 1 0 10212 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1638025753
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_129
timestamp 1638025753
transform 1 0 12972 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1638025753
transform 1 0 12328 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _347_
timestamp 1638025753
transform 1 0 11500 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_135
timestamp 1638025753
transform 1 0 13524 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1638025753
transform -1 0 13892 0 1 13056
box -38 -48 314 592
<< labels >>
rlabel metal5 s 1104 8210 13892 8530 6 VGND
port 0 nsew ground input
rlabel metal4 s 8208 1040 8528 13648 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 4210 13892 4530 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 12210 13892 12530 6 VPWR
port 1 nsew power input
rlabel metal4 s 4208 1040 4528 13648 6 VPWR
port 1 nsew power input
rlabel metal4 s 12208 1040 12528 13648 6 VPWR
port 1 nsew power input
rlabel metal3 s 0 416 800 536 6 clockp[0]
port 2 nsew signal tristate
rlabel metal3 s 0 1232 800 1352 6 clockp[1]
port 3 nsew signal tristate
rlabel metal3 s 0 7896 800 8016 6 dco
port 4 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 div[0]
port 5 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 div[1]
port 6 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 div[2]
port 7 nsew signal input
rlabel metal3 s 0 5040 800 5160 6 div[3]
port 8 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 div[4]
port 9 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 enable
port 10 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 ext_trim[0]
port 11 nsew signal input
rlabel metal2 s 3974 14200 4030 15000 6 ext_trim[10]
port 12 nsew signal input
rlabel metal2 s 5170 14200 5226 15000 6 ext_trim[11]
port 13 nsew signal input
rlabel metal2 s 6274 14200 6330 15000 6 ext_trim[12]
port 14 nsew signal input
rlabel metal2 s 7470 14200 7526 15000 6 ext_trim[13]
port 15 nsew signal input
rlabel metal2 s 8574 14200 8630 15000 6 ext_trim[14]
port 16 nsew signal input
rlabel metal2 s 9770 14200 9826 15000 6 ext_trim[15]
port 17 nsew signal input
rlabel metal2 s 10874 14200 10930 15000 6 ext_trim[16]
port 18 nsew signal input
rlabel metal2 s 12070 14200 12126 15000 6 ext_trim[17]
port 19 nsew signal input
rlabel metal2 s 13174 14200 13230 15000 6 ext_trim[18]
port 20 nsew signal input
rlabel metal2 s 14370 14200 14426 15000 6 ext_trim[19]
port 21 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 ext_trim[1]
port 22 nsew signal input
rlabel metal3 s 14200 13608 15000 13728 6 ext_trim[20]
port 23 nsew signal input
rlabel metal3 s 14200 11160 15000 11280 6 ext_trim[21]
port 24 nsew signal input
rlabel metal3 s 14200 8712 15000 8832 6 ext_trim[22]
port 25 nsew signal input
rlabel metal3 s 14200 6128 15000 6248 6 ext_trim[23]
port 26 nsew signal input
rlabel metal3 s 14200 3680 15000 3800 6 ext_trim[24]
port 27 nsew signal input
rlabel metal3 s 14200 1232 15000 1352 6 ext_trim[25]
port 28 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 ext_trim[2]
port 29 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 ext_trim[3]
port 30 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 ext_trim[4]
port 31 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 ext_trim[5]
port 32 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 ext_trim[6]
port 33 nsew signal input
rlabel metal2 s 570 14200 626 15000 6 ext_trim[7]
port 34 nsew signal input
rlabel metal2 s 1674 14200 1730 15000 6 ext_trim[8]
port 35 nsew signal input
rlabel metal2 s 2870 14200 2926 15000 6 ext_trim[9]
port 36 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 osc
port 37 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 resetb
port 38 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 15000 15000
<< end >>
