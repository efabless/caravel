magic
tech sky130A
magscale 1 2
timestamp 1636983912
<< locali >>
rect 4721 10455 4755 10557
rect 10057 7259 10091 7361
rect 14013 6987 14047 9673
rect 14105 6917 14139 12053
rect 14013 6883 14139 6917
rect 5089 6647 5123 6749
rect 14013 6103 14047 6883
rect 6929 5627 6963 5865
rect 6101 5015 6135 5185
rect 6009 4539 6043 4709
rect 14013 3043 14047 3893
rect 7941 2839 7975 2941
rect 11805 2499 11839 2601
rect 14013 527 14047 3009
<< viali >>
rect 3157 13481 3191 13515
rect 8585 13481 8619 13515
rect 10885 13481 10919 13515
rect 9689 13413 9723 13447
rect 7665 13345 7699 13379
rect 9137 13345 9171 13379
rect 9229 13345 9263 13379
rect 9873 13345 9907 13379
rect 2421 13277 2455 13311
rect 2973 13277 3007 13311
rect 3157 13277 3191 13311
rect 4445 13277 4479 13311
rect 7205 13277 7239 13311
rect 7389 13277 7423 13311
rect 7757 13277 7791 13311
rect 7849 13277 7883 13311
rect 8125 13277 8159 13311
rect 8309 13277 8343 13311
rect 8401 13277 8435 13311
rect 10333 13277 10367 13311
rect 11621 13277 11655 13311
rect 12081 13277 12115 13311
rect 12725 13277 12759 13311
rect 10425 13209 10459 13243
rect 10517 13209 10551 13243
rect 13185 13209 13219 13243
rect 13277 13209 13311 13243
rect 2605 13141 2639 13175
rect 3341 13141 3375 13175
rect 4629 13141 4663 13175
rect 7941 13141 7975 13175
rect 9321 13141 9355 13175
rect 10701 13141 10735 13175
rect 11713 13141 11747 13175
rect 11989 13141 12023 13175
rect 13369 13141 13403 13175
rect 13461 13141 13495 13175
rect 8677 12937 8711 12971
rect 9413 12937 9447 12971
rect 13369 12937 13403 12971
rect 5733 12869 5767 12903
rect 5825 12869 5859 12903
rect 9321 12869 9355 12903
rect 11161 12869 11195 12903
rect 5549 12801 5583 12835
rect 5922 12801 5956 12835
rect 8769 12801 8803 12835
rect 9597 12801 9631 12835
rect 10517 12801 10551 12835
rect 11529 12801 11563 12835
rect 12449 12801 12483 12835
rect 13185 12801 13219 12835
rect 1593 12733 1627 12767
rect 1869 12733 1903 12767
rect 3341 12733 3375 12767
rect 3617 12733 3651 12767
rect 3893 12733 3927 12767
rect 6377 12733 6411 12767
rect 6653 12733 6687 12767
rect 8125 12733 8159 12767
rect 8585 12733 8619 12767
rect 6101 12665 6135 12699
rect 9137 12665 9171 12699
rect 13001 12665 13035 12699
rect 5365 12597 5399 12631
rect 6653 12393 6687 12427
rect 7665 12393 7699 12427
rect 3893 12325 3927 12359
rect 12173 12325 12207 12359
rect 7757 12257 7791 12291
rect 7941 12257 7975 12291
rect 9045 12257 9079 12291
rect 11713 12257 11747 12291
rect 12265 12257 12299 12291
rect 2421 12189 2455 12223
rect 2789 12189 2823 12223
rect 2972 12189 3006 12223
rect 3065 12189 3099 12223
rect 3157 12189 3191 12223
rect 3341 12189 3375 12223
rect 3985 12189 4019 12223
rect 4169 12189 4203 12223
rect 6285 12189 6319 12223
rect 6469 12189 6503 12223
rect 7295 12189 7329 12223
rect 8217 12189 8251 12223
rect 8329 12189 8363 12223
rect 8953 12189 8987 12223
rect 9229 12189 9263 12223
rect 9505 12189 9539 12223
rect 9597 12189 9631 12223
rect 9873 12189 9907 12223
rect 10609 12189 10643 12223
rect 10977 12189 11011 12223
rect 11437 12189 11471 12223
rect 12541 12189 12575 12223
rect 13185 12189 13219 12223
rect 1501 12121 1535 12155
rect 4445 12121 4479 12155
rect 7849 12121 7883 12155
rect 8769 12121 8803 12155
rect 10793 12121 10827 12155
rect 10885 12121 10919 12155
rect 13461 12121 13495 12155
rect 3433 12053 3467 12087
rect 5917 12053 5951 12087
rect 6101 12053 6135 12087
rect 7113 12053 7147 12087
rect 7297 12053 7331 12087
rect 8493 12053 8527 12087
rect 11621 12053 11655 12087
rect 14105 12053 14139 12087
rect 3433 11849 3467 11883
rect 3617 11849 3651 11883
rect 3709 11849 3743 11883
rect 5457 11849 5491 11883
rect 6745 11849 6779 11883
rect 10517 11849 10551 11883
rect 10793 11849 10827 11883
rect 10977 11849 11011 11883
rect 3157 11781 3191 11815
rect 3525 11781 3559 11815
rect 4537 11781 4571 11815
rect 4629 11781 4663 11815
rect 9229 11781 9263 11815
rect 13277 11781 13311 11815
rect 2605 11713 2639 11747
rect 2881 11713 2915 11747
rect 3249 11713 3283 11747
rect 3893 11713 3927 11747
rect 4393 11713 4427 11747
rect 4813 11713 4847 11747
rect 4905 11713 4939 11747
rect 5411 11713 5445 11747
rect 5917 11713 5951 11747
rect 7021 11713 7055 11747
rect 7297 11713 7331 11747
rect 7941 11713 7975 11747
rect 8217 11713 8251 11747
rect 8584 11713 8618 11747
rect 8677 11713 8711 11747
rect 8769 11713 8803 11747
rect 8953 11713 8987 11747
rect 9413 11713 9447 11747
rect 9965 11713 9999 11747
rect 10609 11713 10643 11747
rect 11069 11713 11103 11747
rect 11529 11713 11563 11747
rect 13001 11713 13035 11747
rect 13461 11713 13495 11747
rect 2513 11645 2547 11679
rect 3065 11645 3099 11679
rect 6909 11645 6943 11679
rect 7389 11645 7423 11679
rect 9045 11645 9079 11679
rect 9689 11645 9723 11679
rect 9873 11645 9907 11679
rect 4261 11577 4295 11611
rect 5825 11577 5859 11611
rect 8309 11577 8343 11611
rect 10333 11577 10367 11611
rect 11253 11577 11287 11611
rect 12817 11577 12851 11611
rect 4997 11509 5031 11543
rect 5273 11509 5307 11543
rect 7573 11509 7607 11543
rect 7849 11509 7883 11543
rect 8125 11509 8159 11543
rect 3433 11305 3467 11339
rect 4077 11305 4111 11339
rect 6285 11305 6319 11339
rect 7113 11305 7147 11339
rect 7757 11305 7791 11339
rect 11529 11305 11563 11339
rect 5549 11237 5583 11271
rect 11161 11237 11195 11271
rect 12357 11237 12391 11271
rect 1501 11169 1535 11203
rect 3249 11169 3283 11203
rect 7941 11169 7975 11203
rect 8309 11169 8343 11203
rect 9137 11169 9171 11203
rect 9321 11169 9355 11203
rect 11713 11169 11747 11203
rect 11897 11169 11931 11203
rect 3341 11101 3375 11135
rect 3801 11101 3835 11135
rect 3985 11101 4019 11135
rect 4261 11101 4295 11135
rect 4537 11101 4571 11135
rect 4721 11101 4755 11135
rect 4997 11101 5031 11135
rect 5417 11101 5451 11135
rect 5733 11101 5767 11135
rect 6106 11101 6140 11135
rect 6683 11101 6717 11135
rect 7205 11101 7239 11135
rect 7573 11101 7607 11135
rect 8125 11101 8159 11135
rect 8401 11101 8435 11135
rect 8494 11101 8528 11135
rect 8677 11101 8711 11135
rect 9413 11101 9447 11135
rect 9873 11101 9907 11135
rect 11069 11101 11103 11135
rect 12541 11101 12575 11135
rect 13461 11101 13495 11135
rect 2973 11033 3007 11067
rect 4813 11033 4847 11067
rect 5181 11033 5215 11067
rect 5273 11033 5307 11067
rect 5917 11033 5951 11067
rect 6009 11033 6043 11067
rect 7297 11033 7331 11067
rect 12449 11033 12483 11067
rect 13185 11033 13219 11067
rect 4537 10965 4571 10999
rect 6561 10965 6595 10999
rect 6745 10965 6779 10999
rect 7389 10965 7423 10999
rect 9781 10965 9815 10999
rect 2237 10761 2271 10795
rect 3249 10761 3283 10795
rect 4077 10761 4111 10795
rect 4353 10761 4387 10795
rect 4445 10761 4479 10795
rect 10333 10761 10367 10795
rect 2605 10693 2639 10727
rect 3525 10693 3559 10727
rect 5457 10693 5491 10727
rect 7113 10693 7147 10727
rect 7757 10693 7791 10727
rect 10149 10693 10183 10727
rect 11069 10693 11103 10727
rect 12449 10693 12483 10727
rect 13185 10693 13219 10727
rect 2053 10625 2087 10659
rect 2421 10625 2455 10659
rect 2697 10625 2731 10659
rect 2841 10625 2875 10659
rect 3433 10625 3467 10659
rect 3622 10625 3656 10659
rect 3709 10625 3743 10659
rect 3893 10625 3927 10659
rect 4261 10625 4295 10659
rect 4905 10625 4939 10659
rect 5089 10625 5123 10659
rect 5733 10625 5767 10659
rect 6469 10625 6503 10659
rect 6745 10625 6779 10659
rect 6929 10625 6963 10659
rect 7389 10625 7423 10659
rect 7665 10625 7699 10659
rect 7849 10625 7883 10659
rect 8033 10625 8067 10659
rect 8401 10625 8435 10659
rect 8493 10625 8527 10659
rect 8861 10625 8895 10659
rect 9137 10625 9171 10659
rect 9523 10625 9557 10659
rect 9689 10625 9723 10659
rect 9781 10625 9815 10659
rect 9965 10625 9999 10659
rect 10609 10625 10643 10659
rect 11529 10625 11563 10659
rect 11805 10625 11839 10659
rect 13553 10625 13587 10659
rect 4629 10557 4663 10591
rect 4721 10557 4755 10591
rect 5641 10557 5675 10591
rect 9321 10557 9355 10591
rect 9413 10557 9447 10591
rect 11161 10557 11195 10591
rect 11897 10557 11931 10591
rect 12725 10557 12759 10591
rect 13277 10557 13311 10591
rect 6561 10489 6595 10523
rect 12633 10489 12667 10523
rect 13369 10489 13403 10523
rect 2973 10421 3007 10455
rect 4721 10421 4755 10455
rect 7941 10421 7975 10455
rect 9045 10421 9079 10455
rect 10517 10421 10551 10455
rect 11713 10421 11747 10455
rect 1501 10217 1535 10251
rect 6929 10217 6963 10251
rect 7941 10217 7975 10251
rect 8769 10217 8803 10251
rect 9505 10217 9539 10251
rect 9781 10217 9815 10251
rect 13185 10217 13219 10251
rect 4077 10149 4111 10183
rect 8493 10149 8527 10183
rect 9965 10149 9999 10183
rect 2973 10081 3007 10115
rect 3249 10081 3283 10115
rect 4261 10081 4295 10115
rect 4813 10081 4847 10115
rect 5457 10081 5491 10115
rect 7113 10081 7147 10115
rect 7205 10081 7239 10115
rect 8033 10081 8067 10115
rect 9321 10081 9355 10115
rect 11805 10081 11839 10115
rect 3893 10013 3927 10047
rect 4077 10013 4111 10047
rect 4445 10013 4479 10047
rect 5181 10013 5215 10047
rect 7515 10013 7549 10047
rect 8217 10013 8251 10047
rect 8585 10013 8619 10047
rect 8953 10013 8987 10047
rect 9229 10013 9263 10047
rect 9597 10013 9631 10047
rect 11713 10013 11747 10047
rect 12357 10013 12391 10047
rect 12449 10013 12483 10047
rect 13277 10013 13311 10047
rect 4721 9945 4755 9979
rect 7757 9945 7791 9979
rect 10793 9945 10827 9979
rect 11069 9945 11103 9979
rect 11897 9945 11931 9979
rect 12909 9945 12943 9979
rect 13001 9945 13035 9979
rect 13461 9945 13495 9979
rect 10057 9877 10091 9911
rect 13369 9877 13403 9911
rect 2145 9673 2179 9707
rect 5549 9673 5583 9707
rect 14013 9673 14047 9707
rect 3709 9605 3743 9639
rect 4077 9605 4111 9639
rect 6193 9605 6227 9639
rect 8585 9605 8619 9639
rect 11253 9605 11287 9639
rect 2329 9537 2363 9571
rect 2973 9537 3007 9571
rect 3156 9537 3190 9571
rect 3341 9537 3375 9571
rect 3525 9537 3559 9571
rect 6009 9537 6043 9571
rect 6377 9537 6411 9571
rect 6837 9537 6871 9571
rect 7205 9537 7239 9571
rect 7481 9537 7515 9571
rect 7665 9537 7699 9571
rect 7757 9537 7791 9571
rect 7901 9537 7935 9571
rect 8677 9537 8711 9571
rect 9137 9537 9171 9571
rect 10057 9537 10091 9571
rect 11621 9537 11655 9571
rect 12633 9537 12667 9571
rect 13461 9537 13495 9571
rect 3249 9469 3283 9503
rect 3801 9469 3835 9503
rect 5825 9469 5859 9503
rect 6561 9469 6595 9503
rect 7113 9469 7147 9503
rect 8493 9469 8527 9503
rect 10793 9469 10827 9503
rect 11345 9469 11379 9503
rect 8033 9401 8067 9435
rect 10425 9401 10459 9435
rect 12909 9401 12943 9435
rect 13277 9401 13311 9435
rect 6469 9333 6503 9367
rect 9045 9333 9079 9367
rect 4905 9129 4939 9163
rect 7021 9129 7055 9163
rect 7481 9129 7515 9163
rect 8401 9129 8435 9163
rect 8677 9129 8711 9163
rect 9229 9129 9263 9163
rect 11529 9129 11563 9163
rect 3157 9061 3191 9095
rect 4537 9061 4571 9095
rect 7297 9061 7331 9095
rect 10701 9061 10735 9095
rect 11621 9061 11655 9095
rect 1685 8993 1719 9027
rect 3893 8993 3927 9027
rect 4353 8993 4387 9027
rect 4997 8993 5031 9027
rect 8033 8993 8067 9027
rect 8217 8993 8251 9027
rect 9689 8993 9723 9027
rect 10149 8993 10183 9027
rect 10885 8993 10919 9027
rect 11069 8993 11103 9027
rect 11805 8993 11839 9027
rect 1409 8925 1443 8959
rect 3801 8925 3835 8959
rect 4169 8925 4203 8959
rect 4445 8925 4479 8959
rect 4721 8925 4755 8959
rect 6929 8925 6963 8959
rect 7941 8925 7975 8959
rect 9505 8925 9539 8959
rect 10241 8925 10275 8959
rect 10517 8925 10551 8959
rect 12173 8925 12207 8959
rect 12817 8925 12851 8959
rect 13369 8925 13403 8959
rect 5273 8857 5307 8891
rect 13093 8857 13127 8891
rect 13185 8857 13219 8891
rect 6745 8789 6779 8823
rect 7573 8789 7607 8823
rect 9597 8789 9631 8823
rect 11161 8789 11195 8823
rect 2513 8585 2547 8619
rect 4261 8585 4295 8619
rect 6101 8585 6135 8619
rect 12633 8585 12667 8619
rect 12817 8585 12851 8619
rect 3433 8517 3467 8551
rect 3893 8517 3927 8551
rect 4169 8517 4203 8551
rect 5181 8517 5215 8551
rect 9413 8517 9447 8551
rect 9505 8517 9539 8551
rect 9781 8517 9815 8551
rect 10977 8517 11011 8551
rect 2053 8449 2087 8483
rect 2329 8449 2363 8483
rect 3157 8449 3191 8483
rect 3341 8449 3375 8483
rect 3577 8449 3611 8483
rect 4077 8449 4111 8483
rect 4629 8449 4663 8483
rect 4905 8449 4939 8483
rect 5089 8449 5123 8483
rect 5325 8449 5359 8483
rect 5917 8449 5951 8483
rect 7481 8449 7515 8483
rect 8677 8449 8711 8483
rect 9229 8449 9263 8483
rect 10425 8449 10459 8483
rect 11345 8449 11379 8483
rect 11713 8449 11747 8483
rect 11897 8449 11931 8483
rect 12541 8449 12575 8483
rect 13185 8449 13219 8483
rect 10517 8381 10551 8415
rect 11069 8381 11103 8415
rect 11989 8381 12023 8415
rect 12449 8381 12483 8415
rect 13277 8381 13311 8415
rect 13369 8381 13403 8415
rect 2237 8313 2271 8347
rect 4813 8313 4847 8347
rect 5457 8313 5491 8347
rect 8769 8313 8803 8347
rect 11161 8313 11195 8347
rect 3709 8245 3743 8279
rect 4445 8245 4479 8279
rect 3157 8041 3191 8075
rect 5549 8041 5583 8075
rect 9137 8041 9171 8075
rect 9505 8041 9539 8075
rect 13461 8041 13495 8075
rect 5825 7973 5859 8007
rect 8309 7973 8343 8007
rect 9597 7973 9631 8007
rect 10517 7973 10551 8007
rect 13093 7973 13127 8007
rect 3801 7905 3835 7939
rect 4077 7905 4111 7939
rect 7665 7905 7699 7939
rect 8401 7905 8435 7939
rect 9689 7905 9723 7939
rect 1409 7837 1443 7871
rect 5917 7837 5951 7871
rect 6561 7837 6595 7871
rect 6745 7837 6779 7871
rect 7205 7837 7239 7871
rect 7849 7837 7883 7871
rect 8677 7837 8711 7871
rect 9413 7837 9447 7871
rect 9781 7837 9815 7871
rect 10195 7837 10229 7871
rect 10793 7837 10827 7871
rect 11529 7837 11563 7871
rect 11805 7837 11839 7871
rect 13185 7837 13219 7871
rect 1685 7769 1719 7803
rect 6929 7769 6963 7803
rect 9965 7769 9999 7803
rect 10333 7769 10367 7803
rect 11713 7769 11747 7803
rect 7021 7701 7055 7735
rect 7573 7701 7607 7735
rect 8493 7701 8527 7735
rect 10149 7701 10183 7735
rect 3416 7497 3450 7531
rect 8585 7497 8619 7531
rect 9413 7497 9447 7531
rect 11069 7497 11103 7531
rect 11989 7497 12023 7531
rect 12449 7497 12483 7531
rect 13001 7497 13035 7531
rect 3709 7429 3743 7463
rect 3801 7429 3835 7463
rect 7297 7429 7331 7463
rect 8125 7429 8159 7463
rect 10701 7429 10735 7463
rect 12357 7429 12391 7463
rect 12909 7429 12943 7463
rect 13185 7429 13219 7463
rect 13369 7429 13403 7463
rect 3565 7361 3599 7395
rect 3985 7361 4019 7395
rect 4445 7361 4479 7395
rect 4610 7361 4644 7395
rect 4813 7361 4847 7395
rect 4997 7361 5031 7395
rect 5641 7361 5675 7395
rect 5825 7361 5859 7395
rect 6009 7361 6043 7395
rect 6745 7361 6779 7395
rect 6837 7361 6871 7395
rect 7481 7361 7515 7395
rect 8401 7361 8435 7395
rect 8769 7361 8803 7395
rect 8861 7361 8895 7395
rect 9045 7361 9079 7395
rect 9873 7361 9907 7395
rect 10057 7361 10091 7395
rect 10241 7361 10275 7395
rect 10425 7361 10459 7395
rect 10517 7361 10551 7395
rect 11805 7361 11839 7395
rect 1409 7293 1443 7327
rect 1685 7293 1719 7327
rect 3157 7293 3191 7327
rect 4721 7293 4755 7327
rect 7389 7293 7423 7327
rect 9597 7293 9631 7327
rect 12633 7293 12667 7327
rect 5733 7225 5767 7259
rect 8953 7225 8987 7259
rect 9781 7225 9815 7259
rect 10057 7225 10091 7259
rect 10333 7225 10367 7259
rect 5089 7157 5123 7191
rect 6653 7157 6687 7191
rect 11345 7157 11379 7191
rect 11621 7157 11655 7191
rect 2329 6953 2363 6987
rect 4813 6953 4847 6987
rect 5720 6953 5754 6987
rect 8493 6953 8527 6987
rect 10977 6953 11011 6987
rect 12265 6953 12299 6987
rect 13553 6953 13587 6987
rect 14013 6953 14047 6987
rect 2421 6885 2455 6919
rect 7205 6885 7239 6919
rect 8953 6885 8987 6919
rect 9597 6885 9631 6919
rect 11529 6885 11563 6919
rect 5457 6817 5491 6851
rect 7849 6817 7883 6851
rect 8033 6817 8067 6851
rect 9505 6817 9539 6851
rect 9689 6817 9723 6851
rect 10425 6817 10459 6851
rect 10517 6817 10551 6851
rect 11621 6817 11655 6851
rect 13001 6817 13035 6851
rect 13093 6817 13127 6851
rect 2145 6749 2179 6783
rect 2605 6749 2639 6783
rect 4072 6749 4106 6783
rect 4445 6749 4479 6783
rect 4813 6749 4847 6783
rect 4997 6749 5031 6783
rect 5089 6749 5123 6783
rect 5365 6749 5399 6783
rect 8401 6749 8435 6783
rect 9321 6749 9355 6783
rect 9781 6749 9815 6783
rect 11069 6749 11103 6783
rect 11713 6749 11747 6783
rect 11897 6749 11931 6783
rect 12357 6749 12391 6783
rect 2789 6681 2823 6715
rect 4169 6681 4203 6715
rect 4261 6681 4295 6715
rect 8217 6681 8251 6715
rect 9137 6681 9171 6715
rect 10057 6681 10091 6715
rect 12909 6681 12943 6715
rect 3885 6613 3919 6647
rect 4629 6613 4663 6647
rect 5089 6613 5123 6647
rect 5273 6613 5307 6647
rect 7389 6613 7423 6647
rect 7757 6613 7791 6647
rect 8769 6613 8803 6647
rect 10609 6613 10643 6647
rect 11989 6613 12023 6647
rect 12541 6613 12575 6647
rect 4905 6409 4939 6443
rect 6009 6409 6043 6443
rect 7849 6409 7883 6443
rect 8861 6409 8895 6443
rect 9781 6409 9815 6443
rect 9965 6409 9999 6443
rect 11897 6409 11931 6443
rect 13277 6409 13311 6443
rect 5733 6341 5767 6375
rect 12541 6341 12575 6375
rect 13185 6341 13219 6375
rect 3433 6273 3467 6307
rect 3617 6273 3651 6307
rect 3893 6273 3927 6307
rect 4123 6273 4157 6307
rect 4629 6273 4663 6307
rect 5089 6273 5123 6307
rect 5181 6273 5215 6307
rect 5365 6273 5399 6307
rect 5513 6273 5547 6307
rect 5641 6273 5675 6307
rect 5871 6273 5905 6307
rect 6377 6273 6411 6307
rect 6653 6273 6687 6307
rect 6745 6273 6779 6307
rect 7297 6273 7331 6307
rect 7481 6273 7515 6307
rect 8217 6273 8251 6307
rect 9045 6273 9079 6307
rect 9321 6273 9355 6307
rect 10425 6273 10459 6307
rect 10701 6273 10735 6307
rect 10793 6273 10827 6307
rect 11161 6273 11195 6307
rect 1409 6205 1443 6239
rect 1685 6205 1719 6239
rect 3709 6205 3743 6239
rect 4261 6205 4295 6239
rect 4353 6205 4387 6239
rect 4741 6205 4775 6239
rect 8309 6205 8343 6239
rect 8493 6205 8527 6239
rect 9229 6205 9263 6239
rect 11345 6205 11379 6239
rect 11989 6205 12023 6239
rect 12081 6205 12115 6239
rect 13369 6205 13403 6239
rect 6929 6137 6963 6171
rect 7113 6137 7147 6171
rect 7665 6137 7699 6171
rect 9141 6137 9175 6171
rect 11529 6137 11563 6171
rect 12725 6137 12759 6171
rect 3157 6069 3191 6103
rect 6469 6069 6503 6103
rect 9505 6069 9539 6103
rect 10057 6069 10091 6103
rect 10333 6069 10367 6103
rect 10977 6069 11011 6103
rect 12817 6069 12851 6103
rect 14013 6069 14047 6103
rect 2237 5865 2271 5899
rect 3893 5865 3927 5899
rect 4261 5865 4295 5899
rect 6101 5865 6135 5899
rect 6745 5865 6779 5899
rect 6929 5865 6963 5899
rect 7205 5865 7239 5899
rect 7849 5865 7883 5899
rect 8033 5865 8067 5899
rect 8217 5865 8251 5899
rect 9597 5865 9631 5899
rect 10517 5865 10551 5899
rect 10701 5865 10735 5899
rect 12265 5865 12299 5899
rect 13461 5865 13495 5899
rect 4537 5797 4571 5831
rect 4905 5797 4939 5831
rect 5365 5797 5399 5831
rect 3985 5729 4019 5763
rect 2053 5661 2087 5695
rect 3157 5661 3191 5695
rect 3617 5661 3651 5695
rect 3893 5661 3927 5695
rect 4721 5661 4755 5695
rect 4813 5661 4847 5695
rect 4997 5661 5031 5695
rect 5497 5661 5531 5695
rect 5917 5661 5951 5695
rect 6377 5661 6411 5695
rect 6561 5661 6595 5695
rect 6653 5661 6687 5695
rect 7481 5797 7515 5831
rect 9321 5797 9355 5831
rect 12449 5797 12483 5831
rect 7757 5729 7791 5763
rect 8401 5729 8435 5763
rect 9229 5729 9263 5763
rect 9965 5729 9999 5763
rect 11345 5729 11379 5763
rect 11621 5729 11655 5763
rect 11805 5729 11839 5763
rect 7113 5661 7147 5695
rect 7849 5661 7883 5695
rect 7941 5661 7975 5695
rect 8493 5661 8527 5695
rect 8953 5661 8987 5695
rect 9137 5661 9171 5695
rect 9413 5661 9447 5695
rect 11897 5661 11931 5695
rect 12541 5661 12575 5695
rect 3525 5593 3559 5627
rect 5641 5593 5675 5627
rect 5733 5593 5767 5627
rect 6009 5593 6043 5627
rect 6929 5593 6963 5627
rect 8217 5593 8251 5627
rect 11161 5593 11195 5627
rect 13001 5593 13035 5627
rect 13093 5593 13127 5627
rect 13277 5593 13311 5627
rect 3249 5525 3283 5559
rect 8677 5525 8711 5559
rect 10057 5525 10091 5559
rect 10149 5525 10183 5559
rect 11069 5525 11103 5559
rect 13185 5525 13219 5559
rect 3157 5321 3191 5355
rect 8953 5321 8987 5355
rect 10149 5321 10183 5355
rect 10977 5321 11011 5355
rect 5641 5253 5675 5287
rect 7297 5253 7331 5287
rect 7665 5253 7699 5287
rect 11529 5253 11563 5287
rect 11897 5253 11931 5287
rect 3801 5185 3835 5219
rect 3893 5185 3927 5219
rect 4169 5185 4203 5219
rect 4261 5185 4295 5219
rect 4445 5185 4479 5219
rect 4537 5185 4571 5219
rect 4630 5185 4664 5219
rect 5273 5185 5307 5219
rect 5457 5185 5491 5219
rect 5825 5185 5859 5219
rect 6009 5185 6043 5219
rect 6101 5185 6135 5219
rect 6653 5185 6687 5219
rect 6745 5185 6779 5219
rect 7113 5185 7147 5219
rect 7481 5185 7515 5219
rect 7757 5185 7791 5219
rect 8217 5185 8251 5219
rect 8677 5185 8711 5219
rect 9229 5185 9263 5219
rect 9505 5185 9539 5219
rect 9965 5185 9999 5219
rect 10333 5185 10367 5219
rect 10517 5185 10551 5219
rect 10609 5185 10643 5219
rect 1409 5117 1443 5151
rect 1685 5117 1719 5151
rect 5549 5117 5583 5151
rect 4905 5049 4939 5083
rect 10790 5175 10824 5209
rect 11345 5185 11379 5219
rect 11713 5185 11747 5219
rect 11989 5185 12023 5219
rect 12909 5185 12943 5219
rect 6837 5117 6871 5151
rect 6929 5117 6963 5151
rect 7849 5117 7883 5151
rect 11253 5117 11287 5151
rect 8493 5049 8527 5083
rect 8585 5049 8619 5083
rect 9689 5049 9723 5083
rect 10425 5049 10459 5083
rect 13277 5049 13311 5083
rect 3617 4981 3651 5015
rect 4077 4981 4111 5015
rect 6101 4981 6135 5015
rect 6469 4981 6503 5015
rect 8401 4981 8435 5015
rect 9597 4981 9631 5015
rect 9781 4981 9815 5015
rect 11161 4981 11195 5015
rect 2237 4777 2271 4811
rect 2513 4777 2547 4811
rect 2973 4777 3007 4811
rect 4537 4777 4571 4811
rect 6193 4777 6227 4811
rect 7849 4777 7883 4811
rect 10793 4777 10827 4811
rect 13369 4777 13403 4811
rect 6009 4709 6043 4743
rect 8769 4709 8803 4743
rect 9689 4709 9723 4743
rect 11529 4709 11563 4743
rect 3065 4641 3099 4675
rect 3985 4641 4019 4675
rect 5256 4641 5290 4675
rect 5549 4641 5583 4675
rect 2053 4573 2087 4607
rect 2697 4573 2731 4607
rect 2789 4573 2823 4607
rect 3433 4573 3467 4607
rect 3617 4573 3651 4607
rect 5457 4573 5491 4607
rect 6377 4641 6411 4675
rect 7021 4641 7055 4675
rect 9045 4641 9079 4675
rect 10425 4641 10459 4675
rect 11069 4641 11103 4675
rect 6469 4573 6503 4607
rect 6565 4573 6599 4607
rect 6653 4573 6687 4607
rect 6837 4573 6871 4607
rect 7205 4573 7239 4607
rect 7389 4573 7423 4607
rect 7481 4573 7515 4607
rect 7757 4573 7791 4607
rect 8401 4573 8435 4607
rect 8585 4573 8619 4607
rect 9321 4573 9355 4607
rect 9965 4573 9999 4607
rect 10149 4573 10183 4607
rect 10333 4573 10367 4607
rect 10517 4573 10551 4607
rect 10609 4573 10643 4607
rect 11713 4573 11747 4607
rect 12449 4573 12483 4607
rect 12633 4573 12667 4607
rect 12909 4573 12943 4607
rect 13185 4573 13219 4607
rect 3249 4505 3283 4539
rect 4813 4505 4847 4539
rect 4997 4505 5031 4539
rect 5341 4505 5375 4539
rect 6009 4505 6043 4539
rect 11621 4505 11655 4539
rect 4077 4437 4111 4471
rect 4169 4437 4203 4471
rect 7573 4437 7607 4471
rect 9229 4437 9263 4471
rect 9873 4437 9907 4471
rect 12725 4437 12759 4471
rect 13093 4437 13127 4471
rect 3525 4233 3559 4267
rect 11161 4233 11195 4267
rect 3893 4165 3927 4199
rect 4537 4165 4571 4199
rect 4629 4165 4663 4199
rect 5457 4165 5491 4199
rect 5549 4165 5583 4199
rect 6101 4165 6135 4199
rect 10517 4165 10551 4199
rect 10701 4165 10735 4199
rect 3341 4097 3375 4131
rect 3663 4097 3697 4131
rect 4440 4097 4474 4131
rect 4813 4097 4847 4131
rect 5181 4097 5215 4131
rect 5329 4097 5363 4131
rect 5687 4097 5721 4131
rect 6193 4097 6227 4131
rect 6377 4097 6411 4131
rect 6653 4097 6687 4131
rect 7849 4097 7883 4131
rect 9229 4097 9263 4131
rect 9413 4097 9447 4131
rect 9965 4097 9999 4131
rect 10057 4097 10091 4131
rect 10241 4097 10275 4131
rect 10425 4097 10459 4131
rect 11253 4097 11287 4131
rect 12173 4097 12207 4131
rect 13277 4097 13311 4131
rect 1409 4029 1443 4063
rect 1685 4029 1719 4063
rect 3433 4029 3467 4063
rect 6469 4029 6503 4063
rect 8217 4029 8251 4063
rect 11621 4029 11655 4063
rect 12449 4029 12483 4063
rect 13001 4029 13035 4063
rect 3893 3961 3927 3995
rect 9597 3961 9631 3995
rect 10149 3961 10183 3995
rect 12081 3961 12115 3995
rect 12909 3961 12943 3995
rect 13093 3961 13127 3995
rect 3157 3893 3191 3927
rect 4261 3893 4295 3927
rect 5825 3893 5859 3927
rect 8769 3893 8803 3927
rect 9045 3893 9079 3927
rect 9781 3893 9815 3927
rect 10701 3893 10735 3927
rect 10885 3893 10919 3927
rect 12265 3893 12299 3927
rect 13553 3893 13587 3927
rect 14013 3893 14047 3927
rect 1593 3689 1627 3723
rect 2421 3689 2455 3723
rect 3065 3689 3099 3723
rect 3341 3689 3375 3723
rect 5917 3689 5951 3723
rect 9413 3689 9447 3723
rect 5181 3621 5215 3655
rect 7481 3621 7515 3655
rect 9505 3621 9539 3655
rect 9597 3621 9631 3655
rect 10609 3621 10643 3655
rect 13277 3621 13311 3655
rect 6377 3553 6411 3587
rect 7021 3553 7055 3587
rect 1777 3485 1811 3519
rect 2237 3485 2271 3519
rect 3157 3485 3191 3519
rect 3617 3485 3651 3519
rect 5181 3485 5215 3519
rect 5365 3485 5399 3519
rect 5549 3485 5583 3519
rect 6101 3485 6135 3519
rect 6193 3485 6227 3519
rect 6469 3485 6503 3519
rect 7849 3485 7883 3519
rect 8401 3485 8435 3519
rect 8769 3485 8803 3519
rect 9321 3485 9355 3519
rect 9731 3485 9765 3519
rect 10425 3485 10459 3519
rect 10517 3485 10551 3519
rect 10701 3485 10735 3519
rect 10977 3485 11011 3519
rect 11989 3485 12023 3519
rect 12909 3485 12943 3519
rect 3433 3417 3467 3451
rect 7573 3417 7607 3451
rect 8033 3417 8067 3451
rect 11713 3417 11747 3451
rect 11897 3417 11931 3451
rect 7665 3349 7699 3383
rect 7941 3349 7975 3383
rect 8309 3349 8343 3383
rect 8493 3349 8527 3383
rect 8585 3349 8619 3383
rect 8953 3349 8987 3383
rect 9965 3349 9999 3383
rect 10241 3349 10275 3383
rect 2881 3145 2915 3179
rect 5365 3145 5399 3179
rect 8033 3145 8067 3179
rect 8401 3145 8435 3179
rect 8493 3145 8527 3179
rect 9873 3145 9907 3179
rect 11253 3145 11287 3179
rect 11897 3145 11931 3179
rect 12541 3145 12575 3179
rect 13461 3145 13495 3179
rect 3525 3077 3559 3111
rect 3893 3077 3927 3111
rect 7573 3077 7607 3111
rect 9045 3077 9079 3111
rect 13369 3077 13403 3111
rect 2513 3009 2547 3043
rect 3019 3009 3053 3043
rect 3157 3009 3191 3043
rect 5825 3009 5859 3043
rect 6837 3009 6871 3043
rect 7757 3009 7791 3043
rect 9229 3009 9263 3043
rect 9413 3009 9447 3043
rect 10609 3009 10643 3043
rect 10701 3009 10735 3043
rect 10885 3009 10919 3043
rect 11069 3009 11103 3043
rect 12909 3009 12943 3043
rect 13001 3009 13035 3043
rect 14013 3009 14047 3043
rect 3433 2941 3467 2975
rect 3617 2941 3651 2975
rect 7941 2941 7975 2975
rect 8585 2941 8619 2975
rect 9597 2941 9631 2975
rect 9781 2941 9815 2975
rect 11989 2941 12023 2975
rect 12081 2941 12115 2975
rect 13093 2941 13127 2975
rect 8861 2873 8895 2907
rect 10425 2873 10459 2907
rect 10793 2873 10827 2907
rect 11529 2873 11563 2907
rect 2697 2805 2731 2839
rect 6009 2805 6043 2839
rect 6377 2805 6411 2839
rect 7941 2805 7975 2839
rect 10241 2805 10275 2839
rect 12449 2805 12483 2839
rect 3341 2601 3375 2635
rect 4629 2601 4663 2635
rect 6653 2601 6687 2635
rect 9137 2601 9171 2635
rect 10517 2601 10551 2635
rect 11805 2601 11839 2635
rect 7481 2533 7515 2567
rect 8125 2533 8159 2567
rect 13461 2533 13495 2567
rect 1593 2465 1627 2499
rect 1869 2465 1903 2499
rect 5181 2465 5215 2499
rect 7021 2465 7055 2499
rect 7573 2465 7607 2499
rect 8769 2465 8803 2499
rect 10241 2465 10275 2499
rect 10977 2465 11011 2499
rect 11713 2465 11747 2499
rect 11805 2465 11839 2499
rect 11989 2465 12023 2499
rect 4169 2397 4203 2431
rect 4445 2397 4479 2431
rect 4905 2397 4939 2431
rect 7665 2397 7699 2431
rect 8033 2397 8067 2431
rect 10057 2397 10091 2431
rect 11161 2397 11195 2431
rect 12265 2397 12299 2431
rect 12725 2397 12759 2431
rect 8309 2329 8343 2363
rect 9321 2329 9355 2363
rect 9505 2329 9539 2363
rect 10609 2329 10643 2363
rect 10793 2329 10827 2363
rect 11621 2329 11655 2363
rect 13185 2329 13219 2363
rect 13277 2329 13311 2363
rect 4353 2261 4387 2295
rect 6837 2261 6871 2295
rect 8033 2261 8067 2295
rect 9597 2261 9631 2295
rect 9965 2261 9999 2295
rect 12173 2261 12207 2295
rect 12633 2261 12667 2295
rect 13369 2261 13403 2295
rect 5549 2057 5583 2091
rect 8953 2057 8987 2091
rect 10977 2057 11011 2091
rect 11345 2057 11379 2091
rect 6193 1989 6227 2023
rect 6837 1989 6871 2023
rect 9965 1989 9999 2023
rect 13277 1989 13311 2023
rect 1409 1921 1443 1955
rect 5181 1921 5215 1955
rect 5487 1921 5521 1955
rect 6009 1921 6043 1955
rect 6469 1921 6503 1955
rect 6653 1921 6687 1955
rect 7205 1921 7239 1955
rect 7297 1921 7331 1955
rect 8769 1921 8803 1955
rect 9321 1921 9355 1955
rect 10241 1921 10275 1955
rect 10517 1921 10551 1955
rect 11529 1921 11563 1955
rect 13001 1921 13035 1955
rect 1685 1853 1719 1887
rect 3157 1853 3191 1887
rect 4905 1853 4939 1887
rect 10701 1853 10735 1887
rect 10885 1853 10919 1887
rect 13461 1853 13495 1887
rect 3433 1785 3467 1819
rect 5917 1785 5951 1819
rect 8585 1785 8619 1819
rect 12817 1785 12851 1819
rect 5365 1717 5399 1751
rect 7021 1717 7055 1751
rect 10333 1717 10367 1751
rect 2237 1513 2271 1547
rect 3433 1513 3467 1547
rect 10517 1513 10551 1547
rect 10793 1513 10827 1547
rect 11805 1513 11839 1547
rect 12173 1513 12207 1547
rect 13369 1513 13403 1547
rect 7573 1445 7607 1479
rect 8585 1445 8619 1479
rect 10241 1445 10275 1479
rect 5365 1377 5399 1411
rect 5825 1377 5859 1411
rect 8677 1377 8711 1411
rect 9505 1377 9539 1411
rect 10333 1377 10367 1411
rect 10977 1377 11011 1411
rect 2053 1309 2087 1343
rect 3249 1309 3283 1343
rect 5641 1309 5675 1343
rect 6009 1309 6043 1343
rect 6193 1309 6227 1343
rect 7021 1309 7055 1343
rect 7757 1309 7791 1343
rect 7941 1309 7975 1343
rect 8125 1309 8159 1343
rect 9781 1309 9815 1343
rect 10701 1309 10735 1343
rect 11713 1309 11747 1343
rect 12357 1309 12391 1343
rect 13093 1309 13127 1343
rect 13277 1309 13311 1343
rect 13553 1309 13587 1343
rect 3525 1241 3559 1275
rect 6469 1241 6503 1275
rect 9321 1241 9355 1275
rect 3893 1173 3927 1207
rect 8953 1173 8987 1207
rect 9413 1173 9447 1207
rect 14013 493 14047 527
<< metal1 >>
rect 1104 13626 13892 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 12214 13626
rect 12266 13574 12278 13626
rect 12330 13574 12342 13626
rect 12394 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 13892 13626
rect 1104 13552 13892 13574
rect 3142 13512 3148 13524
rect 3103 13484 3148 13512
rect 3142 13472 3148 13484
rect 3200 13472 3206 13524
rect 8202 13472 8208 13524
rect 8260 13512 8266 13524
rect 8573 13515 8631 13521
rect 8573 13512 8585 13515
rect 8260 13484 8585 13512
rect 8260 13472 8266 13484
rect 8573 13481 8585 13484
rect 8619 13481 8631 13515
rect 9766 13512 9772 13524
rect 8573 13475 8631 13481
rect 9508 13484 9772 13512
rect 6730 13404 6736 13456
rect 6788 13444 6794 13456
rect 6788 13416 9260 13444
rect 6788 13404 6794 13416
rect 7653 13379 7711 13385
rect 7653 13345 7665 13379
rect 7699 13376 7711 13379
rect 7926 13376 7932 13388
rect 7699 13348 7932 13376
rect 7699 13345 7711 13348
rect 7653 13339 7711 13345
rect 7926 13336 7932 13348
rect 7984 13336 7990 13388
rect 9232 13385 9260 13416
rect 9125 13379 9183 13385
rect 9125 13345 9137 13379
rect 9171 13345 9183 13379
rect 9125 13339 9183 13345
rect 9217 13379 9275 13385
rect 9217 13345 9229 13379
rect 9263 13376 9275 13379
rect 9398 13376 9404 13388
rect 9263 13348 9404 13376
rect 9263 13345 9275 13348
rect 9217 13339 9275 13345
rect 2038 13268 2044 13320
rect 2096 13308 2102 13320
rect 2409 13311 2467 13317
rect 2409 13308 2421 13311
rect 2096 13280 2421 13308
rect 2096 13268 2102 13280
rect 2409 13277 2421 13280
rect 2455 13277 2467 13311
rect 2409 13271 2467 13277
rect 2682 13268 2688 13320
rect 2740 13308 2746 13320
rect 2961 13311 3019 13317
rect 2961 13308 2973 13311
rect 2740 13280 2973 13308
rect 2740 13268 2746 13280
rect 2961 13277 2973 13280
rect 3007 13277 3019 13311
rect 2961 13271 3019 13277
rect 3145 13311 3203 13317
rect 3145 13277 3157 13311
rect 3191 13308 3203 13311
rect 3326 13308 3332 13320
rect 3191 13280 3332 13308
rect 3191 13277 3203 13280
rect 3145 13271 3203 13277
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 4433 13311 4491 13317
rect 4433 13277 4445 13311
rect 4479 13308 4491 13311
rect 6086 13308 6092 13320
rect 4479 13280 6092 13308
rect 4479 13277 4491 13280
rect 4433 13271 4491 13277
rect 6086 13268 6092 13280
rect 6144 13268 6150 13320
rect 6914 13268 6920 13320
rect 6972 13308 6978 13320
rect 7193 13311 7251 13317
rect 7193 13308 7205 13311
rect 6972 13280 7205 13308
rect 6972 13268 6978 13280
rect 7193 13277 7205 13280
rect 7239 13277 7251 13311
rect 7374 13308 7380 13320
rect 7335 13280 7380 13308
rect 7193 13271 7251 13277
rect 7208 13240 7236 13271
rect 7374 13268 7380 13280
rect 7432 13268 7438 13320
rect 7742 13308 7748 13320
rect 7703 13280 7748 13308
rect 7742 13268 7748 13280
rect 7800 13268 7806 13320
rect 7834 13268 7840 13320
rect 7892 13308 7898 13320
rect 8113 13311 8171 13317
rect 7892 13280 7937 13308
rect 7892 13268 7898 13280
rect 8113 13277 8125 13311
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 8297 13311 8355 13317
rect 8297 13277 8309 13311
rect 8343 13277 8355 13311
rect 8297 13271 8355 13277
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13308 8447 13311
rect 8570 13308 8576 13320
rect 8435 13280 8576 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 8128 13240 8156 13271
rect 7208 13212 8156 13240
rect 8312 13240 8340 13271
rect 8570 13268 8576 13280
rect 8628 13268 8634 13320
rect 9140 13308 9168 13339
rect 9398 13336 9404 13348
rect 9456 13336 9462 13388
rect 9508 13308 9536 13484
rect 9766 13472 9772 13484
rect 9824 13512 9830 13524
rect 10870 13512 10876 13524
rect 9824 13484 10876 13512
rect 9824 13472 9830 13484
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 9582 13404 9588 13456
rect 9640 13444 9646 13456
rect 9677 13447 9735 13453
rect 9677 13444 9689 13447
rect 9640 13416 9689 13444
rect 9640 13404 9646 13416
rect 9677 13413 9689 13416
rect 9723 13444 9735 13447
rect 9723 13416 9904 13444
rect 9723 13413 9735 13416
rect 9677 13407 9735 13413
rect 9876 13385 9904 13416
rect 9861 13379 9919 13385
rect 9861 13345 9873 13379
rect 9907 13345 9919 13379
rect 9861 13339 9919 13345
rect 9140 13280 9536 13308
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 11146 13308 11152 13320
rect 10367 13280 11152 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 11146 13268 11152 13280
rect 11204 13308 11210 13320
rect 11609 13311 11667 13317
rect 11609 13308 11621 13311
rect 11204 13280 11621 13308
rect 11204 13268 11210 13280
rect 11609 13277 11621 13280
rect 11655 13277 11667 13311
rect 12066 13308 12072 13320
rect 12027 13280 12072 13308
rect 11609 13271 11667 13277
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 12618 13268 12624 13320
rect 12676 13308 12682 13320
rect 12713 13311 12771 13317
rect 12713 13308 12725 13311
rect 12676 13280 12725 13308
rect 12676 13268 12682 13280
rect 12713 13277 12725 13280
rect 12759 13277 12771 13311
rect 12713 13271 12771 13277
rect 8754 13240 8760 13252
rect 8312 13212 8760 13240
rect 8036 13184 8064 13212
rect 8754 13200 8760 13212
rect 8812 13200 8818 13252
rect 10413 13243 10471 13249
rect 10413 13209 10425 13243
rect 10459 13240 10471 13243
rect 10505 13243 10563 13249
rect 10505 13240 10517 13243
rect 10459 13212 10517 13240
rect 10459 13209 10471 13212
rect 10413 13203 10471 13209
rect 10505 13209 10517 13212
rect 10551 13209 10563 13243
rect 13170 13240 13176 13252
rect 13131 13212 13176 13240
rect 10505 13203 10563 13209
rect 13170 13200 13176 13212
rect 13228 13200 13234 13252
rect 13262 13200 13268 13252
rect 13320 13240 13326 13252
rect 13320 13212 13365 13240
rect 13320 13200 13326 13212
rect 2590 13172 2596 13184
rect 2551 13144 2596 13172
rect 2590 13132 2596 13144
rect 2648 13132 2654 13184
rect 3329 13175 3387 13181
rect 3329 13141 3341 13175
rect 3375 13172 3387 13175
rect 3602 13172 3608 13184
rect 3375 13144 3608 13172
rect 3375 13141 3387 13144
rect 3329 13135 3387 13141
rect 3602 13132 3608 13144
rect 3660 13132 3666 13184
rect 4614 13172 4620 13184
rect 4575 13144 4620 13172
rect 4614 13132 4620 13144
rect 4672 13132 4678 13184
rect 7742 13132 7748 13184
rect 7800 13172 7806 13184
rect 7929 13175 7987 13181
rect 7929 13172 7941 13175
rect 7800 13144 7941 13172
rect 7800 13132 7806 13144
rect 7929 13141 7941 13144
rect 7975 13141 7987 13175
rect 7929 13135 7987 13141
rect 8018 13132 8024 13184
rect 8076 13132 8082 13184
rect 9306 13132 9312 13184
rect 9364 13172 9370 13184
rect 10686 13172 10692 13184
rect 9364 13144 9409 13172
rect 10647 13144 10692 13172
rect 9364 13132 9370 13144
rect 10686 13132 10692 13144
rect 10744 13132 10750 13184
rect 11698 13172 11704 13184
rect 11659 13144 11704 13172
rect 11698 13132 11704 13144
rect 11756 13132 11762 13184
rect 11974 13172 11980 13184
rect 11935 13144 11980 13172
rect 11974 13132 11980 13144
rect 12032 13132 12038 13184
rect 13188 13172 13216 13200
rect 13357 13175 13415 13181
rect 13357 13172 13369 13175
rect 13188 13144 13369 13172
rect 13357 13141 13369 13144
rect 13403 13141 13415 13175
rect 13357 13135 13415 13141
rect 13446 13132 13452 13184
rect 13504 13172 13510 13184
rect 13504 13144 13549 13172
rect 13504 13132 13510 13144
rect 1104 13082 13892 13104
rect 1104 13030 8214 13082
rect 8266 13030 8278 13082
rect 8330 13030 8342 13082
rect 8394 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 13892 13082
rect 1104 13008 13892 13030
rect 7374 12968 7380 12980
rect 3988 12940 7380 12968
rect 3988 12912 4016 12940
rect 2590 12860 2596 12912
rect 2648 12860 2654 12912
rect 3970 12900 3976 12912
rect 3344 12872 3976 12900
rect 1581 12767 1639 12773
rect 1581 12733 1593 12767
rect 1627 12764 1639 12767
rect 1854 12764 1860 12776
rect 1627 12736 1716 12764
rect 1815 12736 1860 12764
rect 1627 12733 1639 12736
rect 1581 12727 1639 12733
rect 1688 12628 1716 12736
rect 1854 12724 1860 12736
rect 1912 12724 1918 12776
rect 3344 12773 3372 12872
rect 3970 12860 3976 12872
rect 4028 12860 4034 12912
rect 4614 12860 4620 12912
rect 4672 12860 4678 12912
rect 5736 12909 5764 12940
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 8110 12928 8116 12980
rect 8168 12968 8174 12980
rect 8665 12971 8723 12977
rect 8665 12968 8677 12971
rect 8168 12940 8677 12968
rect 8168 12928 8174 12940
rect 8665 12937 8677 12940
rect 8711 12937 8723 12971
rect 9398 12968 9404 12980
rect 9359 12940 9404 12968
rect 8665 12931 8723 12937
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 13262 12928 13268 12980
rect 13320 12968 13326 12980
rect 13357 12971 13415 12977
rect 13357 12968 13369 12971
rect 13320 12940 13369 12968
rect 13320 12928 13326 12940
rect 13357 12937 13369 12940
rect 13403 12937 13415 12971
rect 13357 12931 13415 12937
rect 5721 12903 5779 12909
rect 5721 12869 5733 12903
rect 5767 12869 5779 12903
rect 5721 12863 5779 12869
rect 5813 12903 5871 12909
rect 5813 12869 5825 12903
rect 5859 12900 5871 12903
rect 6914 12900 6920 12912
rect 5859 12872 6920 12900
rect 5859 12869 5871 12872
rect 5813 12863 5871 12869
rect 6914 12860 6920 12872
rect 6972 12860 6978 12912
rect 7098 12860 7104 12912
rect 7156 12860 7162 12912
rect 9309 12903 9367 12909
rect 9309 12900 9321 12903
rect 8588 12872 9321 12900
rect 5537 12835 5595 12841
rect 5537 12801 5549 12835
rect 5583 12801 5595 12835
rect 5537 12795 5595 12801
rect 3329 12767 3387 12773
rect 3329 12733 3341 12767
rect 3375 12733 3387 12767
rect 3329 12727 3387 12733
rect 3510 12724 3516 12776
rect 3568 12764 3574 12776
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 3568 12736 3617 12764
rect 3568 12724 3574 12736
rect 3605 12733 3617 12736
rect 3651 12733 3663 12767
rect 3605 12727 3663 12733
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12764 3939 12767
rect 3970 12764 3976 12776
rect 3927 12736 3976 12764
rect 3927 12733 3939 12736
rect 3881 12727 3939 12733
rect 3970 12724 3976 12736
rect 4028 12724 4034 12776
rect 4890 12724 4896 12776
rect 4948 12764 4954 12776
rect 5552 12764 5580 12795
rect 5626 12792 5632 12844
rect 5684 12832 5690 12844
rect 5910 12835 5968 12841
rect 5910 12832 5922 12835
rect 5684 12804 5922 12832
rect 5684 12792 5690 12804
rect 5910 12801 5922 12804
rect 5956 12801 5968 12835
rect 5910 12795 5968 12801
rect 4948 12736 5580 12764
rect 4948 12724 4954 12736
rect 5718 12724 5724 12776
rect 5776 12764 5782 12776
rect 6365 12767 6423 12773
rect 6365 12764 6377 12767
rect 5776 12736 6377 12764
rect 5776 12724 5782 12736
rect 6365 12733 6377 12736
rect 6411 12733 6423 12767
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 6365 12727 6423 12733
rect 6472 12736 6653 12764
rect 6089 12699 6147 12705
rect 6089 12665 6101 12699
rect 6135 12696 6147 12699
rect 6472 12696 6500 12736
rect 6641 12733 6653 12736
rect 6687 12733 6699 12767
rect 6641 12727 6699 12733
rect 8018 12724 8024 12776
rect 8076 12764 8082 12776
rect 8588 12773 8616 12872
rect 9309 12869 9321 12872
rect 9355 12900 9367 12903
rect 9766 12900 9772 12912
rect 9355 12872 9772 12900
rect 9355 12869 9367 12872
rect 9309 12863 9367 12869
rect 9766 12860 9772 12872
rect 9824 12860 9830 12912
rect 11146 12900 11152 12912
rect 11107 12872 11152 12900
rect 11146 12860 11152 12872
rect 11204 12860 11210 12912
rect 8757 12835 8815 12841
rect 8757 12801 8769 12835
rect 8803 12832 8815 12835
rect 8846 12832 8852 12844
rect 8803 12804 8852 12832
rect 8803 12801 8815 12804
rect 8757 12795 8815 12801
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 9582 12832 9588 12844
rect 9543 12804 9588 12832
rect 9582 12792 9588 12804
rect 9640 12792 9646 12844
rect 10502 12832 10508 12844
rect 10463 12804 10508 12832
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 8113 12767 8171 12773
rect 8113 12764 8125 12767
rect 8076 12736 8125 12764
rect 8076 12724 8082 12736
rect 8113 12733 8125 12736
rect 8159 12733 8171 12767
rect 8113 12727 8171 12733
rect 8573 12767 8631 12773
rect 8573 12733 8585 12767
rect 8619 12733 8631 12767
rect 11532 12764 11560 12795
rect 11698 12792 11704 12844
rect 11756 12832 11762 12844
rect 12437 12835 12495 12841
rect 12437 12832 12449 12835
rect 11756 12804 12449 12832
rect 11756 12792 11762 12804
rect 12437 12801 12449 12804
rect 12483 12832 12495 12835
rect 13173 12835 13231 12841
rect 13173 12832 13185 12835
rect 12483 12804 13185 12832
rect 12483 12801 12495 12804
rect 12437 12795 12495 12801
rect 13173 12801 13185 12804
rect 13219 12832 13231 12835
rect 13354 12832 13360 12844
rect 13219 12804 13360 12832
rect 13219 12801 13231 12804
rect 13173 12795 13231 12801
rect 13354 12792 13360 12804
rect 13412 12792 13418 12844
rect 8573 12727 8631 12733
rect 9140 12736 11744 12764
rect 9140 12705 9168 12736
rect 11716 12708 11744 12736
rect 6135 12668 6500 12696
rect 9125 12699 9183 12705
rect 6135 12665 6147 12668
rect 6089 12659 6147 12665
rect 9125 12665 9137 12699
rect 9171 12665 9183 12699
rect 9125 12659 9183 12665
rect 11698 12656 11704 12708
rect 11756 12656 11762 12708
rect 12989 12699 13047 12705
rect 12989 12665 13001 12699
rect 13035 12696 13047 12699
rect 13262 12696 13268 12708
rect 13035 12668 13268 12696
rect 13035 12665 13047 12668
rect 12989 12659 13047 12665
rect 13262 12656 13268 12668
rect 13320 12656 13326 12708
rect 3510 12628 3516 12640
rect 1688 12600 3516 12628
rect 3510 12588 3516 12600
rect 3568 12588 3574 12640
rect 5350 12628 5356 12640
rect 5311 12600 5356 12628
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 1104 12538 13892 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 12214 12538
rect 12266 12486 12278 12538
rect 12330 12486 12342 12538
rect 12394 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 13892 12538
rect 1104 12464 13892 12486
rect 6641 12427 6699 12433
rect 2516 12396 6592 12424
rect 2516 12288 2544 12396
rect 2682 12316 2688 12368
rect 2740 12356 2746 12368
rect 2958 12356 2964 12368
rect 2740 12328 2964 12356
rect 2740 12316 2746 12328
rect 2958 12316 2964 12328
rect 3016 12356 3022 12368
rect 3881 12359 3939 12365
rect 3881 12356 3893 12359
rect 3016 12328 3893 12356
rect 3016 12316 3022 12328
rect 3881 12325 3893 12328
rect 3927 12325 3939 12359
rect 6564 12356 6592 12396
rect 6641 12393 6653 12427
rect 6687 12424 6699 12427
rect 7098 12424 7104 12436
rect 6687 12396 7104 12424
rect 6687 12393 6699 12396
rect 6641 12387 6699 12393
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 7653 12427 7711 12433
rect 7653 12393 7665 12427
rect 7699 12424 7711 12427
rect 8570 12424 8576 12436
rect 7699 12396 8576 12424
rect 7699 12393 7711 12396
rect 7653 12387 7711 12393
rect 8570 12384 8576 12396
rect 8628 12384 8634 12436
rect 9674 12384 9680 12436
rect 9732 12424 9738 12436
rect 9858 12424 9864 12436
rect 9732 12396 9864 12424
rect 9732 12384 9738 12396
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 11974 12356 11980 12368
rect 6564 12328 11980 12356
rect 3881 12319 3939 12325
rect 11974 12316 11980 12328
rect 12032 12316 12038 12368
rect 12066 12316 12072 12368
rect 12124 12356 12130 12368
rect 12161 12359 12219 12365
rect 12161 12356 12173 12359
rect 12124 12328 12173 12356
rect 12124 12316 12130 12328
rect 12161 12325 12173 12328
rect 12207 12356 12219 12359
rect 13262 12356 13268 12368
rect 12207 12328 13268 12356
rect 12207 12325 12219 12328
rect 12161 12319 12219 12325
rect 13262 12316 13268 12328
rect 13320 12316 13326 12368
rect 2424 12260 2544 12288
rect 2424 12229 2452 12260
rect 2866 12248 2872 12300
rect 2924 12288 2930 12300
rect 4522 12288 4528 12300
rect 2924 12260 4528 12288
rect 2924 12248 2930 12260
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12189 2467 12223
rect 2409 12183 2467 12189
rect 2682 12180 2688 12232
rect 2740 12220 2746 12232
rect 2976 12229 3004 12260
rect 4522 12248 4528 12260
rect 4580 12248 4586 12300
rect 7742 12288 7748 12300
rect 7703 12260 7748 12288
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 7926 12288 7932 12300
rect 7887 12260 7932 12288
rect 7926 12248 7932 12260
rect 7984 12288 7990 12300
rect 8754 12288 8760 12300
rect 7984 12260 8248 12288
rect 7984 12248 7990 12260
rect 2777 12223 2835 12229
rect 2777 12220 2789 12223
rect 2740 12192 2789 12220
rect 2740 12180 2746 12192
rect 2777 12189 2789 12192
rect 2823 12189 2835 12223
rect 2777 12183 2835 12189
rect 2960 12223 3018 12229
rect 2960 12189 2972 12223
rect 3006 12189 3018 12223
rect 2960 12183 3018 12189
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12189 3111 12223
rect 3053 12183 3111 12189
rect 1486 12152 1492 12164
rect 1447 12124 1492 12152
rect 1486 12112 1492 12124
rect 1544 12112 1550 12164
rect 3068 12152 3096 12183
rect 3142 12180 3148 12232
rect 3200 12220 3206 12232
rect 3329 12223 3387 12229
rect 3200 12192 3245 12220
rect 3200 12180 3206 12192
rect 3329 12189 3341 12223
rect 3375 12220 3387 12223
rect 3418 12220 3424 12232
rect 3375 12192 3424 12220
rect 3375 12189 3387 12192
rect 3329 12183 3387 12189
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12220 4031 12223
rect 4062 12220 4068 12232
rect 4019 12192 4068 12220
rect 4019 12189 4031 12192
rect 3973 12183 4031 12189
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12189 4215 12223
rect 4157 12183 4215 12189
rect 3234 12152 3240 12164
rect 3068 12124 3240 12152
rect 3234 12112 3240 12124
rect 3292 12112 3298 12164
rect 3510 12112 3516 12164
rect 3568 12152 3574 12164
rect 4172 12152 4200 12183
rect 6086 12180 6092 12232
rect 6144 12220 6150 12232
rect 6273 12223 6331 12229
rect 6273 12220 6285 12223
rect 6144 12192 6285 12220
rect 6144 12180 6150 12192
rect 6273 12189 6285 12192
rect 6319 12220 6331 12223
rect 6457 12223 6515 12229
rect 6457 12220 6469 12223
rect 6319 12192 6469 12220
rect 6319 12189 6331 12192
rect 6273 12183 6331 12189
rect 6457 12189 6469 12192
rect 6503 12189 6515 12223
rect 6457 12183 6515 12189
rect 7283 12223 7341 12229
rect 7283 12189 7295 12223
rect 7329 12220 7341 12223
rect 7374 12220 7380 12232
rect 7329 12192 7380 12220
rect 7329 12189 7341 12192
rect 7283 12183 7341 12189
rect 7374 12180 7380 12192
rect 7432 12180 7438 12232
rect 8220 12229 8248 12260
rect 8404 12260 8760 12288
rect 8205 12223 8263 12229
rect 8205 12189 8217 12223
rect 8251 12189 8263 12223
rect 8317 12223 8375 12229
rect 8317 12220 8329 12223
rect 8205 12183 8263 12189
rect 8312 12189 8329 12220
rect 8363 12220 8375 12223
rect 8404 12220 8432 12260
rect 8754 12248 8760 12260
rect 8812 12248 8818 12300
rect 9030 12288 9036 12300
rect 8991 12260 9036 12288
rect 9030 12248 9036 12260
rect 9088 12248 9094 12300
rect 11698 12288 11704 12300
rect 9232 12260 11100 12288
rect 11659 12260 11704 12288
rect 9232 12229 9260 12260
rect 8941 12223 8999 12229
rect 8941 12220 8953 12223
rect 8363 12192 8432 12220
rect 8496 12192 8953 12220
rect 8363 12189 8375 12192
rect 8312 12183 8375 12189
rect 4430 12152 4436 12164
rect 3568 12124 4200 12152
rect 4391 12124 4436 12152
rect 3568 12112 3574 12124
rect 3421 12087 3479 12093
rect 3421 12053 3433 12087
rect 3467 12084 3479 12087
rect 3786 12084 3792 12096
rect 3467 12056 3792 12084
rect 3467 12053 3479 12056
rect 3421 12047 3479 12053
rect 3786 12044 3792 12056
rect 3844 12044 3850 12096
rect 4172 12084 4200 12124
rect 4430 12112 4436 12124
rect 4488 12112 4494 12164
rect 5658 12124 6132 12152
rect 5718 12084 5724 12096
rect 4172 12056 5724 12084
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 5902 12084 5908 12096
rect 5863 12056 5908 12084
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 6104 12093 6132 12124
rect 6914 12112 6920 12164
rect 6972 12152 6978 12164
rect 7837 12155 7895 12161
rect 7837 12152 7849 12155
rect 6972 12124 7849 12152
rect 6972 12112 6978 12124
rect 7837 12121 7849 12124
rect 7883 12152 7895 12155
rect 8312 12152 8340 12183
rect 7883 12124 8340 12152
rect 7883 12121 7895 12124
rect 7837 12115 7895 12121
rect 6089 12087 6147 12093
rect 6089 12053 6101 12087
rect 6135 12053 6147 12087
rect 6089 12047 6147 12053
rect 7006 12044 7012 12096
rect 7064 12084 7070 12096
rect 7101 12087 7159 12093
rect 7101 12084 7113 12087
rect 7064 12056 7113 12084
rect 7064 12044 7070 12056
rect 7101 12053 7113 12056
rect 7147 12053 7159 12087
rect 7101 12047 7159 12053
rect 7285 12087 7343 12093
rect 7285 12053 7297 12087
rect 7331 12084 7343 12087
rect 8018 12084 8024 12096
rect 7331 12056 8024 12084
rect 7331 12053 7343 12056
rect 7285 12047 7343 12053
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 8496 12093 8524 12192
rect 8941 12189 8953 12192
rect 8987 12189 8999 12223
rect 8941 12183 8999 12189
rect 9217 12223 9275 12229
rect 9217 12189 9229 12223
rect 9263 12189 9275 12223
rect 9217 12183 9275 12189
rect 9493 12223 9551 12229
rect 9493 12189 9505 12223
rect 9539 12189 9551 12223
rect 9493 12183 9551 12189
rect 8570 12112 8576 12164
rect 8628 12152 8634 12164
rect 8757 12155 8815 12161
rect 8757 12152 8769 12155
rect 8628 12124 8769 12152
rect 8628 12112 8634 12124
rect 8757 12121 8769 12124
rect 8803 12152 8815 12155
rect 9232 12152 9260 12183
rect 8803 12124 9260 12152
rect 9508 12152 9536 12183
rect 9582 12180 9588 12232
rect 9640 12220 9646 12232
rect 9861 12223 9919 12229
rect 9640 12192 9685 12220
rect 9640 12180 9646 12192
rect 9861 12189 9873 12223
rect 9907 12220 9919 12223
rect 9950 12220 9956 12232
rect 9907 12192 9956 12220
rect 9907 12189 9919 12192
rect 9861 12183 9919 12189
rect 9950 12180 9956 12192
rect 10008 12180 10014 12232
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12220 10655 12223
rect 10686 12220 10692 12232
rect 10643 12192 10692 12220
rect 10643 12189 10655 12192
rect 10597 12183 10655 12189
rect 10686 12180 10692 12192
rect 10744 12220 10750 12232
rect 10965 12223 11023 12229
rect 10965 12220 10977 12223
rect 10744 12192 10977 12220
rect 10744 12180 10750 12192
rect 10965 12189 10977 12192
rect 11011 12189 11023 12223
rect 10965 12183 11023 12189
rect 9674 12152 9680 12164
rect 9508 12124 9680 12152
rect 8803 12121 8815 12124
rect 8757 12115 8815 12121
rect 9674 12112 9680 12124
rect 9732 12112 9738 12164
rect 10502 12112 10508 12164
rect 10560 12152 10566 12164
rect 10781 12155 10839 12161
rect 10781 12152 10793 12155
rect 10560 12124 10793 12152
rect 10560 12112 10566 12124
rect 10781 12121 10793 12124
rect 10827 12121 10839 12155
rect 10781 12115 10839 12121
rect 8481 12087 8539 12093
rect 8481 12053 8493 12087
rect 8527 12084 8539 12087
rect 8662 12084 8668 12096
rect 8527 12056 8668 12084
rect 8527 12053 8539 12056
rect 8481 12047 8539 12053
rect 8662 12044 8668 12056
rect 8720 12044 8726 12096
rect 10796 12084 10824 12115
rect 10870 12112 10876 12164
rect 10928 12152 10934 12164
rect 11072 12152 11100 12260
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 12253 12291 12311 12297
rect 12253 12257 12265 12291
rect 12299 12288 12311 12291
rect 13446 12288 13452 12300
rect 12299 12260 13452 12288
rect 12299 12257 12311 12260
rect 12253 12251 12311 12257
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 11422 12220 11428 12232
rect 11383 12192 11428 12220
rect 11422 12180 11428 12192
rect 11480 12180 11486 12232
rect 12529 12223 12587 12229
rect 12529 12189 12541 12223
rect 12575 12220 12587 12223
rect 12618 12220 12624 12232
rect 12575 12192 12624 12220
rect 12575 12189 12587 12192
rect 12529 12183 12587 12189
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 13170 12220 13176 12232
rect 13131 12192 13176 12220
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 10928 12124 10973 12152
rect 11072 12124 11652 12152
rect 10928 12112 10934 12124
rect 11624 12096 11652 12124
rect 10962 12084 10968 12096
rect 10796 12056 10968 12084
rect 10962 12044 10968 12056
rect 11020 12044 11026 12096
rect 11606 12084 11612 12096
rect 11567 12056 11612 12084
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 12636 12084 12664 12180
rect 13354 12112 13360 12164
rect 13412 12152 13418 12164
rect 13449 12155 13507 12161
rect 13449 12152 13461 12155
rect 13412 12124 13461 12152
rect 13412 12112 13418 12124
rect 13449 12121 13461 12124
rect 13495 12121 13507 12155
rect 13449 12115 13507 12121
rect 14093 12087 14151 12093
rect 14093 12084 14105 12087
rect 12636 12056 14105 12084
rect 14093 12053 14105 12056
rect 14139 12053 14151 12087
rect 14093 12047 14151 12053
rect 1104 11994 13892 12016
rect 1104 11942 8214 11994
rect 8266 11942 8278 11994
rect 8330 11942 8342 11994
rect 8394 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 13892 11994
rect 1104 11920 13892 11942
rect 1854 11840 1860 11892
rect 1912 11880 1918 11892
rect 3421 11883 3479 11889
rect 3421 11880 3433 11883
rect 1912 11852 3433 11880
rect 1912 11840 1918 11852
rect 3421 11849 3433 11852
rect 3467 11849 3479 11883
rect 3602 11880 3608 11892
rect 3515 11852 3608 11880
rect 3421 11843 3479 11849
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 3697 11883 3755 11889
rect 3697 11849 3709 11883
rect 3743 11880 3755 11883
rect 5445 11883 5503 11889
rect 5445 11880 5457 11883
rect 3743 11852 4384 11880
rect 3743 11849 3755 11852
rect 3697 11843 3755 11849
rect 3050 11812 3056 11824
rect 2884 11784 3056 11812
rect 2593 11747 2651 11753
rect 2593 11713 2605 11747
rect 2639 11744 2651 11747
rect 2774 11744 2780 11756
rect 2639 11716 2780 11744
rect 2639 11713 2651 11716
rect 2593 11707 2651 11713
rect 2774 11704 2780 11716
rect 2832 11704 2838 11756
rect 2884 11753 2912 11784
rect 3050 11772 3056 11784
rect 3108 11772 3114 11824
rect 3145 11815 3203 11821
rect 3145 11781 3157 11815
rect 3191 11812 3203 11815
rect 3513 11815 3571 11821
rect 3513 11812 3525 11815
rect 3191 11784 3525 11812
rect 3191 11781 3203 11784
rect 3145 11775 3203 11781
rect 3513 11781 3525 11784
rect 3559 11781 3571 11815
rect 3513 11775 3571 11781
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11713 2927 11747
rect 2869 11707 2927 11713
rect 2958 11704 2964 11756
rect 3016 11744 3022 11756
rect 3237 11747 3295 11753
rect 3237 11744 3249 11747
rect 3016 11716 3249 11744
rect 3016 11704 3022 11716
rect 3237 11713 3249 11716
rect 3283 11713 3295 11747
rect 3237 11707 3295 11713
rect 2501 11679 2559 11685
rect 2501 11645 2513 11679
rect 2547 11676 2559 11679
rect 3053 11679 3111 11685
rect 3053 11676 3065 11679
rect 2547 11648 3065 11676
rect 2547 11645 2559 11648
rect 2501 11639 2559 11645
rect 3053 11645 3065 11648
rect 3099 11676 3111 11679
rect 3326 11676 3332 11688
rect 3099 11648 3332 11676
rect 3099 11645 3111 11648
rect 3053 11639 3111 11645
rect 3326 11636 3332 11648
rect 3384 11636 3390 11688
rect 3620 11676 3648 11840
rect 4356 11756 4384 11852
rect 4540 11852 5457 11880
rect 4540 11821 4568 11852
rect 5445 11849 5457 11852
rect 5491 11849 5503 11883
rect 5445 11843 5503 11849
rect 4525 11815 4583 11821
rect 4525 11781 4537 11815
rect 4571 11781 4583 11815
rect 4525 11775 4583 11781
rect 4614 11772 4620 11824
rect 4672 11812 4678 11824
rect 5460 11812 5488 11843
rect 5902 11840 5908 11892
rect 5960 11840 5966 11892
rect 6733 11883 6791 11889
rect 6733 11849 6745 11883
rect 6779 11880 6791 11883
rect 10505 11883 10563 11889
rect 6779 11852 9168 11880
rect 6779 11849 6791 11852
rect 6733 11843 6791 11849
rect 5920 11812 5948 11840
rect 4672 11784 5120 11812
rect 5460 11784 6132 11812
rect 4672 11772 4678 11784
rect 3878 11744 3884 11756
rect 3839 11716 3884 11744
rect 3878 11704 3884 11716
rect 3936 11704 3942 11756
rect 4338 11704 4344 11756
rect 4396 11753 4402 11756
rect 4396 11747 4439 11753
rect 4427 11713 4439 11747
rect 4798 11744 4804 11756
rect 4759 11716 4804 11744
rect 4396 11707 4439 11713
rect 4396 11704 4402 11707
rect 4798 11704 4804 11716
rect 4856 11704 4862 11756
rect 4893 11747 4951 11753
rect 4893 11713 4905 11747
rect 4939 11713 4951 11747
rect 5092 11744 5120 11784
rect 5350 11744 5356 11756
rect 5092 11716 5356 11744
rect 4893 11707 4951 11713
rect 4908 11676 4936 11707
rect 5350 11704 5356 11716
rect 5408 11753 5414 11756
rect 5408 11747 5457 11753
rect 5408 11713 5411 11747
rect 5445 11744 5457 11747
rect 5905 11747 5963 11753
rect 5905 11744 5917 11747
rect 5445 11716 5917 11744
rect 5445 11713 5457 11716
rect 5408 11707 5457 11713
rect 5905 11713 5917 11716
rect 5951 11744 5963 11747
rect 5994 11744 6000 11756
rect 5951 11716 6000 11744
rect 5951 11713 5963 11716
rect 5905 11707 5963 11713
rect 5408 11704 5414 11707
rect 5994 11704 6000 11716
rect 6052 11704 6058 11756
rect 3620 11648 4936 11676
rect 4249 11611 4307 11617
rect 4249 11577 4261 11611
rect 4295 11608 4307 11611
rect 4430 11608 4436 11620
rect 4295 11580 4436 11608
rect 4295 11577 4307 11580
rect 4249 11571 4307 11577
rect 4430 11568 4436 11580
rect 4488 11568 4494 11620
rect 5166 11568 5172 11620
rect 5224 11608 5230 11620
rect 5813 11611 5871 11617
rect 5224 11580 5488 11608
rect 5224 11568 5230 11580
rect 4982 11540 4988 11552
rect 4943 11512 4988 11540
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 5258 11540 5264 11552
rect 5219 11512 5264 11540
rect 5258 11500 5264 11512
rect 5316 11500 5322 11552
rect 5460 11540 5488 11580
rect 5813 11577 5825 11611
rect 5859 11608 5871 11611
rect 6104 11608 6132 11784
rect 8110 11772 8116 11824
rect 8168 11812 8174 11824
rect 9030 11812 9036 11824
rect 8168 11784 9036 11812
rect 8168 11772 8174 11784
rect 7006 11744 7012 11756
rect 6967 11716 7012 11744
rect 7006 11704 7012 11716
rect 7064 11744 7070 11756
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 7064 11716 7297 11744
rect 7064 11704 7070 11716
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11744 7987 11747
rect 8205 11747 8263 11753
rect 7975 11716 8064 11744
rect 7975 11713 7987 11716
rect 7929 11707 7987 11713
rect 6897 11679 6955 11685
rect 6897 11645 6909 11679
rect 6943 11676 6955 11679
rect 7374 11676 7380 11688
rect 6943 11648 7380 11676
rect 6943 11645 6955 11648
rect 6897 11639 6955 11645
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 8036 11620 8064 11716
rect 8205 11713 8217 11747
rect 8251 11713 8263 11747
rect 8205 11707 8263 11713
rect 8220 11676 8248 11707
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 8956 11753 8984 11784
rect 9030 11772 9036 11784
rect 9088 11772 9094 11824
rect 8572 11747 8630 11753
rect 8572 11744 8584 11747
rect 8536 11716 8584 11744
rect 8536 11704 8542 11716
rect 8572 11713 8584 11716
rect 8618 11713 8630 11747
rect 8572 11707 8630 11713
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 8757 11747 8815 11753
rect 8757 11713 8769 11747
rect 8803 11713 8815 11747
rect 8757 11707 8815 11713
rect 8941 11747 8999 11753
rect 8941 11713 8953 11747
rect 8987 11713 8999 11747
rect 9140 11744 9168 11852
rect 10505 11849 10517 11883
rect 10551 11880 10563 11883
rect 10686 11880 10692 11892
rect 10551 11852 10692 11880
rect 10551 11849 10563 11852
rect 10505 11843 10563 11849
rect 9217 11815 9275 11821
rect 9217 11781 9229 11815
rect 9263 11812 9275 11815
rect 9674 11812 9680 11824
rect 9263 11784 9680 11812
rect 9263 11781 9275 11784
rect 9217 11775 9275 11781
rect 9674 11772 9680 11784
rect 9732 11812 9738 11824
rect 10520 11812 10548 11843
rect 10686 11840 10692 11852
rect 10744 11840 10750 11892
rect 10781 11883 10839 11889
rect 10781 11849 10793 11883
rect 10827 11849 10839 11883
rect 10962 11880 10968 11892
rect 10923 11852 10968 11880
rect 10781 11843 10839 11849
rect 9732 11784 10548 11812
rect 9732 11772 9738 11784
rect 9401 11747 9459 11753
rect 9401 11744 9413 11747
rect 9140 11716 9413 11744
rect 8941 11707 8999 11713
rect 9401 11713 9413 11716
rect 9447 11744 9459 11747
rect 9582 11744 9588 11756
rect 9447 11716 9588 11744
rect 9447 11713 9459 11716
rect 9401 11707 9459 11713
rect 8220 11648 8616 11676
rect 7926 11608 7932 11620
rect 5859 11580 6132 11608
rect 7576 11580 7932 11608
rect 5859 11577 5871 11580
rect 5813 11571 5871 11577
rect 7576 11549 7604 11580
rect 7926 11568 7932 11580
rect 7984 11568 7990 11620
rect 8018 11568 8024 11620
rect 8076 11608 8082 11620
rect 8297 11611 8355 11617
rect 8297 11608 8309 11611
rect 8076 11580 8309 11608
rect 8076 11568 8082 11580
rect 8297 11577 8309 11580
rect 8343 11577 8355 11611
rect 8297 11571 8355 11577
rect 7561 11543 7619 11549
rect 7561 11540 7573 11543
rect 5460 11512 7573 11540
rect 7561 11509 7573 11512
rect 7607 11509 7619 11543
rect 7834 11540 7840 11552
rect 7795 11512 7840 11540
rect 7561 11503 7619 11509
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 8113 11543 8171 11549
rect 8113 11509 8125 11543
rect 8159 11540 8171 11543
rect 8202 11540 8208 11552
rect 8159 11512 8208 11540
rect 8159 11509 8171 11512
rect 8113 11503 8171 11509
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8588 11540 8616 11648
rect 8680 11620 8708 11707
rect 8772 11676 8800 11707
rect 9582 11704 9588 11716
rect 9640 11704 9646 11756
rect 9766 11744 9772 11756
rect 9692 11716 9772 11744
rect 9692 11685 9720 11716
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11744 10011 11747
rect 10134 11744 10140 11756
rect 9999 11716 10140 11744
rect 9999 11713 10011 11716
rect 9953 11707 10011 11713
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 10502 11704 10508 11756
rect 10560 11744 10566 11756
rect 10597 11747 10655 11753
rect 10597 11744 10609 11747
rect 10560 11716 10609 11744
rect 10560 11704 10566 11716
rect 10597 11713 10609 11716
rect 10643 11713 10655 11747
rect 10796 11744 10824 11843
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 13262 11812 13268 11824
rect 13223 11784 13268 11812
rect 13262 11772 13268 11784
rect 13320 11772 13326 11824
rect 10870 11744 10876 11756
rect 10796 11716 10876 11744
rect 10597 11707 10655 11713
rect 10870 11704 10876 11716
rect 10928 11704 10934 11756
rect 11054 11744 11060 11756
rect 11015 11716 11060 11744
rect 11054 11704 11060 11716
rect 11112 11704 11118 11756
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 12989 11747 13047 11753
rect 12989 11713 13001 11747
rect 13035 11744 13047 11747
rect 13446 11744 13452 11756
rect 13035 11716 13452 11744
rect 13035 11713 13047 11716
rect 12989 11707 13047 11713
rect 9033 11679 9091 11685
rect 9033 11676 9045 11679
rect 8772 11648 9045 11676
rect 8662 11568 8668 11620
rect 8720 11568 8726 11620
rect 8772 11540 8800 11648
rect 9033 11645 9045 11648
rect 9079 11645 9091 11679
rect 9033 11639 9091 11645
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11645 9735 11679
rect 9858 11676 9864 11688
rect 9819 11648 9864 11676
rect 9677 11639 9735 11645
rect 9858 11636 9864 11648
rect 9916 11636 9922 11688
rect 11532 11676 11560 11707
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 11882 11676 11888 11688
rect 10336 11648 11888 11676
rect 10336 11617 10364 11648
rect 11882 11636 11888 11648
rect 11940 11636 11946 11688
rect 10321 11611 10379 11617
rect 10321 11577 10333 11611
rect 10367 11577 10379 11611
rect 10321 11571 10379 11577
rect 10778 11568 10784 11620
rect 10836 11608 10842 11620
rect 11241 11611 11299 11617
rect 11241 11608 11253 11611
rect 10836 11580 11253 11608
rect 10836 11568 10842 11580
rect 11241 11577 11253 11580
rect 11287 11577 11299 11611
rect 12802 11608 12808 11620
rect 12763 11580 12808 11608
rect 11241 11571 11299 11577
rect 12802 11568 12808 11580
rect 12860 11568 12866 11620
rect 8588 11512 8800 11540
rect 9950 11500 9956 11552
rect 10008 11540 10014 11552
rect 10962 11540 10968 11552
rect 10008 11512 10968 11540
rect 10008 11500 10014 11512
rect 10962 11500 10968 11512
rect 11020 11540 11026 11552
rect 11422 11540 11428 11552
rect 11020 11512 11428 11540
rect 11020 11500 11026 11512
rect 11422 11500 11428 11512
rect 11480 11500 11486 11552
rect 1104 11450 13892 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 12214 11450
rect 12266 11398 12278 11450
rect 12330 11398 12342 11450
rect 12394 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 13892 11450
rect 1104 11376 13892 11398
rect 3142 11296 3148 11348
rect 3200 11336 3206 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 3200 11308 3433 11336
rect 3200 11296 3206 11308
rect 3421 11305 3433 11308
rect 3467 11305 3479 11339
rect 3421 11299 3479 11305
rect 3326 11268 3332 11280
rect 3252 11240 3332 11268
rect 1489 11203 1547 11209
rect 1489 11169 1501 11203
rect 1535 11200 1547 11203
rect 2590 11200 2596 11212
rect 1535 11172 2596 11200
rect 1535 11169 1547 11172
rect 1489 11163 1547 11169
rect 2590 11160 2596 11172
rect 2648 11160 2654 11212
rect 3252 11209 3280 11240
rect 3326 11228 3332 11240
rect 3384 11228 3390 11280
rect 3237 11203 3295 11209
rect 3237 11169 3249 11203
rect 3283 11169 3295 11203
rect 3436 11200 3464 11299
rect 3970 11296 3976 11348
rect 4028 11336 4034 11348
rect 4065 11339 4123 11345
rect 4065 11336 4077 11339
rect 4028 11308 4077 11336
rect 4028 11296 4034 11308
rect 4065 11305 4077 11308
rect 4111 11305 4123 11339
rect 4065 11299 4123 11305
rect 6273 11339 6331 11345
rect 6273 11305 6285 11339
rect 6319 11336 6331 11339
rect 6914 11336 6920 11348
rect 6319 11308 6920 11336
rect 6319 11305 6331 11308
rect 6273 11299 6331 11305
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 7006 11296 7012 11348
rect 7064 11336 7070 11348
rect 7101 11339 7159 11345
rect 7101 11336 7113 11339
rect 7064 11308 7113 11336
rect 7064 11296 7070 11308
rect 7101 11305 7113 11308
rect 7147 11305 7159 11339
rect 7101 11299 7159 11305
rect 7374 11296 7380 11348
rect 7432 11336 7438 11348
rect 7745 11339 7803 11345
rect 7745 11336 7757 11339
rect 7432 11308 7757 11336
rect 7432 11296 7438 11308
rect 7745 11305 7757 11308
rect 7791 11305 7803 11339
rect 7745 11299 7803 11305
rect 7926 11296 7932 11348
rect 7984 11336 7990 11348
rect 7984 11308 9260 11336
rect 7984 11296 7990 11308
rect 5442 11228 5448 11280
rect 5500 11268 5506 11280
rect 5537 11271 5595 11277
rect 5537 11268 5549 11271
rect 5500 11240 5549 11268
rect 5500 11228 5506 11240
rect 5537 11237 5549 11240
rect 5583 11237 5595 11271
rect 5537 11231 5595 11237
rect 5828 11240 6132 11268
rect 3436 11172 4292 11200
rect 3237 11163 3295 11169
rect 3326 11092 3332 11144
rect 3384 11132 3390 11144
rect 3786 11132 3792 11144
rect 3384 11104 3429 11132
rect 3747 11104 3792 11132
rect 3384 11092 3390 11104
rect 3786 11092 3792 11104
rect 3844 11092 3850 11144
rect 3878 11092 3884 11144
rect 3936 11132 3942 11144
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3936 11104 3985 11132
rect 3936 11092 3942 11104
rect 3973 11101 3985 11104
rect 4019 11132 4031 11135
rect 4062 11132 4068 11144
rect 4019 11104 4068 11132
rect 4019 11101 4031 11104
rect 3973 11095 4031 11101
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 4264 11141 4292 11172
rect 4338 11160 4344 11212
rect 4396 11200 4402 11212
rect 4396 11172 4936 11200
rect 4396 11160 4402 11172
rect 4908 11144 4936 11172
rect 5258 11160 5264 11212
rect 5316 11200 5322 11212
rect 5316 11172 5764 11200
rect 5316 11160 5322 11172
rect 4249 11135 4307 11141
rect 4249 11101 4261 11135
rect 4295 11101 4307 11135
rect 4249 11095 4307 11101
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11132 4583 11135
rect 4614 11132 4620 11144
rect 4571 11104 4620 11132
rect 4571 11101 4583 11104
rect 4525 11095 4583 11101
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 4706 11092 4712 11144
rect 4764 11132 4770 11144
rect 4764 11104 4809 11132
rect 4764 11092 4770 11104
rect 4890 11092 4896 11144
rect 4948 11132 4954 11144
rect 4985 11135 5043 11141
rect 4985 11132 4997 11135
rect 4948 11104 4997 11132
rect 4948 11092 4954 11104
rect 4985 11101 4997 11104
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 5405 11135 5463 11141
rect 5405 11101 5417 11135
rect 5451 11132 5463 11135
rect 5626 11132 5632 11144
rect 5451 11104 5632 11132
rect 5451 11101 5463 11104
rect 5405 11095 5463 11101
rect 5626 11092 5632 11104
rect 5684 11092 5690 11144
rect 5736 11141 5764 11172
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11101 5779 11135
rect 5721 11095 5779 11101
rect 2222 11024 2228 11076
rect 2280 11024 2286 11076
rect 2958 11064 2964 11076
rect 2919 11036 2964 11064
rect 2958 11024 2964 11036
rect 3016 11024 3022 11076
rect 4632 11064 4660 11092
rect 4801 11067 4859 11073
rect 4801 11064 4813 11067
rect 4632 11036 4813 11064
rect 4801 11033 4813 11036
rect 4847 11033 4859 11067
rect 5166 11064 5172 11076
rect 5127 11036 5172 11064
rect 4801 11027 4859 11033
rect 5166 11024 5172 11036
rect 5224 11024 5230 11076
rect 5261 11067 5319 11073
rect 5261 11033 5273 11067
rect 5307 11064 5319 11067
rect 5828 11064 5856 11240
rect 5902 11160 5908 11212
rect 5960 11160 5966 11212
rect 6104 11200 6132 11240
rect 7834 11228 7840 11280
rect 7892 11268 7898 11280
rect 7892 11240 8524 11268
rect 7892 11228 7898 11240
rect 6104 11172 6224 11200
rect 5920 11132 5948 11160
rect 6094 11135 6152 11141
rect 6094 11132 6106 11135
rect 5920 11104 6106 11132
rect 6094 11101 6106 11104
rect 6140 11101 6152 11135
rect 6094 11095 6152 11101
rect 5307 11036 5856 11064
rect 5905 11067 5963 11073
rect 5307 11033 5319 11036
rect 5261 11027 5319 11033
rect 5905 11033 5917 11067
rect 5951 11033 5963 11067
rect 5905 11027 5963 11033
rect 750 10956 756 11008
rect 808 10996 814 11008
rect 2774 10996 2780 11008
rect 808 10968 2780 10996
rect 808 10956 814 10968
rect 2774 10956 2780 10968
rect 2832 10956 2838 11008
rect 3326 10956 3332 11008
rect 3384 10996 3390 11008
rect 4246 10996 4252 11008
rect 3384 10968 4252 10996
rect 3384 10956 3390 10968
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 4525 10999 4583 11005
rect 4525 10965 4537 10999
rect 4571 10996 4583 10999
rect 4890 10996 4896 11008
rect 4571 10968 4896 10996
rect 4571 10965 4583 10968
rect 4525 10959 4583 10965
rect 4890 10956 4896 10968
rect 4948 10996 4954 11008
rect 5920 10996 5948 11027
rect 5994 11024 6000 11076
rect 6052 11064 6058 11076
rect 6196 11064 6224 11172
rect 7098 11160 7104 11212
rect 7156 11200 7162 11212
rect 7929 11203 7987 11209
rect 7929 11200 7941 11203
rect 7156 11172 7941 11200
rect 7156 11160 7162 11172
rect 7929 11169 7941 11172
rect 7975 11169 7987 11203
rect 7929 11163 7987 11169
rect 8202 11160 8208 11212
rect 8260 11200 8266 11212
rect 8297 11203 8355 11209
rect 8297 11200 8309 11203
rect 8260 11172 8309 11200
rect 8260 11160 8266 11172
rect 8297 11169 8309 11172
rect 8343 11169 8355 11203
rect 8297 11163 8355 11169
rect 6546 11092 6552 11144
rect 6604 11132 6610 11144
rect 6671 11135 6729 11141
rect 6671 11132 6683 11135
rect 6604 11104 6683 11132
rect 6604 11092 6610 11104
rect 6671 11101 6683 11104
rect 6717 11132 6729 11135
rect 7006 11132 7012 11144
rect 6717 11104 7012 11132
rect 6717 11101 6729 11104
rect 6671 11095 6729 11101
rect 7006 11092 7012 11104
rect 7064 11092 7070 11144
rect 7190 11132 7196 11144
rect 7151 11104 7196 11132
rect 7190 11092 7196 11104
rect 7248 11132 7254 11144
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 7248 11104 7573 11132
rect 7248 11092 7254 11104
rect 7561 11101 7573 11104
rect 7607 11101 7619 11135
rect 8110 11132 8116 11144
rect 8071 11104 8116 11132
rect 7561 11095 7619 11101
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 8496 11141 8524 11240
rect 9125 11203 9183 11209
rect 9125 11169 9137 11203
rect 9171 11169 9183 11203
rect 9232 11200 9260 11308
rect 9858 11296 9864 11348
rect 9916 11336 9922 11348
rect 11517 11339 11575 11345
rect 11517 11336 11529 11339
rect 9916 11308 11529 11336
rect 9916 11296 9922 11308
rect 11517 11305 11529 11308
rect 11563 11305 11575 11339
rect 11517 11299 11575 11305
rect 11054 11228 11060 11280
rect 11112 11268 11118 11280
rect 11149 11271 11207 11277
rect 11149 11268 11161 11271
rect 11112 11240 11161 11268
rect 11112 11228 11118 11240
rect 11149 11237 11161 11240
rect 11195 11237 11207 11271
rect 11149 11231 11207 11237
rect 12345 11271 12403 11277
rect 12345 11237 12357 11271
rect 12391 11268 12403 11271
rect 12434 11268 12440 11280
rect 12391 11240 12440 11268
rect 12391 11237 12403 11240
rect 12345 11231 12403 11237
rect 12434 11228 12440 11240
rect 12492 11268 12498 11280
rect 12802 11268 12808 11280
rect 12492 11240 12808 11268
rect 12492 11228 12498 11240
rect 12802 11228 12808 11240
rect 12860 11228 12866 11280
rect 9309 11203 9367 11209
rect 9309 11200 9321 11203
rect 9232 11172 9321 11200
rect 9125 11163 9183 11169
rect 9309 11169 9321 11172
rect 9355 11169 9367 11203
rect 9309 11163 9367 11169
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 8482 11135 8540 11141
rect 8482 11101 8494 11135
rect 8528 11101 8540 11135
rect 8482 11095 8540 11101
rect 8665 11135 8723 11141
rect 8665 11101 8677 11135
rect 8711 11132 8723 11135
rect 8754 11132 8760 11144
rect 8711 11104 8760 11132
rect 8711 11101 8723 11104
rect 8665 11095 8723 11101
rect 6914 11064 6920 11076
rect 6052 11036 6097 11064
rect 6196 11036 6920 11064
rect 6052 11024 6058 11036
rect 4948 10968 5948 10996
rect 6549 10999 6607 11005
rect 4948 10956 4954 10968
rect 6549 10965 6561 10999
rect 6595 10996 6607 10999
rect 6638 10996 6644 11008
rect 6595 10968 6644 10996
rect 6595 10965 6607 10968
rect 6549 10959 6607 10965
rect 6638 10956 6644 10968
rect 6696 10956 6702 11008
rect 6748 11005 6776 11036
rect 6914 11024 6920 11036
rect 6972 11064 6978 11076
rect 7285 11067 7343 11073
rect 7285 11064 7297 11067
rect 6972 11036 7297 11064
rect 6972 11024 6978 11036
rect 7285 11033 7297 11036
rect 7331 11033 7343 11067
rect 8404 11064 8432 11095
rect 8754 11092 8760 11104
rect 8812 11092 8818 11144
rect 9140 11064 9168 11163
rect 9674 11160 9680 11212
rect 9732 11200 9738 11212
rect 11701 11203 11759 11209
rect 11701 11200 11713 11203
rect 9732 11172 11713 11200
rect 9732 11160 9738 11172
rect 11701 11169 11713 11172
rect 11747 11169 11759 11203
rect 11882 11200 11888 11212
rect 11843 11172 11888 11200
rect 11701 11163 11759 11169
rect 11882 11160 11888 11172
rect 11940 11160 11946 11212
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11132 9459 11135
rect 9766 11132 9772 11144
rect 9447 11104 9772 11132
rect 9447 11101 9459 11104
rect 9401 11095 9459 11101
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 9861 11135 9919 11141
rect 9861 11101 9873 11135
rect 9907 11101 9919 11135
rect 9861 11095 9919 11101
rect 11057 11135 11115 11141
rect 11057 11101 11069 11135
rect 11103 11101 11115 11135
rect 11057 11095 11115 11101
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11132 12587 11135
rect 12710 11132 12716 11144
rect 12575 11104 12716 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 9674 11064 9680 11076
rect 8404 11036 8616 11064
rect 9140 11036 9680 11064
rect 7285 11027 7343 11033
rect 8588 11008 8616 11036
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 6733 10999 6791 11005
rect 6733 10965 6745 10999
rect 6779 10965 6791 10999
rect 6733 10959 6791 10965
rect 7006 10956 7012 11008
rect 7064 10996 7070 11008
rect 7377 10999 7435 11005
rect 7377 10996 7389 10999
rect 7064 10968 7389 10996
rect 7064 10956 7070 10968
rect 7377 10965 7389 10968
rect 7423 10965 7435 10999
rect 7377 10959 7435 10965
rect 8570 10956 8576 11008
rect 8628 10956 8634 11008
rect 9769 10999 9827 11005
rect 9769 10965 9781 10999
rect 9815 10996 9827 10999
rect 9876 10996 9904 11095
rect 10594 10996 10600 11008
rect 9815 10968 10600 10996
rect 9815 10965 9827 10968
rect 9769 10959 9827 10965
rect 10594 10956 10600 10968
rect 10652 10956 10658 11008
rect 10686 10956 10692 11008
rect 10744 10996 10750 11008
rect 11072 10996 11100 11095
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 13446 11132 13452 11144
rect 13407 11104 13452 11132
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 12437 11067 12495 11073
rect 12437 11033 12449 11067
rect 12483 11064 12495 11067
rect 12802 11064 12808 11076
rect 12483 11036 12808 11064
rect 12483 11033 12495 11036
rect 12437 11027 12495 11033
rect 12802 11024 12808 11036
rect 12860 11024 12866 11076
rect 13170 11064 13176 11076
rect 13131 11036 13176 11064
rect 13170 11024 13176 11036
rect 13228 11024 13234 11076
rect 10744 10968 11100 10996
rect 10744 10956 10750 10968
rect 1104 10906 13892 10928
rect 1104 10854 8214 10906
rect 8266 10854 8278 10906
rect 8330 10854 8342 10906
rect 8394 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 13892 10906
rect 1104 10832 13892 10854
rect 2222 10792 2228 10804
rect 2183 10764 2228 10792
rect 2222 10752 2228 10764
rect 2280 10752 2286 10804
rect 2958 10752 2964 10804
rect 3016 10792 3022 10804
rect 3237 10795 3295 10801
rect 3237 10792 3249 10795
rect 3016 10764 3249 10792
rect 3016 10752 3022 10764
rect 3237 10761 3249 10764
rect 3283 10761 3295 10795
rect 4062 10792 4068 10804
rect 3237 10755 3295 10761
rect 3528 10764 3924 10792
rect 4023 10764 4068 10792
rect 2590 10724 2596 10736
rect 2551 10696 2596 10724
rect 2590 10684 2596 10696
rect 2648 10684 2654 10736
rect 3528 10733 3556 10764
rect 3513 10727 3571 10733
rect 3513 10693 3525 10727
rect 3559 10693 3571 10727
rect 3786 10724 3792 10736
rect 3513 10687 3571 10693
rect 3727 10696 3792 10724
rect 2038 10656 2044 10668
rect 1999 10628 2044 10656
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 2406 10656 2412 10668
rect 2367 10628 2412 10656
rect 2406 10616 2412 10628
rect 2464 10616 2470 10668
rect 2866 10665 2872 10668
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10625 2743 10659
rect 2685 10619 2743 10625
rect 2829 10659 2872 10665
rect 2829 10625 2841 10659
rect 2829 10619 2872 10625
rect 1486 10548 1492 10600
rect 1544 10588 1550 10600
rect 2700 10588 2728 10619
rect 2866 10616 2872 10619
rect 2924 10616 2930 10668
rect 3142 10616 3148 10668
rect 3200 10616 3206 10668
rect 3326 10616 3332 10668
rect 3384 10654 3390 10668
rect 3421 10659 3479 10665
rect 3421 10654 3433 10659
rect 3384 10626 3433 10654
rect 3384 10616 3390 10626
rect 3421 10625 3433 10626
rect 3467 10625 3479 10659
rect 3603 10656 3609 10668
rect 3661 10665 3667 10668
rect 3727 10665 3755 10696
rect 3786 10684 3792 10696
rect 3844 10684 3850 10736
rect 3896 10724 3924 10764
rect 4062 10752 4068 10764
rect 4120 10752 4126 10804
rect 4246 10752 4252 10804
rect 4304 10792 4310 10804
rect 4341 10795 4399 10801
rect 4341 10792 4353 10795
rect 4304 10764 4353 10792
rect 4304 10752 4310 10764
rect 4341 10761 4353 10764
rect 4387 10761 4399 10795
rect 4341 10755 4399 10761
rect 4433 10795 4491 10801
rect 4433 10761 4445 10795
rect 4479 10792 4491 10795
rect 4982 10792 4988 10804
rect 4479 10764 4988 10792
rect 4479 10761 4491 10764
rect 4433 10755 4491 10761
rect 3970 10724 3976 10736
rect 3896 10696 3976 10724
rect 3970 10684 3976 10696
rect 4028 10724 4034 10736
rect 4448 10724 4476 10755
rect 4982 10752 4988 10764
rect 5040 10752 5046 10804
rect 7834 10752 7840 10804
rect 7892 10792 7898 10804
rect 8754 10792 8760 10804
rect 7892 10764 8760 10792
rect 7892 10752 7898 10764
rect 8754 10752 8760 10764
rect 8812 10752 8818 10804
rect 9122 10752 9128 10804
rect 9180 10792 9186 10804
rect 10318 10792 10324 10804
rect 9180 10764 10324 10792
rect 9180 10752 9186 10764
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 4028 10696 4476 10724
rect 5445 10727 5503 10733
rect 4028 10684 4034 10696
rect 5445 10693 5457 10727
rect 5491 10724 5503 10727
rect 7101 10727 7159 10733
rect 5491 10696 7052 10724
rect 5491 10693 5503 10696
rect 5445 10687 5503 10693
rect 3568 10628 3609 10656
rect 3421 10619 3479 10625
rect 3603 10616 3609 10628
rect 3661 10619 3668 10665
rect 3697 10659 3755 10665
rect 3697 10625 3709 10659
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 3881 10659 3939 10665
rect 3881 10625 3893 10659
rect 3927 10625 3939 10659
rect 3881 10619 3939 10625
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10656 4307 10659
rect 4522 10656 4528 10668
rect 4295 10628 4528 10656
rect 4295 10625 4307 10628
rect 4249 10619 4307 10625
rect 3661 10616 3667 10619
rect 3050 10588 3056 10600
rect 1544 10560 3056 10588
rect 1544 10548 1550 10560
rect 3050 10548 3056 10560
rect 3108 10548 3114 10600
rect 3160 10588 3188 10616
rect 3727 10588 3755 10619
rect 3160 10560 3755 10588
rect 3786 10548 3792 10600
rect 3844 10588 3850 10600
rect 3896 10588 3924 10619
rect 4522 10616 4528 10628
rect 4580 10616 4586 10668
rect 4890 10656 4896 10668
rect 4851 10628 4896 10656
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10656 5135 10659
rect 5258 10656 5264 10668
rect 5123 10628 5264 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 5258 10616 5264 10628
rect 5316 10656 5322 10668
rect 5721 10659 5779 10665
rect 5721 10656 5733 10659
rect 5316 10628 5733 10656
rect 5316 10616 5322 10628
rect 5721 10625 5733 10628
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 5810 10616 5816 10668
rect 5868 10656 5874 10668
rect 6457 10659 6515 10665
rect 6457 10656 6469 10659
rect 5868 10628 6469 10656
rect 5868 10616 5874 10628
rect 6457 10625 6469 10628
rect 6503 10625 6515 10659
rect 6457 10619 6515 10625
rect 4338 10588 4344 10600
rect 3844 10560 4344 10588
rect 3844 10548 3850 10560
rect 4338 10548 4344 10560
rect 4396 10548 4402 10600
rect 4617 10591 4675 10597
rect 4617 10557 4629 10591
rect 4663 10588 4675 10591
rect 4709 10591 4767 10597
rect 4709 10588 4721 10591
rect 4663 10560 4721 10588
rect 4663 10557 4675 10560
rect 4617 10551 4675 10557
rect 4709 10557 4721 10560
rect 4755 10557 4767 10591
rect 4908 10588 4936 10616
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 4908 10560 5641 10588
rect 4709 10551 4767 10557
rect 5629 10557 5641 10560
rect 5675 10557 5687 10591
rect 6472 10588 6500 10619
rect 6546 10616 6552 10668
rect 6604 10656 6610 10668
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 6604 10628 6745 10656
rect 6604 10616 6610 10628
rect 6733 10625 6745 10628
rect 6779 10625 6791 10659
rect 6914 10656 6920 10668
rect 6875 10628 6920 10656
rect 6733 10619 6791 10625
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 7024 10656 7052 10696
rect 7101 10693 7113 10727
rect 7147 10724 7159 10727
rect 7190 10724 7196 10736
rect 7147 10696 7196 10724
rect 7147 10693 7159 10696
rect 7101 10687 7159 10693
rect 7190 10684 7196 10696
rect 7248 10684 7254 10736
rect 7745 10727 7803 10733
rect 7745 10693 7757 10727
rect 7791 10724 7803 10727
rect 10134 10724 10140 10736
rect 7791 10696 9720 10724
rect 10095 10696 10140 10724
rect 7791 10693 7803 10696
rect 7745 10687 7803 10693
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 7024 10628 7389 10656
rect 7377 10625 7389 10628
rect 7423 10656 7435 10659
rect 7466 10656 7472 10668
rect 7423 10628 7472 10656
rect 7423 10625 7435 10628
rect 7377 10619 7435 10625
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 7650 10656 7656 10668
rect 7611 10628 7656 10656
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 7834 10656 7840 10668
rect 7795 10628 7840 10656
rect 7834 10616 7840 10628
rect 7892 10616 7898 10668
rect 8018 10656 8024 10668
rect 7979 10628 8024 10656
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 8386 10656 8392 10668
rect 8347 10628 8392 10656
rect 8386 10616 8392 10628
rect 8444 10616 8450 10668
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10625 8539 10659
rect 8481 10619 8539 10625
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10656 8907 10659
rect 9030 10656 9036 10668
rect 8895 10628 9036 10656
rect 8895 10625 8907 10628
rect 8849 10619 8907 10625
rect 8496 10588 8524 10619
rect 9030 10616 9036 10628
rect 9088 10616 9094 10668
rect 9122 10616 9128 10668
rect 9180 10656 9186 10668
rect 9692 10665 9720 10696
rect 10134 10684 10140 10696
rect 10192 10684 10198 10736
rect 11054 10724 11060 10736
rect 11015 10696 11060 10724
rect 11054 10684 11060 10696
rect 11112 10684 11118 10736
rect 12434 10724 12440 10736
rect 12395 10696 12440 10724
rect 12434 10684 12440 10696
rect 12492 10684 12498 10736
rect 13170 10724 13176 10736
rect 13131 10696 13176 10724
rect 13170 10684 13176 10696
rect 13228 10684 13234 10736
rect 9511 10659 9569 10665
rect 9180 10628 9225 10656
rect 9180 10616 9186 10628
rect 9511 10625 9523 10659
rect 9557 10656 9569 10659
rect 9677 10659 9735 10665
rect 9557 10628 9628 10656
rect 9557 10625 9569 10628
rect 9511 10619 9569 10625
rect 6472 10560 8524 10588
rect 5629 10551 5687 10557
rect 9214 10548 9220 10600
rect 9272 10588 9278 10600
rect 9309 10591 9367 10597
rect 9309 10588 9321 10591
rect 9272 10560 9321 10588
rect 9272 10548 9278 10560
rect 9309 10557 9321 10560
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 9401 10591 9459 10597
rect 9401 10557 9413 10591
rect 9447 10557 9459 10591
rect 9600 10588 9628 10628
rect 9677 10625 9689 10659
rect 9723 10625 9735 10659
rect 9677 10619 9735 10625
rect 9766 10616 9772 10668
rect 9824 10656 9830 10668
rect 9824 10628 9869 10656
rect 9824 10616 9830 10628
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 10594 10656 10600 10668
rect 10008 10628 10053 10656
rect 10555 10628 10600 10656
rect 10008 10616 10014 10628
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 10686 10616 10692 10668
rect 10744 10656 10750 10668
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 10744 10628 11529 10656
rect 10744 10616 10750 10628
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 11606 10616 11612 10668
rect 11664 10656 11670 10668
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 11664 10628 11805 10656
rect 11664 10616 11670 10628
rect 11793 10625 11805 10628
rect 11839 10625 11851 10659
rect 11793 10619 11851 10625
rect 13446 10616 13452 10668
rect 13504 10656 13510 10668
rect 13541 10659 13599 10665
rect 13541 10656 13553 10659
rect 13504 10628 13553 10656
rect 13504 10616 13510 10628
rect 13541 10625 13553 10628
rect 13587 10625 13599 10659
rect 13541 10619 13599 10625
rect 11149 10591 11207 10597
rect 9600 10560 10548 10588
rect 9401 10551 9459 10557
rect 2314 10480 2320 10532
rect 2372 10520 2378 10532
rect 6549 10523 6607 10529
rect 2372 10492 6500 10520
rect 2372 10480 2378 10492
rect 2958 10452 2964 10464
rect 2919 10424 2964 10452
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 3602 10412 3608 10464
rect 3660 10452 3666 10464
rect 4709 10455 4767 10461
rect 4709 10452 4721 10455
rect 3660 10424 4721 10452
rect 3660 10412 3666 10424
rect 4709 10421 4721 10424
rect 4755 10452 4767 10455
rect 5166 10452 5172 10464
rect 4755 10424 5172 10452
rect 4755 10421 4767 10424
rect 4709 10415 4767 10421
rect 5166 10412 5172 10424
rect 5224 10452 5230 10464
rect 5534 10452 5540 10464
rect 5224 10424 5540 10452
rect 5224 10412 5230 10424
rect 5534 10412 5540 10424
rect 5592 10452 5598 10464
rect 6362 10452 6368 10464
rect 5592 10424 6368 10452
rect 5592 10412 5598 10424
rect 6362 10412 6368 10424
rect 6420 10412 6426 10464
rect 6472 10452 6500 10492
rect 6549 10489 6561 10523
rect 6595 10520 6607 10523
rect 9416 10520 9444 10551
rect 6595 10492 9444 10520
rect 6595 10489 6607 10492
rect 6549 10483 6607 10489
rect 10520 10464 10548 10560
rect 11149 10557 11161 10591
rect 11195 10588 11207 10591
rect 11885 10591 11943 10597
rect 11885 10588 11897 10591
rect 11195 10560 11897 10588
rect 11195 10557 11207 10560
rect 11149 10551 11207 10557
rect 11885 10557 11897 10560
rect 11931 10557 11943 10591
rect 12710 10588 12716 10600
rect 12671 10560 12716 10588
rect 11885 10551 11943 10557
rect 12710 10548 12716 10560
rect 12768 10548 12774 10600
rect 13265 10591 13323 10597
rect 13265 10557 13277 10591
rect 13311 10557 13323 10591
rect 13265 10551 13323 10557
rect 12618 10520 12624 10532
rect 12579 10492 12624 10520
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 13280 10520 13308 10551
rect 13357 10523 13415 10529
rect 13357 10520 13369 10523
rect 13280 10492 13369 10520
rect 13357 10489 13369 10492
rect 13403 10489 13415 10523
rect 13357 10483 13415 10489
rect 7006 10452 7012 10464
rect 6472 10424 7012 10452
rect 7006 10412 7012 10424
rect 7064 10412 7070 10464
rect 7926 10452 7932 10464
rect 7887 10424 7932 10452
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 8386 10412 8392 10464
rect 8444 10452 8450 10464
rect 9033 10455 9091 10461
rect 9033 10452 9045 10455
rect 8444 10424 9045 10452
rect 8444 10412 8450 10424
rect 9033 10421 9045 10424
rect 9079 10421 9091 10455
rect 10502 10452 10508 10464
rect 10463 10424 10508 10452
rect 9033 10415 9091 10421
rect 10502 10412 10508 10424
rect 10560 10412 10566 10464
rect 11701 10455 11759 10461
rect 11701 10421 11713 10455
rect 11747 10452 11759 10455
rect 11790 10452 11796 10464
rect 11747 10424 11796 10452
rect 11747 10421 11759 10424
rect 11701 10415 11759 10421
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 1104 10362 13892 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 12214 10362
rect 12266 10310 12278 10362
rect 12330 10310 12342 10362
rect 12394 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 13892 10362
rect 1104 10288 13892 10310
rect 1486 10248 1492 10260
rect 1447 10220 1492 10248
rect 1486 10208 1492 10220
rect 1544 10208 1550 10260
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 6914 10248 6920 10260
rect 2832 10220 6776 10248
rect 6875 10220 6920 10248
rect 2832 10208 2838 10220
rect 3878 10140 3884 10192
rect 3936 10140 3942 10192
rect 4062 10180 4068 10192
rect 4023 10152 4068 10180
rect 4062 10140 4068 10152
rect 4120 10140 4126 10192
rect 4614 10180 4620 10192
rect 4264 10152 4620 10180
rect 2958 10112 2964 10124
rect 2919 10084 2964 10112
rect 2958 10072 2964 10084
rect 3016 10072 3022 10124
rect 3237 10115 3295 10121
rect 3237 10081 3249 10115
rect 3283 10112 3295 10115
rect 3418 10112 3424 10124
rect 3283 10084 3424 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 3896 10112 3924 10140
rect 4264 10121 4292 10152
rect 4614 10140 4620 10152
rect 4672 10140 4678 10192
rect 6748 10180 6776 10220
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 7650 10248 7656 10260
rect 7392 10220 7656 10248
rect 7392 10180 7420 10220
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 7800 10220 7941 10248
rect 7800 10208 7806 10220
rect 7929 10217 7941 10220
rect 7975 10248 7987 10251
rect 8202 10248 8208 10260
rect 7975 10220 8208 10248
rect 7975 10217 7987 10220
rect 7929 10211 7987 10217
rect 8202 10208 8208 10220
rect 8260 10248 8266 10260
rect 8757 10251 8815 10257
rect 8757 10248 8769 10251
rect 8260 10220 8769 10248
rect 8260 10208 8266 10220
rect 8757 10217 8769 10220
rect 8803 10248 8815 10251
rect 8938 10248 8944 10260
rect 8803 10220 8944 10248
rect 8803 10217 8815 10220
rect 8757 10211 8815 10217
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 9030 10208 9036 10260
rect 9088 10248 9094 10260
rect 9493 10251 9551 10257
rect 9493 10248 9505 10251
rect 9088 10220 9505 10248
rect 9088 10208 9094 10220
rect 9493 10217 9505 10220
rect 9539 10217 9551 10251
rect 9493 10211 9551 10217
rect 9769 10251 9827 10257
rect 9769 10217 9781 10251
rect 9815 10248 9827 10251
rect 10502 10248 10508 10260
rect 9815 10220 10508 10248
rect 9815 10217 9827 10220
rect 9769 10211 9827 10217
rect 6748 10152 7420 10180
rect 7466 10140 7472 10192
rect 7524 10180 7530 10192
rect 8481 10183 8539 10189
rect 7524 10152 8432 10180
rect 7524 10140 7530 10152
rect 4249 10115 4307 10121
rect 3896 10084 4200 10112
rect 3602 10004 3608 10056
rect 3660 10044 3666 10056
rect 3881 10047 3939 10053
rect 3881 10044 3893 10047
rect 3660 10016 3893 10044
rect 3660 10004 3666 10016
rect 3881 10013 3893 10016
rect 3927 10013 3939 10047
rect 3881 10007 3939 10013
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 4028 10016 4077 10044
rect 4028 10004 4034 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4172 10044 4200 10084
rect 4249 10081 4261 10115
rect 4295 10081 4307 10115
rect 4249 10075 4307 10081
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10112 4859 10115
rect 4890 10112 4896 10124
rect 4847 10084 4896 10112
rect 4847 10081 4859 10084
rect 4801 10075 4859 10081
rect 4890 10072 4896 10084
rect 4948 10072 4954 10124
rect 5442 10112 5448 10124
rect 5403 10084 5448 10112
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 6638 10072 6644 10124
rect 6696 10112 6702 10124
rect 7101 10115 7159 10121
rect 7101 10112 7113 10115
rect 6696 10084 7113 10112
rect 6696 10072 6702 10084
rect 7101 10081 7113 10084
rect 7147 10081 7159 10115
rect 7101 10075 7159 10081
rect 7193 10115 7251 10121
rect 7193 10081 7205 10115
rect 7239 10112 7251 10115
rect 7374 10112 7380 10124
rect 7239 10084 7380 10112
rect 7239 10081 7251 10084
rect 7193 10075 7251 10081
rect 7374 10072 7380 10084
rect 7432 10072 7438 10124
rect 8036 10121 8064 10152
rect 8021 10115 8079 10121
rect 8021 10081 8033 10115
rect 8067 10081 8079 10115
rect 8404 10112 8432 10152
rect 8481 10149 8493 10183
rect 8527 10180 8539 10183
rect 8570 10180 8576 10192
rect 8527 10152 8576 10180
rect 8527 10149 8539 10152
rect 8481 10143 8539 10149
rect 8570 10140 8576 10152
rect 8628 10140 8634 10192
rect 9214 10180 9220 10192
rect 8680 10152 9220 10180
rect 8680 10112 8708 10152
rect 9214 10140 9220 10152
rect 9272 10140 9278 10192
rect 8404 10084 8708 10112
rect 8021 10075 8079 10081
rect 8754 10072 8760 10124
rect 8812 10112 8818 10124
rect 9309 10115 9367 10121
rect 9309 10112 9321 10115
rect 8812 10084 9321 10112
rect 8812 10072 8818 10084
rect 9309 10081 9321 10084
rect 9355 10081 9367 10115
rect 9309 10075 9367 10081
rect 4433 10047 4491 10053
rect 4433 10044 4445 10047
rect 4172 10016 4445 10044
rect 4065 10007 4123 10013
rect 4433 10013 4445 10016
rect 4479 10013 4491 10047
rect 5166 10044 5172 10056
rect 5127 10016 5172 10044
rect 4433 10007 4491 10013
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 7282 10004 7288 10056
rect 7340 10044 7346 10056
rect 7503 10047 7561 10053
rect 7503 10044 7515 10047
rect 7340 10016 7515 10044
rect 7340 10004 7346 10016
rect 7503 10013 7515 10016
rect 7549 10013 7561 10047
rect 8202 10044 8208 10056
rect 8163 10016 8208 10044
rect 7503 10007 7561 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 8386 10004 8392 10056
rect 8444 10044 8450 10056
rect 8573 10047 8631 10053
rect 8573 10044 8585 10047
rect 8444 10016 8585 10044
rect 8444 10004 8450 10016
rect 8573 10013 8585 10016
rect 8619 10013 8631 10047
rect 8573 10007 8631 10013
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 9585 10047 9643 10053
rect 9585 10013 9597 10047
rect 9631 10044 9643 10047
rect 9784 10044 9812 10211
rect 10502 10208 10508 10220
rect 10560 10208 10566 10260
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 13173 10251 13231 10257
rect 13173 10248 13185 10251
rect 12860 10220 13185 10248
rect 12860 10208 12866 10220
rect 13173 10217 13185 10220
rect 13219 10217 13231 10251
rect 13173 10211 13231 10217
rect 9953 10183 10011 10189
rect 9953 10149 9965 10183
rect 9999 10180 10011 10183
rect 10042 10180 10048 10192
rect 9999 10152 10048 10180
rect 9999 10149 10011 10152
rect 9953 10143 10011 10149
rect 9631 10016 9812 10044
rect 9631 10013 9643 10016
rect 9585 10007 9643 10013
rect 2222 9936 2228 9988
rect 2280 9936 2286 9988
rect 4709 9979 4767 9985
rect 4709 9945 4721 9979
rect 4755 9976 4767 9979
rect 5718 9976 5724 9988
rect 4755 9948 5724 9976
rect 4755 9945 4767 9948
rect 4709 9939 4767 9945
rect 5718 9936 5724 9948
rect 5776 9936 5782 9988
rect 5902 9936 5908 9988
rect 5960 9936 5966 9988
rect 7006 9936 7012 9988
rect 7064 9976 7070 9988
rect 7745 9979 7803 9985
rect 7745 9976 7757 9979
rect 7064 9948 7757 9976
rect 7064 9936 7070 9948
rect 7745 9945 7757 9948
rect 7791 9976 7803 9979
rect 8956 9976 8984 10007
rect 7791 9948 8984 9976
rect 9232 9976 9260 10007
rect 9968 9976 9996 10143
rect 10042 10140 10048 10152
rect 10100 10140 10106 10192
rect 11790 10112 11796 10124
rect 11751 10084 11796 10112
rect 11790 10072 11796 10084
rect 11848 10072 11854 10124
rect 11698 10044 11704 10056
rect 11659 10016 11704 10044
rect 11698 10004 11704 10016
rect 11756 10044 11762 10056
rect 12345 10047 12403 10053
rect 12345 10044 12357 10047
rect 11756 10016 12357 10044
rect 11756 10004 11762 10016
rect 12345 10013 12357 10016
rect 12391 10013 12403 10047
rect 12345 10007 12403 10013
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 12492 10016 12537 10044
rect 12492 10004 12498 10016
rect 13170 10004 13176 10056
rect 13228 10044 13234 10056
rect 13265 10047 13323 10053
rect 13265 10044 13277 10047
rect 13228 10016 13277 10044
rect 13228 10004 13234 10016
rect 13265 10013 13277 10016
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 9232 9948 9996 9976
rect 7791 9945 7803 9948
rect 7745 9939 7803 9945
rect 3510 9868 3516 9920
rect 3568 9908 3574 9920
rect 7190 9908 7196 9920
rect 3568 9880 7196 9908
rect 3568 9868 3574 9880
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 7466 9868 7472 9920
rect 7524 9908 7530 9920
rect 9232 9908 9260 9948
rect 10686 9936 10692 9988
rect 10744 9976 10750 9988
rect 10781 9979 10839 9985
rect 10781 9976 10793 9979
rect 10744 9948 10793 9976
rect 10744 9936 10750 9948
rect 10781 9945 10793 9948
rect 10827 9945 10839 9979
rect 10781 9939 10839 9945
rect 11057 9979 11115 9985
rect 11057 9945 11069 9979
rect 11103 9976 11115 9979
rect 11606 9976 11612 9988
rect 11103 9948 11612 9976
rect 11103 9945 11115 9948
rect 11057 9939 11115 9945
rect 11606 9936 11612 9948
rect 11664 9976 11670 9988
rect 11885 9979 11943 9985
rect 11885 9976 11897 9979
rect 11664 9948 11897 9976
rect 11664 9936 11670 9948
rect 11885 9945 11897 9948
rect 11931 9945 11943 9979
rect 12894 9976 12900 9988
rect 12855 9948 12900 9976
rect 11885 9939 11943 9945
rect 12894 9936 12900 9948
rect 12952 9936 12958 9988
rect 12989 9979 13047 9985
rect 12989 9945 13001 9979
rect 13035 9976 13047 9979
rect 13449 9979 13507 9985
rect 13449 9976 13461 9979
rect 13035 9948 13461 9976
rect 13035 9945 13047 9948
rect 12989 9939 13047 9945
rect 13449 9945 13461 9948
rect 13495 9945 13507 9979
rect 13449 9939 13507 9945
rect 7524 9880 9260 9908
rect 7524 9868 7530 9880
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 10045 9911 10103 9917
rect 10045 9908 10057 9911
rect 9732 9880 10057 9908
rect 9732 9868 9738 9880
rect 10045 9877 10057 9880
rect 10091 9877 10103 9911
rect 13354 9908 13360 9920
rect 13315 9880 13360 9908
rect 10045 9871 10103 9877
rect 13354 9868 13360 9880
rect 13412 9868 13418 9920
rect 1104 9818 13892 9840
rect 1104 9766 8214 9818
rect 8266 9766 8278 9818
rect 8330 9766 8342 9818
rect 8394 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 13892 9818
rect 1104 9744 13892 9766
rect 2133 9707 2191 9713
rect 2133 9673 2145 9707
rect 2179 9704 2191 9707
rect 2222 9704 2228 9716
rect 2179 9676 2228 9704
rect 2179 9673 2191 9676
rect 2133 9667 2191 9673
rect 2222 9664 2228 9676
rect 2280 9664 2286 9716
rect 3970 9704 3976 9716
rect 3344 9676 3976 9704
rect 2866 9596 2872 9648
rect 2924 9636 2930 9648
rect 3234 9636 3240 9648
rect 2924 9608 3240 9636
rect 2924 9596 2930 9608
rect 2038 9528 2044 9580
rect 2096 9568 2102 9580
rect 2976 9577 3004 9608
rect 3234 9596 3240 9608
rect 3292 9596 3298 9648
rect 2317 9571 2375 9577
rect 2317 9568 2329 9571
rect 2096 9540 2329 9568
rect 2096 9528 2102 9540
rect 2317 9537 2329 9540
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9537 3019 9571
rect 3142 9568 3148 9580
rect 3103 9540 3148 9568
rect 2961 9531 3019 9537
rect 3142 9528 3148 9540
rect 3200 9528 3206 9580
rect 3344 9577 3372 9676
rect 3970 9664 3976 9676
rect 4028 9664 4034 9716
rect 5534 9704 5540 9716
rect 5495 9676 5540 9704
rect 5534 9664 5540 9676
rect 5592 9664 5598 9716
rect 7190 9664 7196 9716
rect 7248 9704 7254 9716
rect 14001 9707 14059 9713
rect 7248 9676 7420 9704
rect 7248 9664 7254 9676
rect 3697 9639 3755 9645
rect 3697 9605 3709 9639
rect 3743 9636 3755 9639
rect 4065 9639 4123 9645
rect 4065 9636 4077 9639
rect 3743 9608 4077 9636
rect 3743 9605 3755 9608
rect 3697 9599 3755 9605
rect 4065 9605 4077 9608
rect 4111 9605 4123 9639
rect 4065 9599 4123 9605
rect 4798 9596 4804 9648
rect 4856 9596 4862 9648
rect 6181 9639 6239 9645
rect 6181 9605 6193 9639
rect 6227 9636 6239 9639
rect 6638 9636 6644 9648
rect 6227 9608 6644 9636
rect 6227 9605 6239 9608
rect 6181 9599 6239 9605
rect 6638 9596 6644 9608
rect 6696 9596 6702 9648
rect 7282 9636 7288 9648
rect 6748 9608 7288 9636
rect 3329 9571 3387 9577
rect 3329 9537 3341 9571
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 3513 9571 3571 9577
rect 3513 9537 3525 9571
rect 3559 9568 3571 9571
rect 3602 9568 3608 9580
rect 3559 9540 3608 9568
rect 3559 9537 3571 9540
rect 3513 9531 3571 9537
rect 3602 9528 3608 9540
rect 3660 9528 3666 9580
rect 5994 9568 6000 9580
rect 5955 9540 6000 9568
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9568 6423 9571
rect 6748 9568 6776 9608
rect 7282 9596 7288 9608
rect 7340 9596 7346 9648
rect 7392 9636 7420 9676
rect 14001 9673 14013 9707
rect 14047 9704 14059 9707
rect 14182 9704 14188 9716
rect 14047 9676 14188 9704
rect 14047 9673 14059 9676
rect 14001 9667 14059 9673
rect 14182 9664 14188 9676
rect 14240 9664 14246 9716
rect 8386 9636 8392 9648
rect 7392 9608 8392 9636
rect 8386 9596 8392 9608
rect 8444 9636 8450 9648
rect 8573 9639 8631 9645
rect 8573 9636 8585 9639
rect 8444 9608 8585 9636
rect 8444 9596 8450 9608
rect 8573 9605 8585 9608
rect 8619 9605 8631 9639
rect 8573 9599 8631 9605
rect 11241 9639 11299 9645
rect 11241 9605 11253 9639
rect 11287 9636 11299 9639
rect 13354 9636 13360 9648
rect 11287 9608 13360 9636
rect 11287 9605 11299 9608
rect 11241 9599 11299 9605
rect 13354 9596 13360 9608
rect 13412 9596 13418 9648
rect 6411 9540 6776 9568
rect 6825 9571 6883 9577
rect 6411 9537 6423 9540
rect 6365 9531 6423 9537
rect 6825 9537 6837 9571
rect 6871 9568 6883 9571
rect 7006 9568 7012 9580
rect 6871 9540 7012 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 3237 9503 3295 9509
rect 3237 9469 3249 9503
rect 3283 9469 3295 9503
rect 3237 9463 3295 9469
rect 3252 9364 3280 9463
rect 3418 9460 3424 9512
rect 3476 9500 3482 9512
rect 3789 9503 3847 9509
rect 3789 9500 3801 9503
rect 3476 9472 3801 9500
rect 3476 9460 3482 9472
rect 3789 9469 3801 9472
rect 3835 9500 3847 9503
rect 5350 9500 5356 9512
rect 3835 9472 5356 9500
rect 3835 9469 3847 9472
rect 3789 9463 3847 9469
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 5813 9503 5871 9509
rect 5813 9469 5825 9503
rect 5859 9500 5871 9503
rect 6380 9500 6408 9531
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 7190 9568 7196 9580
rect 7151 9540 7196 9568
rect 7190 9528 7196 9540
rect 7248 9568 7254 9580
rect 7469 9571 7527 9577
rect 7469 9568 7481 9571
rect 7248 9540 7481 9568
rect 7248 9528 7254 9540
rect 7469 9537 7481 9540
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 7653 9571 7711 9577
rect 7653 9537 7665 9571
rect 7699 9537 7711 9571
rect 7653 9531 7711 9537
rect 6546 9500 6552 9512
rect 5859 9472 6408 9500
rect 6507 9472 6552 9500
rect 5859 9469 5871 9472
rect 5813 9463 5871 9469
rect 6546 9460 6552 9472
rect 6604 9460 6610 9512
rect 6638 9460 6644 9512
rect 6696 9500 6702 9512
rect 7101 9503 7159 9509
rect 7101 9500 7113 9503
rect 6696 9472 7113 9500
rect 6696 9460 6702 9472
rect 7101 9469 7113 9472
rect 7147 9500 7159 9503
rect 7668 9500 7696 9531
rect 7742 9528 7748 9580
rect 7800 9568 7806 9580
rect 7889 9571 7947 9577
rect 7800 9540 7845 9568
rect 7800 9528 7806 9540
rect 7889 9537 7901 9571
rect 7935 9568 7972 9571
rect 8018 9568 8024 9580
rect 7935 9540 8024 9568
rect 7935 9537 7947 9540
rect 7889 9531 7947 9537
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 8665 9571 8723 9577
rect 8665 9537 8677 9571
rect 8711 9568 8723 9571
rect 8938 9568 8944 9580
rect 8711 9540 8944 9568
rect 8711 9537 8723 9540
rect 8665 9531 8723 9537
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 9125 9571 9183 9577
rect 9125 9568 9137 9571
rect 9048 9540 9137 9568
rect 8478 9500 8484 9512
rect 7147 9472 7696 9500
rect 8439 9472 8484 9500
rect 7147 9469 7159 9472
rect 7101 9463 7159 9469
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 5994 9392 6000 9444
rect 6052 9432 6058 9444
rect 7374 9432 7380 9444
rect 6052 9404 7380 9432
rect 6052 9392 6058 9404
rect 7374 9392 7380 9404
rect 7432 9432 7438 9444
rect 8021 9435 8079 9441
rect 8021 9432 8033 9435
rect 7432 9404 8033 9432
rect 7432 9392 7438 9404
rect 8021 9401 8033 9404
rect 8067 9401 8079 9435
rect 8021 9395 8079 9401
rect 9048 9376 9076 9540
rect 9125 9537 9137 9540
rect 9171 9537 9183 9571
rect 10042 9568 10048 9580
rect 10003 9540 10048 9568
rect 9125 9531 9183 9537
rect 10042 9528 10048 9540
rect 10100 9528 10106 9580
rect 11514 9528 11520 9580
rect 11572 9568 11578 9580
rect 11609 9571 11667 9577
rect 11609 9568 11621 9571
rect 11572 9540 11621 9568
rect 11572 9528 11578 9540
rect 11609 9537 11621 9540
rect 11655 9568 11667 9571
rect 12434 9568 12440 9580
rect 11655 9540 12440 9568
rect 11655 9537 11667 9540
rect 11609 9531 11667 9537
rect 12434 9528 12440 9540
rect 12492 9528 12498 9580
rect 12618 9568 12624 9580
rect 12579 9540 12624 9568
rect 12618 9528 12624 9540
rect 12676 9568 12682 9580
rect 13078 9568 13084 9580
rect 12676 9540 13084 9568
rect 12676 9528 12682 9540
rect 13078 9528 13084 9540
rect 13136 9568 13142 9580
rect 13449 9571 13507 9577
rect 13449 9568 13461 9571
rect 13136 9540 13461 9568
rect 13136 9528 13142 9540
rect 13449 9537 13461 9540
rect 13495 9537 13507 9571
rect 13449 9531 13507 9537
rect 10594 9460 10600 9512
rect 10652 9500 10658 9512
rect 10781 9503 10839 9509
rect 10781 9500 10793 9503
rect 10652 9472 10793 9500
rect 10652 9460 10658 9472
rect 10781 9469 10793 9472
rect 10827 9469 10839 9503
rect 10781 9463 10839 9469
rect 11333 9503 11391 9509
rect 11333 9469 11345 9503
rect 11379 9500 11391 9503
rect 11379 9472 13308 9500
rect 11379 9469 11391 9472
rect 11333 9463 11391 9469
rect 10413 9435 10471 9441
rect 10413 9401 10425 9435
rect 10459 9432 10471 9435
rect 10502 9432 10508 9444
rect 10459 9404 10508 9432
rect 10459 9401 10471 9404
rect 10413 9395 10471 9401
rect 10502 9392 10508 9404
rect 10560 9392 10566 9444
rect 12894 9432 12900 9444
rect 12855 9404 12900 9432
rect 12894 9392 12900 9404
rect 12952 9392 12958 9444
rect 13280 9441 13308 9472
rect 13265 9435 13323 9441
rect 13265 9401 13277 9435
rect 13311 9401 13323 9435
rect 13265 9395 13323 9401
rect 4062 9364 4068 9376
rect 3252 9336 4068 9364
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 6454 9364 6460 9376
rect 6415 9336 6460 9364
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 6546 9324 6552 9376
rect 6604 9364 6610 9376
rect 7466 9364 7472 9376
rect 6604 9336 7472 9364
rect 6604 9324 6610 9336
rect 7466 9324 7472 9336
rect 7524 9324 7530 9376
rect 9030 9364 9036 9376
rect 8991 9336 9036 9364
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 1104 9274 13892 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 12214 9274
rect 12266 9222 12278 9274
rect 12330 9222 12342 9274
rect 12394 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 13892 9274
rect 1104 9200 13892 9222
rect 4798 9120 4804 9172
rect 4856 9160 4862 9172
rect 4893 9163 4951 9169
rect 4893 9160 4905 9163
rect 4856 9132 4905 9160
rect 4856 9120 4862 9132
rect 4893 9129 4905 9132
rect 4939 9129 4951 9163
rect 6638 9160 6644 9172
rect 4893 9123 4951 9129
rect 5092 9132 6644 9160
rect 3142 9092 3148 9104
rect 3055 9064 3148 9092
rect 3142 9052 3148 9064
rect 3200 9092 3206 9104
rect 4525 9095 4583 9101
rect 3200 9064 4476 9092
rect 3200 9052 3206 9064
rect 1673 9027 1731 9033
rect 1673 8993 1685 9027
rect 1719 9024 1731 9027
rect 3881 9027 3939 9033
rect 3881 9024 3893 9027
rect 1719 8996 3893 9024
rect 1719 8993 1731 8996
rect 1673 8987 1731 8993
rect 3881 8993 3893 8996
rect 3927 8993 3939 9027
rect 3881 8987 3939 8993
rect 4062 8984 4068 9036
rect 4120 9024 4126 9036
rect 4341 9027 4399 9033
rect 4341 9024 4353 9027
rect 4120 8996 4353 9024
rect 4120 8984 4126 8996
rect 4341 8993 4353 8996
rect 4387 8993 4399 9027
rect 4341 8987 4399 8993
rect 4448 8968 4476 9064
rect 4525 9061 4537 9095
rect 4571 9092 4583 9095
rect 5092 9092 5120 9132
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 7009 9163 7067 9169
rect 7009 9129 7021 9163
rect 7055 9160 7067 9163
rect 7190 9160 7196 9172
rect 7055 9132 7196 9160
rect 7055 9129 7067 9132
rect 7009 9123 7067 9129
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 7466 9160 7472 9172
rect 7427 9132 7472 9160
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 8386 9160 8392 9172
rect 8347 9132 8392 9160
rect 8386 9120 8392 9132
rect 8444 9120 8450 9172
rect 8478 9120 8484 9172
rect 8536 9160 8542 9172
rect 8665 9163 8723 9169
rect 8665 9160 8677 9163
rect 8536 9132 8677 9160
rect 8536 9120 8542 9132
rect 8665 9129 8677 9132
rect 8711 9160 8723 9163
rect 9217 9163 9275 9169
rect 9217 9160 9229 9163
rect 8711 9132 9229 9160
rect 8711 9129 8723 9132
rect 8665 9123 8723 9129
rect 9217 9129 9229 9132
rect 9263 9160 9275 9163
rect 9674 9160 9680 9172
rect 9263 9132 9680 9160
rect 9263 9129 9275 9132
rect 9217 9123 9275 9129
rect 9674 9120 9680 9132
rect 9732 9160 9738 9172
rect 11514 9160 11520 9172
rect 9732 9132 10824 9160
rect 11475 9132 11520 9160
rect 9732 9120 9738 9132
rect 4571 9064 5120 9092
rect 4571 9061 4583 9064
rect 4525 9055 4583 9061
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 3786 8956 3792 8968
rect 3747 8928 3792 8956
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8925 4215 8959
rect 4430 8956 4436 8968
rect 4391 8928 4436 8956
rect 4157 8919 4215 8925
rect 2406 8848 2412 8900
rect 2464 8848 2470 8900
rect 4172 8888 4200 8919
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 4540 8888 4568 9055
rect 6914 9052 6920 9104
rect 6972 9092 6978 9104
rect 7285 9095 7343 9101
rect 7285 9092 7297 9095
rect 6972 9064 7297 9092
rect 6972 9052 6978 9064
rect 7285 9061 7297 9064
rect 7331 9092 7343 9095
rect 7331 9064 8064 9092
rect 7331 9061 7343 9064
rect 7285 9055 7343 9061
rect 4985 9027 5043 9033
rect 4985 8993 4997 9027
rect 5031 9024 5043 9027
rect 5350 9024 5356 9036
rect 5031 8996 5356 9024
rect 5031 8993 5043 8996
rect 4985 8987 5043 8993
rect 5350 8984 5356 8996
rect 5408 8984 5414 9036
rect 8036 9033 8064 9064
rect 8021 9027 8079 9033
rect 8021 8993 8033 9027
rect 8067 8993 8079 9027
rect 8021 8987 8079 8993
rect 8205 9027 8263 9033
rect 8205 8993 8217 9027
rect 8251 9024 8263 9027
rect 8496 9024 8524 9120
rect 10686 9092 10692 9104
rect 10647 9064 10692 9092
rect 10686 9052 10692 9064
rect 10744 9052 10750 9104
rect 10796 9092 10824 9132
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 11609 9095 11667 9101
rect 11609 9092 11621 9095
rect 10796 9064 11621 9092
rect 8251 8996 8524 9024
rect 8251 8993 8263 8996
rect 8205 8987 8263 8993
rect 9030 8984 9036 9036
rect 9088 9024 9094 9036
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 9088 8996 9689 9024
rect 9088 8984 9094 8996
rect 9677 8993 9689 8996
rect 9723 8993 9735 9027
rect 9677 8987 9735 8993
rect 10137 9027 10195 9033
rect 10137 8993 10149 9027
rect 10183 9024 10195 9027
rect 10796 9024 10824 9064
rect 11609 9061 11621 9064
rect 11655 9092 11667 9095
rect 12618 9092 12624 9104
rect 11655 9064 12624 9092
rect 11655 9061 11667 9064
rect 11609 9055 11667 9061
rect 12618 9052 12624 9064
rect 12676 9052 12682 9104
rect 13354 9092 13360 9104
rect 12820 9064 13360 9092
rect 10870 9024 10876 9036
rect 10183 8996 10548 9024
rect 10783 8996 10876 9024
rect 10183 8993 10195 8996
rect 10137 8987 10195 8993
rect 10520 8968 10548 8996
rect 10870 8984 10876 8996
rect 10928 8984 10934 9036
rect 11057 9027 11115 9033
rect 11057 8993 11069 9027
rect 11103 9024 11115 9027
rect 11238 9024 11244 9036
rect 11103 8996 11244 9024
rect 11103 8993 11115 8996
rect 11057 8987 11115 8993
rect 11238 8984 11244 8996
rect 11296 9024 11302 9036
rect 11793 9027 11851 9033
rect 11793 9024 11805 9027
rect 11296 8996 11805 9024
rect 11296 8984 11302 8996
rect 11793 8993 11805 8996
rect 11839 8993 11851 9027
rect 11793 8987 11851 8993
rect 4614 8916 4620 8968
rect 4672 8956 4678 8968
rect 4709 8959 4767 8965
rect 4709 8956 4721 8959
rect 4672 8928 4721 8956
rect 4672 8916 4678 8928
rect 4709 8925 4721 8928
rect 4755 8925 4767 8959
rect 6917 8959 6975 8965
rect 6917 8956 6929 8959
rect 4709 8919 4767 8925
rect 6748 8928 6929 8956
rect 5258 8888 5264 8900
rect 4172 8860 4568 8888
rect 5219 8860 5264 8888
rect 5258 8848 5264 8860
rect 5316 8848 5322 8900
rect 5994 8848 6000 8900
rect 6052 8848 6058 8900
rect 6748 8888 6776 8928
rect 6917 8925 6929 8928
rect 6963 8925 6975 8959
rect 6917 8919 6975 8925
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8956 7987 8959
rect 8570 8956 8576 8968
rect 7975 8928 8576 8956
rect 7975 8925 7987 8928
rect 7929 8919 7987 8925
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 9493 8959 9551 8965
rect 9493 8925 9505 8959
rect 9539 8956 9551 8959
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 9539 8928 10241 8956
rect 9539 8925 9551 8928
rect 9493 8919 9551 8925
rect 10229 8925 10241 8928
rect 10275 8925 10287 8959
rect 10502 8956 10508 8968
rect 10463 8928 10508 8956
rect 10229 8919 10287 8925
rect 10502 8916 10508 8928
rect 10560 8916 10566 8968
rect 10594 8916 10600 8968
rect 10652 8956 10658 8968
rect 12820 8965 12848 9064
rect 13354 9052 13360 9064
rect 13412 9052 13418 9104
rect 12161 8959 12219 8965
rect 12161 8956 12173 8959
rect 10652 8928 12173 8956
rect 10652 8916 10658 8928
rect 12161 8925 12173 8928
rect 12207 8925 12219 8959
rect 12161 8919 12219 8925
rect 12805 8959 12863 8965
rect 12805 8925 12817 8959
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 12894 8916 12900 8968
rect 12952 8956 12958 8968
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 12952 8928 13369 8956
rect 12952 8916 12958 8928
rect 13357 8925 13369 8928
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 8018 8888 8024 8900
rect 6748 8860 8024 8888
rect 6748 8832 6776 8860
rect 8018 8848 8024 8860
rect 8076 8848 8082 8900
rect 13078 8888 13084 8900
rect 13039 8860 13084 8888
rect 13078 8848 13084 8860
rect 13136 8848 13142 8900
rect 13170 8848 13176 8900
rect 13228 8888 13234 8900
rect 13228 8860 13273 8888
rect 13228 8848 13234 8860
rect 3786 8780 3792 8832
rect 3844 8820 3850 8832
rect 4890 8820 4896 8832
rect 3844 8792 4896 8820
rect 3844 8780 3850 8792
rect 4890 8780 4896 8792
rect 4948 8780 4954 8832
rect 6730 8820 6736 8832
rect 6691 8792 6736 8820
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 7466 8780 7472 8832
rect 7524 8820 7530 8832
rect 7561 8823 7619 8829
rect 7561 8820 7573 8823
rect 7524 8792 7573 8820
rect 7524 8780 7530 8792
rect 7561 8789 7573 8792
rect 7607 8789 7619 8823
rect 9582 8820 9588 8832
rect 9543 8792 9588 8820
rect 7561 8783 7619 8789
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 11146 8780 11152 8832
rect 11204 8820 11210 8832
rect 11204 8792 11249 8820
rect 11204 8780 11210 8792
rect 1104 8730 13892 8752
rect 1104 8678 8214 8730
rect 8266 8678 8278 8730
rect 8330 8678 8342 8730
rect 8394 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 13892 8730
rect 1104 8656 13892 8678
rect 2406 8576 2412 8628
rect 2464 8616 2470 8628
rect 2501 8619 2559 8625
rect 2501 8616 2513 8619
rect 2464 8588 2513 8616
rect 2464 8576 2470 8588
rect 2501 8585 2513 8588
rect 2547 8585 2559 8619
rect 2501 8579 2559 8585
rect 3786 8576 3792 8628
rect 3844 8616 3850 8628
rect 4249 8619 4307 8625
rect 4249 8616 4261 8619
rect 3844 8588 4261 8616
rect 3844 8576 3850 8588
rect 4249 8585 4261 8588
rect 4295 8585 4307 8619
rect 4249 8579 4307 8585
rect 4614 8576 4620 8628
rect 4672 8616 4678 8628
rect 5902 8616 5908 8628
rect 4672 8588 5908 8616
rect 4672 8576 4678 8588
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 6089 8619 6147 8625
rect 6089 8616 6101 8619
rect 6052 8588 6101 8616
rect 6052 8576 6058 8588
rect 6089 8585 6101 8588
rect 6135 8585 6147 8619
rect 10042 8616 10048 8628
rect 6089 8579 6147 8585
rect 9508 8588 10048 8616
rect 3418 8548 3424 8560
rect 3331 8520 3424 8548
rect 3418 8508 3424 8520
rect 3476 8548 3482 8560
rect 3881 8551 3939 8557
rect 3881 8548 3893 8551
rect 3476 8520 3893 8548
rect 3476 8508 3482 8520
rect 3881 8517 3893 8520
rect 3927 8517 3939 8551
rect 3881 8511 3939 8517
rect 4157 8551 4215 8557
rect 4157 8517 4169 8551
rect 4203 8548 4215 8551
rect 4706 8548 4712 8560
rect 4203 8520 4712 8548
rect 4203 8517 4215 8520
rect 4157 8511 4215 8517
rect 2038 8480 2044 8492
rect 1999 8452 2044 8480
rect 2038 8440 2044 8452
rect 2096 8480 2102 8492
rect 2317 8483 2375 8489
rect 2317 8480 2329 8483
rect 2096 8452 2329 8480
rect 2096 8440 2102 8452
rect 2317 8449 2329 8452
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8480 3203 8483
rect 3234 8480 3240 8492
rect 3191 8452 3240 8480
rect 3191 8449 3203 8452
rect 3145 8443 3203 8449
rect 2222 8344 2228 8356
rect 2183 8316 2228 8344
rect 2222 8304 2228 8316
rect 2280 8304 2286 8356
rect 2332 8344 2360 8443
rect 3234 8440 3240 8452
rect 3292 8440 3298 8492
rect 3329 8483 3387 8489
rect 3329 8449 3341 8483
rect 3375 8449 3387 8483
rect 3329 8443 3387 8449
rect 3565 8483 3623 8489
rect 3565 8449 3577 8483
rect 3611 8480 3623 8483
rect 3694 8480 3700 8492
rect 3611 8452 3700 8480
rect 3611 8449 3623 8452
rect 3565 8443 3623 8449
rect 3344 8412 3372 8443
rect 3694 8440 3700 8452
rect 3752 8480 3758 8492
rect 3970 8480 3976 8492
rect 3752 8452 3976 8480
rect 3752 8440 3758 8452
rect 3970 8440 3976 8452
rect 4028 8480 4034 8492
rect 4065 8483 4123 8489
rect 4065 8480 4077 8483
rect 4028 8452 4077 8480
rect 4028 8440 4034 8452
rect 4065 8449 4077 8452
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4172 8412 4200 8511
rect 4706 8508 4712 8520
rect 4764 8508 4770 8560
rect 5169 8551 5227 8557
rect 5169 8517 5181 8551
rect 5215 8548 5227 8551
rect 6730 8548 6736 8560
rect 5215 8520 6736 8548
rect 5215 8517 5227 8520
rect 5169 8511 5227 8517
rect 6730 8508 6736 8520
rect 6788 8508 6794 8560
rect 9508 8557 9536 8588
rect 10042 8576 10048 8588
rect 10100 8616 10106 8628
rect 12618 8616 12624 8628
rect 10100 8588 11376 8616
rect 12579 8588 12624 8616
rect 10100 8576 10106 8588
rect 9401 8551 9459 8557
rect 9401 8517 9413 8551
rect 9447 8548 9459 8551
rect 9493 8551 9551 8557
rect 9493 8548 9505 8551
rect 9447 8520 9505 8548
rect 9447 8517 9459 8520
rect 9401 8511 9459 8517
rect 9493 8517 9505 8520
rect 9539 8517 9551 8551
rect 9493 8511 9551 8517
rect 9582 8508 9588 8560
rect 9640 8548 9646 8560
rect 9769 8551 9827 8557
rect 9769 8548 9781 8551
rect 9640 8520 9781 8548
rect 9640 8508 9646 8520
rect 9769 8517 9781 8520
rect 9815 8548 9827 8551
rect 10965 8551 11023 8557
rect 10965 8548 10977 8551
rect 9815 8520 10977 8548
rect 9815 8517 9827 8520
rect 9769 8511 9827 8517
rect 10965 8517 10977 8520
rect 11011 8517 11023 8551
rect 10965 8511 11023 8517
rect 4614 8480 4620 8492
rect 3344 8384 4200 8412
rect 4356 8452 4620 8480
rect 4356 8344 4384 8452
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 4890 8480 4896 8492
rect 4851 8452 4896 8480
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 5350 8489 5356 8492
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5313 8483 5356 8489
rect 5313 8449 5325 8483
rect 5313 8443 5356 8449
rect 4430 8372 4436 8424
rect 4488 8412 4494 8424
rect 5092 8412 5120 8443
rect 5350 8440 5356 8443
rect 5408 8440 5414 8492
rect 5902 8480 5908 8492
rect 5863 8452 5908 8480
rect 5902 8440 5908 8452
rect 5960 8480 5966 8492
rect 7190 8480 7196 8492
rect 5960 8452 7196 8480
rect 5960 8440 5966 8452
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 7466 8480 7472 8492
rect 7427 8452 7472 8480
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 8662 8480 8668 8492
rect 8623 8452 8668 8480
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 11348 8489 11376 8588
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 12710 8576 12716 8628
rect 12768 8616 12774 8628
rect 12805 8619 12863 8625
rect 12805 8616 12817 8619
rect 12768 8588 12817 8616
rect 12768 8576 12774 8588
rect 12805 8585 12817 8588
rect 12851 8585 12863 8619
rect 12805 8579 12863 8585
rect 12636 8548 12664 8576
rect 12894 8548 12900 8560
rect 12636 8520 12900 8548
rect 12894 8508 12900 8520
rect 12952 8548 12958 8560
rect 12952 8520 13308 8548
rect 12952 8508 12958 8520
rect 9217 8483 9275 8489
rect 9217 8480 9229 8483
rect 8772 8452 9229 8480
rect 7742 8412 7748 8424
rect 4488 8384 7748 8412
rect 4488 8372 4494 8384
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 8772 8356 8800 8452
rect 9217 8449 9229 8452
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8480 10471 8483
rect 11333 8483 11391 8489
rect 10459 8452 10548 8480
rect 10459 8449 10471 8452
rect 10413 8443 10471 8449
rect 10520 8424 10548 8452
rect 11333 8449 11345 8483
rect 11379 8449 11391 8483
rect 11333 8443 11391 8449
rect 11514 8440 11520 8492
rect 11572 8480 11578 8492
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 11572 8452 11713 8480
rect 11572 8440 11578 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 12529 8483 12587 8489
rect 12529 8480 12541 8483
rect 11931 8452 12541 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 12529 8449 12541 8452
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 13078 8440 13084 8492
rect 13136 8480 13142 8492
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 13136 8452 13185 8480
rect 13136 8440 13142 8452
rect 13173 8449 13185 8452
rect 13219 8449 13231 8483
rect 13280 8480 13308 8520
rect 13280 8452 13400 8480
rect 13173 8443 13231 8449
rect 10502 8412 10508 8424
rect 10463 8384 10508 8412
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 11057 8415 11115 8421
rect 11057 8381 11069 8415
rect 11103 8381 11115 8415
rect 11057 8375 11115 8381
rect 4798 8344 4804 8356
rect 2332 8316 4384 8344
rect 4759 8316 4804 8344
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 5258 8304 5264 8356
rect 5316 8344 5322 8356
rect 5445 8347 5503 8353
rect 5445 8344 5457 8347
rect 5316 8316 5457 8344
rect 5316 8304 5322 8316
rect 5445 8313 5457 8316
rect 5491 8313 5503 8347
rect 8754 8344 8760 8356
rect 8715 8316 8760 8344
rect 5445 8307 5503 8313
rect 8754 8304 8760 8316
rect 8812 8304 8818 8356
rect 11072 8344 11100 8375
rect 11790 8372 11796 8424
rect 11848 8412 11854 8424
rect 11977 8415 12035 8421
rect 11977 8412 11989 8415
rect 11848 8384 11989 8412
rect 11848 8372 11854 8384
rect 11977 8381 11989 8384
rect 12023 8381 12035 8415
rect 11977 8375 12035 8381
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8412 12495 8415
rect 12618 8412 12624 8424
rect 12483 8384 12624 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 12618 8372 12624 8384
rect 12676 8372 12682 8424
rect 13262 8412 13268 8424
rect 13223 8384 13268 8412
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 13372 8421 13400 8452
rect 13357 8415 13415 8421
rect 13357 8381 13369 8415
rect 13403 8381 13415 8415
rect 13357 8375 13415 8381
rect 11149 8347 11207 8353
rect 11149 8344 11161 8347
rect 11072 8316 11161 8344
rect 11149 8313 11161 8316
rect 11195 8313 11207 8347
rect 11149 8307 11207 8313
rect 3697 8279 3755 8285
rect 3697 8245 3709 8279
rect 3743 8276 3755 8279
rect 4062 8276 4068 8288
rect 3743 8248 4068 8276
rect 3743 8245 3755 8248
rect 3697 8239 3755 8245
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 4433 8279 4491 8285
rect 4433 8245 4445 8279
rect 4479 8276 4491 8279
rect 4614 8276 4620 8288
rect 4479 8248 4620 8276
rect 4479 8245 4491 8248
rect 4433 8239 4491 8245
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 1104 8186 13892 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 12214 8186
rect 12266 8134 12278 8186
rect 12330 8134 12342 8186
rect 12394 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 13892 8186
rect 1104 8112 13892 8134
rect 3145 8075 3203 8081
rect 3145 8041 3157 8075
rect 3191 8072 3203 8075
rect 3418 8072 3424 8084
rect 3191 8044 3424 8072
rect 3191 8041 3203 8044
rect 3145 8035 3203 8041
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 4706 8032 4712 8084
rect 4764 8072 4770 8084
rect 5537 8075 5595 8081
rect 5537 8072 5549 8075
rect 4764 8044 5549 8072
rect 4764 8032 4770 8044
rect 5537 8041 5549 8044
rect 5583 8041 5595 8075
rect 5537 8035 5595 8041
rect 9125 8075 9183 8081
rect 9125 8041 9137 8075
rect 9171 8072 9183 8075
rect 9306 8072 9312 8084
rect 9171 8044 9312 8072
rect 9171 8041 9183 8044
rect 9125 8035 9183 8041
rect 9306 8032 9312 8044
rect 9364 8032 9370 8084
rect 9493 8075 9551 8081
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 9950 8072 9956 8084
rect 9539 8044 9956 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 5074 7964 5080 8016
rect 5132 8004 5138 8016
rect 5813 8007 5871 8013
rect 5813 8004 5825 8007
rect 5132 7976 5825 8004
rect 5132 7964 5138 7976
rect 5813 7973 5825 7976
rect 5859 7973 5871 8007
rect 5813 7967 5871 7973
rect 8297 8007 8355 8013
rect 8297 7973 8309 8007
rect 8343 8004 8355 8007
rect 8754 8004 8760 8016
rect 8343 7976 8760 8004
rect 8343 7973 8355 7976
rect 8297 7967 8355 7973
rect 8754 7964 8760 7976
rect 8812 7964 8818 8016
rect 9214 7964 9220 8016
rect 9272 8004 9278 8016
rect 9508 8004 9536 8035
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 13262 8032 13268 8084
rect 13320 8072 13326 8084
rect 13449 8075 13507 8081
rect 13449 8072 13461 8075
rect 13320 8044 13461 8072
rect 13320 8032 13326 8044
rect 13449 8041 13461 8044
rect 13495 8041 13507 8075
rect 13449 8035 13507 8041
rect 9272 7976 9536 8004
rect 9585 8007 9643 8013
rect 9272 7964 9278 7976
rect 9585 7973 9597 8007
rect 9631 8004 9643 8007
rect 10042 8004 10048 8016
rect 9631 7976 10048 8004
rect 9631 7973 9643 7976
rect 9585 7967 9643 7973
rect 10042 7964 10048 7976
rect 10100 7964 10106 8016
rect 10505 8007 10563 8013
rect 10505 7973 10517 8007
rect 10551 8004 10563 8007
rect 11146 8004 11152 8016
rect 10551 7976 11152 8004
rect 10551 7973 10563 7976
rect 10505 7967 10563 7973
rect 11146 7964 11152 7976
rect 11204 7964 11210 8016
rect 12618 7964 12624 8016
rect 12676 8004 12682 8016
rect 13081 8007 13139 8013
rect 13081 8004 13093 8007
rect 12676 7976 13093 8004
rect 12676 7964 12682 7976
rect 13081 7973 13093 7976
rect 13127 7973 13139 8007
rect 13081 7967 13139 7973
rect 3789 7939 3847 7945
rect 3789 7936 3801 7939
rect 1412 7908 3801 7936
rect 1412 7880 1440 7908
rect 3789 7905 3801 7908
rect 3835 7905 3847 7939
rect 4062 7936 4068 7948
rect 4023 7908 4068 7936
rect 3789 7899 3847 7905
rect 4062 7896 4068 7908
rect 4120 7896 4126 7948
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 5350 7936 5356 7948
rect 4212 7908 5356 7936
rect 4212 7896 4218 7908
rect 5350 7896 5356 7908
rect 5408 7936 5414 7948
rect 7653 7939 7711 7945
rect 5408 7908 5948 7936
rect 5408 7896 5414 7908
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 5920 7877 5948 7908
rect 7653 7905 7665 7939
rect 7699 7936 7711 7939
rect 8389 7939 8447 7945
rect 8389 7936 8401 7939
rect 7699 7908 8401 7936
rect 7699 7905 7711 7908
rect 7653 7899 7711 7905
rect 8389 7905 8401 7908
rect 8435 7905 8447 7939
rect 8389 7899 8447 7905
rect 9490 7896 9496 7948
rect 9548 7936 9554 7948
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 9548 7908 9689 7936
rect 9548 7896 9554 7908
rect 9677 7905 9689 7908
rect 9723 7936 9735 7939
rect 9723 7908 10226 7936
rect 9723 7905 9735 7908
rect 9677 7899 9735 7905
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7837 5963 7871
rect 5905 7831 5963 7837
rect 6454 7828 6460 7880
rect 6512 7868 6518 7880
rect 6549 7871 6607 7877
rect 6549 7868 6561 7871
rect 6512 7840 6561 7868
rect 6512 7828 6518 7840
rect 6549 7837 6561 7840
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7868 6791 7871
rect 7098 7868 7104 7880
rect 6779 7840 7104 7868
rect 6779 7837 6791 7840
rect 6733 7831 6791 7837
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 7190 7828 7196 7880
rect 7248 7868 7254 7880
rect 7248 7840 7293 7868
rect 7248 7828 7254 7840
rect 7466 7828 7472 7880
rect 7524 7868 7530 7880
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7524 7840 7849 7868
rect 7524 7828 7530 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 8662 7868 8668 7880
rect 8623 7840 8668 7868
rect 7837 7831 7895 7837
rect 8662 7828 8668 7840
rect 8720 7828 8726 7880
rect 8938 7828 8944 7880
rect 8996 7868 9002 7880
rect 9398 7868 9404 7880
rect 8996 7840 9404 7868
rect 8996 7828 9002 7840
rect 9398 7828 9404 7840
rect 9456 7828 9462 7880
rect 10198 7877 10226 7908
rect 9769 7871 9827 7877
rect 9769 7837 9781 7871
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 10183 7871 10241 7877
rect 10183 7837 10195 7871
rect 10229 7837 10241 7871
rect 10183 7831 10241 7837
rect 1670 7800 1676 7812
rect 1631 7772 1676 7800
rect 1670 7760 1676 7772
rect 1728 7760 1734 7812
rect 2222 7760 2228 7812
rect 2280 7760 2286 7812
rect 4798 7760 4804 7812
rect 4856 7760 4862 7812
rect 6638 7760 6644 7812
rect 6696 7800 6702 7812
rect 6917 7803 6975 7809
rect 6917 7800 6929 7803
rect 6696 7772 6929 7800
rect 6696 7760 6702 7772
rect 6917 7769 6929 7772
rect 6963 7769 6975 7803
rect 6917 7763 6975 7769
rect 9122 7760 9128 7812
rect 9180 7800 9186 7812
rect 9784 7800 9812 7831
rect 10686 7828 10692 7880
rect 10744 7868 10750 7880
rect 10781 7871 10839 7877
rect 10781 7868 10793 7871
rect 10744 7840 10793 7868
rect 10744 7828 10750 7840
rect 10781 7837 10793 7840
rect 10827 7837 10839 7871
rect 11514 7868 11520 7880
rect 11475 7840 11520 7868
rect 10781 7831 10839 7837
rect 11514 7828 11520 7840
rect 11572 7828 11578 7880
rect 11790 7868 11796 7880
rect 11751 7840 11796 7868
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 13170 7868 13176 7880
rect 13131 7840 13176 7868
rect 13170 7828 13176 7840
rect 13228 7828 13234 7880
rect 9180 7772 9812 7800
rect 9953 7803 10011 7809
rect 9180 7760 9186 7772
rect 9953 7769 9965 7803
rect 9999 7800 10011 7803
rect 10042 7800 10048 7812
rect 9999 7772 10048 7800
rect 9999 7769 10011 7772
rect 9953 7763 10011 7769
rect 10042 7760 10048 7772
rect 10100 7760 10106 7812
rect 10318 7800 10324 7812
rect 10279 7772 10324 7800
rect 10318 7760 10324 7772
rect 10376 7760 10382 7812
rect 11701 7803 11759 7809
rect 11701 7769 11713 7803
rect 11747 7800 11759 7803
rect 13188 7800 13216 7828
rect 11747 7772 13216 7800
rect 11747 7769 11759 7772
rect 11701 7763 11759 7769
rect 11808 7744 11836 7772
rect 7006 7732 7012 7744
rect 6967 7704 7012 7732
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7558 7732 7564 7744
rect 7519 7704 7564 7732
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 7650 7692 7656 7744
rect 7708 7732 7714 7744
rect 8481 7735 8539 7741
rect 8481 7732 8493 7735
rect 7708 7704 8493 7732
rect 7708 7692 7714 7704
rect 8481 7701 8493 7704
rect 8527 7701 8539 7735
rect 8481 7695 8539 7701
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 10137 7735 10195 7741
rect 10137 7732 10149 7735
rect 8812 7704 10149 7732
rect 8812 7692 8818 7704
rect 10137 7701 10149 7704
rect 10183 7701 10195 7735
rect 10137 7695 10195 7701
rect 11790 7692 11796 7744
rect 11848 7692 11854 7744
rect 1104 7642 13892 7664
rect 1104 7590 8214 7642
rect 8266 7590 8278 7642
rect 8330 7590 8342 7642
rect 8394 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 13892 7642
rect 1104 7568 13892 7590
rect 1670 7488 1676 7540
rect 1728 7528 1734 7540
rect 3404 7531 3462 7537
rect 3404 7528 3416 7531
rect 1728 7500 3416 7528
rect 1728 7488 1734 7500
rect 3404 7497 3416 7500
rect 3450 7497 3462 7531
rect 3404 7491 3462 7497
rect 3510 7488 3516 7540
rect 3568 7528 3574 7540
rect 4062 7528 4068 7540
rect 3568 7500 4068 7528
rect 3568 7488 3574 7500
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 4614 7488 4620 7540
rect 4672 7488 4678 7540
rect 7926 7528 7932 7540
rect 4908 7500 7932 7528
rect 2314 7420 2320 7472
rect 2372 7420 2378 7472
rect 3697 7463 3755 7469
rect 3697 7460 3709 7463
rect 3436 7432 3709 7460
rect 3436 7404 3464 7432
rect 3697 7429 3709 7432
rect 3743 7429 3755 7463
rect 3697 7423 3755 7429
rect 3786 7420 3792 7472
rect 3844 7460 3850 7472
rect 4632 7460 4660 7488
rect 3844 7432 3889 7460
rect 4448 7432 4660 7460
rect 3844 7420 3850 7432
rect 3418 7352 3424 7404
rect 3476 7352 3482 7404
rect 3510 7352 3516 7404
rect 3568 7401 3574 7404
rect 3568 7395 3611 7401
rect 3599 7361 3611 7395
rect 3568 7355 3611 7361
rect 3568 7352 3574 7355
rect 1394 7324 1400 7336
rect 1355 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7284 1458 7336
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 2406 7324 2412 7336
rect 1719 7296 2412 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 3142 7324 3148 7336
rect 3055 7296 3148 7324
rect 3142 7284 3148 7296
rect 3200 7324 3206 7336
rect 3804 7324 3832 7420
rect 3970 7392 3976 7404
rect 3931 7364 3976 7392
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 4448 7401 4476 7432
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7361 4491 7395
rect 4598 7395 4656 7401
rect 4598 7392 4610 7395
rect 4433 7355 4491 7361
rect 4540 7364 4610 7392
rect 3200 7296 3832 7324
rect 3200 7284 3206 7296
rect 4540 7256 4568 7364
rect 4598 7361 4610 7364
rect 4644 7361 4656 7395
rect 4598 7355 4656 7361
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7392 4859 7395
rect 4908 7392 4936 7500
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 8570 7528 8576 7540
rect 8531 7500 8576 7528
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 9398 7528 9404 7540
rect 9359 7500 9404 7528
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 10870 7488 10876 7540
rect 10928 7528 10934 7540
rect 11057 7531 11115 7537
rect 11057 7528 11069 7531
rect 10928 7500 11069 7528
rect 10928 7488 10934 7500
rect 11057 7497 11069 7500
rect 11103 7497 11115 7531
rect 11057 7491 11115 7497
rect 11882 7488 11888 7540
rect 11940 7528 11946 7540
rect 11977 7531 12035 7537
rect 11977 7528 11989 7531
rect 11940 7500 11989 7528
rect 11940 7488 11946 7500
rect 11977 7497 11989 7500
rect 12023 7497 12035 7531
rect 11977 7491 12035 7497
rect 12437 7531 12495 7537
rect 12437 7497 12449 7531
rect 12483 7528 12495 7531
rect 12802 7528 12808 7540
rect 12483 7500 12808 7528
rect 12483 7497 12495 7500
rect 12437 7491 12495 7497
rect 12802 7488 12808 7500
rect 12860 7528 12866 7540
rect 12989 7531 13047 7537
rect 12989 7528 13001 7531
rect 12860 7500 13001 7528
rect 12860 7488 12866 7500
rect 12989 7497 13001 7500
rect 13035 7497 13047 7531
rect 12989 7491 13047 7497
rect 6454 7460 6460 7472
rect 5000 7432 6460 7460
rect 5000 7401 5028 7432
rect 6454 7420 6460 7432
rect 6512 7420 6518 7472
rect 7285 7463 7343 7469
rect 7285 7429 7297 7463
rect 7331 7460 7343 7463
rect 7558 7460 7564 7472
rect 7331 7432 7564 7460
rect 7331 7429 7343 7432
rect 7285 7423 7343 7429
rect 7558 7420 7564 7432
rect 7616 7460 7622 7472
rect 8113 7463 8171 7469
rect 8113 7460 8125 7463
rect 7616 7432 8125 7460
rect 7616 7420 7622 7432
rect 8113 7429 8125 7432
rect 8159 7429 8171 7463
rect 9306 7460 9312 7472
rect 8113 7423 8171 7429
rect 8864 7432 9312 7460
rect 4847 7364 4936 7392
rect 4985 7395 5043 7401
rect 4847 7361 4859 7364
rect 4801 7355 4859 7361
rect 4985 7361 4997 7395
rect 5031 7361 5043 7395
rect 4985 7355 5043 7361
rect 5074 7352 5080 7404
rect 5132 7392 5138 7404
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 5132 7364 5641 7392
rect 5132 7352 5138 7364
rect 5629 7361 5641 7364
rect 5675 7361 5687 7395
rect 5810 7392 5816 7404
rect 5771 7364 5816 7392
rect 5629 7355 5687 7361
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 5994 7392 6000 7404
rect 5955 7364 6000 7392
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 6730 7392 6736 7404
rect 6691 7364 6736 7392
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 7466 7392 7472 7404
rect 6871 7364 7472 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 8386 7392 8392 7404
rect 8347 7364 8392 7392
rect 8386 7352 8392 7364
rect 8444 7392 8450 7404
rect 8662 7392 8668 7404
rect 8444 7364 8668 7392
rect 8444 7352 8450 7364
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 8864 7401 8892 7432
rect 9306 7420 9312 7432
rect 9364 7420 9370 7472
rect 9416 7460 9444 7488
rect 9582 7460 9588 7472
rect 9416 7432 9588 7460
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 8849 7395 8907 7401
rect 8849 7361 8861 7395
rect 8895 7361 8907 7395
rect 8849 7355 8907 7361
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7392 9091 7395
rect 9416 7392 9444 7432
rect 9582 7420 9588 7432
rect 9640 7420 9646 7472
rect 9950 7420 9956 7472
rect 10008 7460 10014 7472
rect 10318 7460 10324 7472
rect 10008 7432 10324 7460
rect 10008 7420 10014 7432
rect 10318 7420 10324 7432
rect 10376 7460 10382 7472
rect 10689 7463 10747 7469
rect 10376 7432 10548 7460
rect 10376 7420 10382 7432
rect 9079 7364 9444 7392
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 4706 7324 4712 7336
rect 4667 7296 4712 7324
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 4890 7324 4896 7336
rect 4816 7296 4896 7324
rect 4816 7256 4844 7296
rect 4890 7284 4896 7296
rect 4948 7324 4954 7336
rect 6638 7324 6644 7336
rect 4948 7296 6644 7324
rect 4948 7284 4954 7296
rect 6638 7284 6644 7296
rect 6696 7284 6702 7336
rect 7377 7327 7435 7333
rect 7377 7293 7389 7327
rect 7423 7324 7435 7327
rect 7650 7324 7656 7336
rect 7423 7296 7656 7324
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 7650 7284 7656 7296
rect 7708 7284 7714 7336
rect 8772 7324 8800 7355
rect 9766 7352 9772 7404
rect 9824 7352 9830 7404
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 10042 7392 10048 7404
rect 9907 7364 10048 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 10042 7352 10048 7364
rect 10100 7352 10106 7404
rect 10520 7401 10548 7432
rect 10689 7429 10701 7463
rect 10735 7460 10747 7463
rect 12345 7463 12403 7469
rect 12345 7460 12357 7463
rect 10735 7432 12357 7460
rect 10735 7429 10747 7432
rect 10689 7423 10747 7429
rect 12345 7429 12357 7432
rect 12391 7429 12403 7463
rect 12894 7460 12900 7472
rect 12855 7432 12900 7460
rect 12345 7423 12403 7429
rect 12894 7420 12900 7432
rect 12952 7460 12958 7472
rect 13173 7463 13231 7469
rect 13173 7460 13185 7463
rect 12952 7432 13185 7460
rect 12952 7420 12958 7432
rect 13173 7429 13185 7432
rect 13219 7460 13231 7463
rect 13357 7463 13415 7469
rect 13357 7460 13369 7463
rect 13219 7432 13369 7460
rect 13219 7429 13231 7432
rect 13173 7423 13231 7429
rect 13357 7429 13369 7432
rect 13403 7429 13415 7463
rect 13357 7423 13415 7429
rect 10229 7395 10287 7401
rect 10229 7361 10241 7395
rect 10275 7361 10287 7395
rect 10229 7355 10287 7361
rect 10413 7395 10471 7401
rect 10413 7361 10425 7395
rect 10459 7361 10471 7395
rect 10413 7355 10471 7361
rect 10505 7395 10563 7401
rect 10505 7361 10517 7395
rect 10551 7361 10563 7395
rect 11790 7392 11796 7404
rect 11751 7364 11796 7392
rect 10505 7355 10563 7361
rect 9122 7324 9128 7336
rect 8680 7296 9128 7324
rect 8680 7268 8708 7296
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 9306 7284 9312 7336
rect 9364 7324 9370 7336
rect 9585 7327 9643 7333
rect 9585 7324 9597 7327
rect 9364 7296 9597 7324
rect 9364 7284 9370 7296
rect 9585 7293 9597 7296
rect 9631 7324 9643 7327
rect 9784 7324 9812 7352
rect 10244 7324 10272 7355
rect 9631 7296 10272 7324
rect 9631 7293 9643 7296
rect 9585 7287 9643 7293
rect 5718 7256 5724 7268
rect 4540 7228 4844 7256
rect 5679 7228 5724 7256
rect 5718 7216 5724 7228
rect 5776 7216 5782 7268
rect 8662 7256 8668 7268
rect 6656 7228 8668 7256
rect 4982 7148 4988 7200
rect 5040 7188 5046 7200
rect 5077 7191 5135 7197
rect 5077 7188 5089 7191
rect 5040 7160 5089 7188
rect 5040 7148 5046 7160
rect 5077 7157 5089 7160
rect 5123 7157 5135 7191
rect 5077 7151 5135 7157
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 6362 7188 6368 7200
rect 5868 7160 6368 7188
rect 5868 7148 5874 7160
rect 6362 7148 6368 7160
rect 6420 7188 6426 7200
rect 6656 7197 6684 7228
rect 8662 7216 8668 7228
rect 8720 7216 8726 7268
rect 8941 7259 8999 7265
rect 8941 7225 8953 7259
rect 8987 7256 8999 7259
rect 9030 7256 9036 7268
rect 8987 7228 9036 7256
rect 8987 7225 8999 7228
rect 8941 7219 8999 7225
rect 9030 7216 9036 7228
rect 9088 7216 9094 7268
rect 9769 7259 9827 7265
rect 9769 7225 9781 7259
rect 9815 7256 9827 7259
rect 9858 7256 9864 7268
rect 9815 7228 9864 7256
rect 9815 7225 9827 7228
rect 9769 7219 9827 7225
rect 9858 7216 9864 7228
rect 9916 7216 9922 7268
rect 10045 7259 10103 7265
rect 10045 7225 10057 7259
rect 10091 7256 10103 7259
rect 10226 7256 10232 7268
rect 10091 7228 10232 7256
rect 10091 7225 10103 7228
rect 10045 7219 10103 7225
rect 10226 7216 10232 7228
rect 10284 7256 10290 7268
rect 10321 7259 10379 7265
rect 10321 7256 10333 7259
rect 10284 7228 10333 7256
rect 10284 7216 10290 7228
rect 10321 7225 10333 7228
rect 10367 7225 10379 7259
rect 10321 7219 10379 7225
rect 6641 7191 6699 7197
rect 6641 7188 6653 7191
rect 6420 7160 6653 7188
rect 6420 7148 6426 7160
rect 6641 7157 6653 7160
rect 6687 7157 6699 7191
rect 9876 7188 9904 7216
rect 10428 7188 10456 7355
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 12621 7327 12679 7333
rect 12621 7293 12633 7327
rect 12667 7324 12679 7327
rect 12912 7324 12940 7420
rect 12667 7296 12940 7324
rect 12667 7293 12679 7296
rect 12621 7287 12679 7293
rect 11330 7188 11336 7200
rect 9876 7160 10456 7188
rect 11291 7160 11336 7188
rect 6641 7151 6699 7157
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11606 7188 11612 7200
rect 11567 7160 11612 7188
rect 11606 7148 11612 7160
rect 11664 7148 11670 7200
rect 1104 7098 13892 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 12214 7098
rect 12266 7046 12278 7098
rect 12330 7046 12342 7098
rect 12394 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 13892 7098
rect 1104 7024 13892 7046
rect 2314 6984 2320 6996
rect 2275 6956 2320 6984
rect 2314 6944 2320 6956
rect 2372 6944 2378 6996
rect 5718 6993 5724 6996
rect 4801 6987 4859 6993
rect 4801 6984 4813 6987
rect 4540 6956 4813 6984
rect 4540 6928 4568 6956
rect 4801 6953 4813 6956
rect 4847 6953 4859 6987
rect 4801 6947 4859 6953
rect 5708 6987 5724 6993
rect 5708 6953 5720 6987
rect 5708 6947 5724 6953
rect 5718 6944 5724 6947
rect 5776 6944 5782 6996
rect 8481 6987 8539 6993
rect 8481 6953 8493 6987
rect 8527 6984 8539 6987
rect 9490 6984 9496 6996
rect 8527 6956 9496 6984
rect 8527 6953 8539 6956
rect 8481 6947 8539 6953
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 10962 6984 10968 6996
rect 10923 6956 10968 6984
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 12253 6987 12311 6993
rect 12253 6953 12265 6987
rect 12299 6984 12311 6987
rect 12894 6984 12900 6996
rect 12299 6956 12900 6984
rect 12299 6953 12311 6956
rect 12253 6947 12311 6953
rect 12894 6944 12900 6956
rect 12952 6944 12958 6996
rect 13541 6987 13599 6993
rect 13541 6984 13553 6987
rect 13004 6956 13553 6984
rect 2406 6916 2412 6928
rect 2367 6888 2412 6916
rect 2406 6876 2412 6888
rect 2464 6876 2470 6928
rect 4522 6876 4528 6928
rect 4580 6876 4586 6928
rect 6730 6876 6736 6928
rect 6788 6916 6794 6928
rect 7193 6919 7251 6925
rect 7193 6916 7205 6919
rect 6788 6888 7205 6916
rect 6788 6876 6794 6888
rect 7193 6885 7205 6888
rect 7239 6916 7251 6919
rect 7239 6888 7972 6916
rect 7239 6885 7251 6888
rect 7193 6879 7251 6885
rect 3970 6808 3976 6860
rect 4028 6808 4034 6860
rect 4614 6848 4620 6860
rect 4356 6820 4620 6848
rect 2038 6740 2044 6792
rect 2096 6780 2102 6792
rect 2133 6783 2191 6789
rect 2133 6780 2145 6783
rect 2096 6752 2145 6780
rect 2096 6740 2102 6752
rect 2133 6749 2145 6752
rect 2179 6749 2191 6783
rect 2133 6743 2191 6749
rect 2593 6783 2651 6789
rect 2593 6749 2605 6783
rect 2639 6780 2651 6783
rect 3142 6780 3148 6792
rect 2639 6752 3148 6780
rect 2639 6749 2651 6752
rect 2593 6743 2651 6749
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 3988 6780 4016 6808
rect 3896 6752 4016 6780
rect 4060 6783 4118 6789
rect 2777 6715 2835 6721
rect 2777 6681 2789 6715
rect 2823 6712 2835 6715
rect 3896 6712 3924 6752
rect 4060 6749 4072 6783
rect 4106 6780 4118 6783
rect 4356 6780 4384 6820
rect 4614 6808 4620 6820
rect 4672 6808 4678 6860
rect 4890 6848 4896 6860
rect 4744 6820 4896 6848
rect 4106 6752 4384 6780
rect 4433 6783 4491 6789
rect 4106 6749 4118 6752
rect 4060 6743 4118 6749
rect 4433 6749 4445 6783
rect 4479 6780 4491 6783
rect 4744 6780 4772 6820
rect 4890 6808 4896 6820
rect 4948 6808 4954 6860
rect 5166 6848 5172 6860
rect 5000 6820 5172 6848
rect 5000 6789 5028 6820
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 5442 6808 5448 6860
rect 5500 6848 5506 6860
rect 5500 6820 5545 6848
rect 5500 6808 5506 6820
rect 7742 6808 7748 6860
rect 7800 6848 7806 6860
rect 7837 6851 7895 6857
rect 7837 6848 7849 6851
rect 7800 6820 7849 6848
rect 7800 6808 7806 6820
rect 7837 6817 7849 6820
rect 7883 6817 7895 6851
rect 7837 6811 7895 6817
rect 4479 6752 4772 6780
rect 4801 6783 4859 6789
rect 4479 6749 4491 6752
rect 4433 6743 4491 6749
rect 4801 6749 4813 6783
rect 4847 6749 4859 6783
rect 4801 6743 4859 6749
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5258 6780 5264 6792
rect 5123 6752 5264 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 4157 6715 4215 6721
rect 4157 6712 4169 6715
rect 2823 6684 3924 6712
rect 3988 6684 4169 6712
rect 2823 6681 2835 6684
rect 2777 6675 2835 6681
rect 3988 6656 4016 6684
rect 4157 6681 4169 6684
rect 4203 6681 4215 6715
rect 4157 6675 4215 6681
rect 4249 6715 4307 6721
rect 4249 6681 4261 6715
rect 4295 6712 4307 6715
rect 4816 6712 4844 6743
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 5353 6783 5411 6789
rect 5353 6749 5365 6783
rect 5399 6749 5411 6783
rect 7944 6780 7972 6888
rect 8386 6876 8392 6928
rect 8444 6916 8450 6928
rect 8941 6919 8999 6925
rect 8941 6916 8953 6919
rect 8444 6888 8953 6916
rect 8444 6876 8450 6888
rect 8941 6885 8953 6888
rect 8987 6885 8999 6919
rect 8941 6879 8999 6885
rect 9030 6876 9036 6928
rect 9088 6916 9094 6928
rect 9585 6919 9643 6925
rect 9585 6916 9597 6919
rect 9088 6888 9597 6916
rect 9088 6876 9094 6888
rect 9585 6885 9597 6888
rect 9631 6916 9643 6919
rect 10226 6916 10232 6928
rect 9631 6888 10232 6916
rect 9631 6885 9643 6888
rect 9585 6879 9643 6885
rect 10226 6876 10232 6888
rect 10284 6876 10290 6928
rect 10870 6916 10876 6928
rect 10428 6888 10876 6916
rect 8018 6808 8024 6860
rect 8076 6848 8082 6860
rect 8076 6820 8121 6848
rect 8076 6808 8082 6820
rect 9398 6808 9404 6860
rect 9456 6848 9462 6860
rect 9493 6851 9551 6857
rect 9493 6848 9505 6851
rect 9456 6820 9505 6848
rect 9456 6808 9462 6820
rect 9493 6817 9505 6820
rect 9539 6817 9551 6851
rect 9493 6811 9551 6817
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 9950 6848 9956 6860
rect 9723 6820 9956 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 9950 6808 9956 6820
rect 10008 6808 10014 6860
rect 10318 6808 10324 6860
rect 10376 6848 10382 6860
rect 10428 6857 10456 6888
rect 10870 6876 10876 6888
rect 10928 6876 10934 6928
rect 11514 6916 11520 6928
rect 11475 6888 11520 6916
rect 11514 6876 11520 6888
rect 11572 6876 11578 6928
rect 10413 6851 10471 6857
rect 10413 6848 10425 6851
rect 10376 6820 10425 6848
rect 10376 6808 10382 6820
rect 10413 6817 10425 6820
rect 10459 6817 10471 6851
rect 10413 6811 10471 6817
rect 10505 6851 10563 6857
rect 10505 6817 10517 6851
rect 10551 6848 10563 6851
rect 11330 6848 11336 6860
rect 10551 6820 11336 6848
rect 10551 6817 10563 6820
rect 10505 6811 10563 6817
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 11606 6848 11612 6860
rect 11567 6820 11612 6848
rect 11606 6808 11612 6820
rect 11664 6808 11670 6860
rect 8389 6783 8447 6789
rect 8389 6780 8401 6783
rect 7944 6752 8401 6780
rect 5353 6743 5411 6749
rect 8389 6749 8401 6752
rect 8435 6780 8447 6783
rect 8754 6780 8760 6792
rect 8435 6752 8760 6780
rect 8435 6749 8447 6752
rect 8389 6743 8447 6749
rect 5166 6712 5172 6724
rect 4295 6684 5172 6712
rect 4295 6681 4307 6684
rect 4249 6675 4307 6681
rect 3878 6653 3884 6656
rect 3873 6644 3884 6653
rect 3839 6616 3884 6644
rect 3873 6607 3884 6616
rect 3878 6604 3884 6607
rect 3936 6604 3942 6656
rect 3970 6604 3976 6656
rect 4028 6604 4034 6656
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 4264 6644 4292 6675
rect 5166 6672 5172 6684
rect 5224 6672 5230 6724
rect 5368 6712 5396 6743
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 8956 6752 9321 6780
rect 5626 6712 5632 6724
rect 5368 6684 5632 6712
rect 5626 6672 5632 6684
rect 5684 6672 5690 6724
rect 7006 6712 7012 6724
rect 6946 6684 7012 6712
rect 7006 6672 7012 6684
rect 7064 6672 7070 6724
rect 7926 6672 7932 6724
rect 7984 6712 7990 6724
rect 8205 6715 8263 6721
rect 8205 6712 8217 6715
rect 7984 6684 8217 6712
rect 7984 6672 7990 6684
rect 8205 6681 8217 6684
rect 8251 6681 8263 6715
rect 8205 6675 8263 6681
rect 8662 6672 8668 6724
rect 8720 6712 8726 6724
rect 8956 6712 8984 6752
rect 9309 6749 9321 6752
rect 9355 6749 9367 6783
rect 9766 6780 9772 6792
rect 9727 6752 9772 6780
rect 9309 6743 9367 6749
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 10686 6740 10692 6792
rect 10744 6780 10750 6792
rect 11057 6783 11115 6789
rect 11057 6780 11069 6783
rect 10744 6752 11069 6780
rect 10744 6740 10750 6752
rect 11057 6749 11069 6752
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 11146 6740 11152 6792
rect 11204 6780 11210 6792
rect 11701 6783 11759 6789
rect 11701 6780 11713 6783
rect 11204 6752 11713 6780
rect 11204 6740 11210 6752
rect 11701 6749 11713 6752
rect 11747 6749 11759 6783
rect 11701 6743 11759 6749
rect 11790 6740 11796 6792
rect 11848 6780 11854 6792
rect 11885 6783 11943 6789
rect 11885 6780 11897 6783
rect 11848 6752 11897 6780
rect 11848 6740 11854 6752
rect 11885 6749 11897 6752
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 12066 6740 12072 6792
rect 12124 6780 12130 6792
rect 12345 6783 12403 6789
rect 12345 6780 12357 6783
rect 12124 6752 12357 6780
rect 12124 6740 12130 6752
rect 12345 6749 12357 6752
rect 12391 6749 12403 6783
rect 12912 6780 12940 6944
rect 13004 6857 13032 6956
rect 13541 6953 13553 6956
rect 13587 6984 13599 6987
rect 14001 6987 14059 6993
rect 14001 6984 14013 6987
rect 13587 6956 14013 6984
rect 13587 6953 13599 6956
rect 13541 6947 13599 6953
rect 14001 6953 14013 6956
rect 14047 6953 14059 6987
rect 14001 6947 14059 6953
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6817 13047 6851
rect 12989 6811 13047 6817
rect 13081 6851 13139 6857
rect 13081 6817 13093 6851
rect 13127 6817 13139 6851
rect 13081 6811 13139 6817
rect 13096 6780 13124 6811
rect 13354 6780 13360 6792
rect 12912 6752 13360 6780
rect 12345 6743 12403 6749
rect 13354 6740 13360 6752
rect 13412 6740 13418 6792
rect 9122 6712 9128 6724
rect 8720 6684 8984 6712
rect 9083 6684 9128 6712
rect 8720 6672 8726 6684
rect 9122 6672 9128 6684
rect 9180 6672 9186 6724
rect 9490 6672 9496 6724
rect 9548 6712 9554 6724
rect 9858 6712 9864 6724
rect 9548 6684 9864 6712
rect 9548 6672 9554 6684
rect 9646 6656 9674 6684
rect 9858 6672 9864 6684
rect 9916 6672 9922 6724
rect 10045 6715 10103 6721
rect 10045 6681 10057 6715
rect 10091 6712 10103 6715
rect 12897 6715 12955 6721
rect 12897 6712 12909 6715
rect 10091 6684 12909 6712
rect 10091 6681 10103 6684
rect 10045 6675 10103 6681
rect 12897 6681 12909 6684
rect 12943 6681 12955 6715
rect 12897 6675 12955 6681
rect 4120 6616 4292 6644
rect 4617 6647 4675 6653
rect 4120 6604 4126 6616
rect 4617 6613 4629 6647
rect 4663 6644 4675 6647
rect 5077 6647 5135 6653
rect 5077 6644 5089 6647
rect 4663 6616 5089 6644
rect 4663 6613 4675 6616
rect 4617 6607 4675 6613
rect 5077 6613 5089 6616
rect 5123 6613 5135 6647
rect 5077 6607 5135 6613
rect 5261 6647 5319 6653
rect 5261 6613 5273 6647
rect 5307 6644 5319 6647
rect 5718 6644 5724 6656
rect 5307 6616 5724 6644
rect 5307 6613 5319 6616
rect 5261 6607 5319 6613
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 7374 6644 7380 6656
rect 7335 6616 7380 6644
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 7742 6644 7748 6656
rect 7703 6616 7748 6644
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 8018 6604 8024 6656
rect 8076 6644 8082 6656
rect 8570 6644 8576 6656
rect 8076 6616 8576 6644
rect 8076 6604 8082 6616
rect 8570 6604 8576 6616
rect 8628 6644 8634 6656
rect 8757 6647 8815 6653
rect 8757 6644 8769 6647
rect 8628 6616 8769 6644
rect 8628 6604 8634 6616
rect 8757 6613 8769 6616
rect 8803 6644 8815 6647
rect 8938 6644 8944 6656
rect 8803 6616 8944 6644
rect 8803 6613 8815 6616
rect 8757 6607 8815 6613
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 9646 6616 9680 6656
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 10134 6604 10140 6656
rect 10192 6644 10198 6656
rect 10597 6647 10655 6653
rect 10597 6644 10609 6647
rect 10192 6616 10609 6644
rect 10192 6604 10198 6616
rect 10597 6613 10609 6616
rect 10643 6613 10655 6647
rect 11974 6644 11980 6656
rect 11935 6616 11980 6644
rect 10597 6607 10655 6613
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12529 6647 12587 6653
rect 12529 6613 12541 6647
rect 12575 6644 12587 6647
rect 12618 6644 12624 6656
rect 12575 6616 12624 6644
rect 12575 6613 12587 6616
rect 12529 6607 12587 6613
rect 12618 6604 12624 6616
rect 12676 6604 12682 6656
rect 1104 6554 13892 6576
rect 1104 6502 8214 6554
rect 8266 6502 8278 6554
rect 8330 6502 8342 6554
rect 8394 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 13892 6554
rect 1104 6480 13892 6502
rect 3888 6412 4103 6440
rect 2222 6332 2228 6384
rect 2280 6332 2286 6384
rect 3418 6304 3424 6316
rect 3379 6276 3424 6304
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 3602 6304 3608 6316
rect 3563 6276 3608 6304
rect 3602 6264 3608 6276
rect 3660 6264 3666 6316
rect 3888 6313 3916 6412
rect 4075 6372 4103 6412
rect 4890 6400 4896 6452
rect 4948 6440 4954 6452
rect 4948 6412 4993 6440
rect 4948 6400 4954 6412
rect 5074 6400 5080 6452
rect 5132 6400 5138 6452
rect 5994 6440 6000 6452
rect 5955 6412 6000 6440
rect 5994 6400 6000 6412
rect 6052 6400 6058 6452
rect 7466 6400 7472 6452
rect 7524 6440 7530 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 7524 6412 7849 6440
rect 7524 6400 7530 6412
rect 7837 6409 7849 6412
rect 7883 6409 7895 6443
rect 8846 6440 8852 6452
rect 8807 6412 8852 6440
rect 7837 6403 7895 6409
rect 8846 6400 8852 6412
rect 8904 6400 8910 6452
rect 8938 6400 8944 6452
rect 8996 6440 9002 6452
rect 9769 6443 9827 6449
rect 9769 6440 9781 6443
rect 8996 6412 9781 6440
rect 8996 6400 9002 6412
rect 9769 6409 9781 6412
rect 9815 6440 9827 6443
rect 9953 6443 10011 6449
rect 9953 6440 9965 6443
rect 9815 6412 9965 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 9953 6409 9965 6412
rect 9999 6440 10011 6443
rect 10318 6440 10324 6452
rect 9999 6412 10324 6440
rect 9999 6409 10011 6412
rect 9953 6403 10011 6409
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 11885 6443 11943 6449
rect 11885 6440 11897 6443
rect 10428 6412 11897 6440
rect 5092 6372 5120 6400
rect 5718 6372 5724 6384
rect 4075 6344 5120 6372
rect 5679 6344 5724 6372
rect 5718 6332 5724 6344
rect 5776 6332 5782 6384
rect 7098 6332 7104 6384
rect 7156 6372 7162 6384
rect 7742 6372 7748 6384
rect 7156 6344 7748 6372
rect 7156 6332 7162 6344
rect 7742 6332 7748 6344
rect 7800 6332 7806 6384
rect 10428 6372 10456 6412
rect 11885 6409 11897 6412
rect 11931 6409 11943 6443
rect 11885 6403 11943 6409
rect 11974 6400 11980 6452
rect 12032 6440 12038 6452
rect 13262 6440 13268 6452
rect 12032 6412 12664 6440
rect 13223 6412 13268 6440
rect 12032 6400 12038 6412
rect 11054 6372 11060 6384
rect 7852 6344 10456 6372
rect 4154 6313 4160 6316
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6273 3939 6307
rect 3881 6267 3939 6273
rect 4111 6307 4160 6313
rect 4111 6273 4123 6307
rect 4157 6273 4160 6307
rect 4111 6267 4160 6273
rect 4154 6264 4160 6267
rect 4212 6264 4218 6316
rect 4522 6304 4528 6316
rect 4264 6276 4528 6304
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 3697 6239 3755 6245
rect 3697 6236 3709 6239
rect 1719 6208 3709 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 3697 6205 3709 6208
rect 3743 6205 3755 6239
rect 3697 6199 3755 6205
rect 3786 6196 3792 6248
rect 3844 6236 3850 6248
rect 4264 6245 4292 6276
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6273 5135 6307
rect 5077 6267 5135 6273
rect 4249 6239 4307 6245
rect 4249 6236 4261 6239
rect 3844 6208 4261 6236
rect 3844 6196 3850 6208
rect 4249 6205 4261 6208
rect 4295 6205 4307 6239
rect 4249 6199 4307 6205
rect 4341 6239 4399 6245
rect 4341 6205 4353 6239
rect 4387 6236 4399 6239
rect 4632 6236 4660 6267
rect 4729 6239 4787 6245
rect 4729 6236 4741 6239
rect 4387 6208 4660 6236
rect 4387 6205 4399 6208
rect 4341 6199 4399 6205
rect 4724 6205 4741 6236
rect 4775 6205 4787 6239
rect 4724 6199 4787 6205
rect 3878 6128 3884 6180
rect 3936 6168 3942 6180
rect 4356 6168 4384 6199
rect 3936 6140 4384 6168
rect 3936 6128 3942 6140
rect 4522 6128 4528 6180
rect 4580 6168 4586 6180
rect 4724 6168 4752 6199
rect 4580 6140 4752 6168
rect 4580 6128 4586 6140
rect 3145 6103 3203 6109
rect 3145 6069 3157 6103
rect 3191 6100 3203 6103
rect 3970 6100 3976 6112
rect 3191 6072 3976 6100
rect 3191 6069 3203 6072
rect 3145 6063 3203 6069
rect 3970 6060 3976 6072
rect 4028 6100 4034 6112
rect 5092 6100 5120 6267
rect 5166 6264 5172 6316
rect 5224 6304 5230 6316
rect 5350 6304 5356 6316
rect 5224 6276 5269 6304
rect 5311 6276 5356 6304
rect 5224 6264 5230 6276
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 5501 6307 5559 6313
rect 5501 6273 5513 6307
rect 5547 6304 5559 6307
rect 5547 6273 5580 6304
rect 5501 6267 5580 6273
rect 5552 6236 5580 6267
rect 5626 6264 5632 6316
rect 5684 6304 5690 6316
rect 5859 6307 5917 6313
rect 5684 6276 5729 6304
rect 5684 6264 5690 6276
rect 5859 6273 5871 6307
rect 5905 6304 5917 6307
rect 6086 6304 6092 6316
rect 5905 6276 6092 6304
rect 5905 6273 5917 6276
rect 5859 6267 5917 6273
rect 6086 6264 6092 6276
rect 6144 6264 6150 6316
rect 6362 6304 6368 6316
rect 6323 6276 6368 6304
rect 6362 6264 6368 6276
rect 6420 6264 6426 6316
rect 6638 6304 6644 6316
rect 6599 6276 6644 6304
rect 6638 6264 6644 6276
rect 6696 6264 6702 6316
rect 6730 6264 6736 6316
rect 6788 6304 6794 6316
rect 6788 6276 6833 6304
rect 6788 6264 6794 6276
rect 7190 6264 7196 6316
rect 7248 6304 7254 6316
rect 7285 6307 7343 6313
rect 7285 6304 7297 6307
rect 7248 6276 7297 6304
rect 7248 6264 7254 6276
rect 7285 6273 7297 6276
rect 7331 6273 7343 6307
rect 7466 6304 7472 6316
rect 7427 6276 7472 6304
rect 7285 6267 7343 6273
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 6270 6236 6276 6248
rect 5552 6208 6276 6236
rect 6270 6196 6276 6208
rect 6328 6196 6334 6248
rect 7852 6236 7880 6344
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 8260 6276 8305 6304
rect 8260 6264 8266 6276
rect 8386 6264 8392 6316
rect 8444 6304 8450 6316
rect 9030 6304 9036 6316
rect 8444 6276 9036 6304
rect 8444 6264 8450 6276
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9306 6304 9312 6316
rect 9267 6276 9312 6304
rect 9306 6264 9312 6276
rect 9364 6264 9370 6316
rect 10428 6313 10456 6344
rect 10704 6344 11060 6372
rect 10704 6313 10732 6344
rect 11054 6332 11060 6344
rect 11112 6332 11118 6384
rect 12526 6372 12532 6384
rect 11164 6344 12434 6372
rect 12487 6344 12532 6372
rect 11164 6313 11192 6344
rect 10413 6307 10471 6313
rect 10413 6273 10425 6307
rect 10459 6273 10471 6307
rect 10413 6267 10471 6273
rect 10689 6307 10747 6313
rect 10689 6273 10701 6307
rect 10735 6273 10747 6307
rect 10689 6267 10747 6273
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6304 10839 6307
rect 11149 6307 11207 6313
rect 11149 6304 11161 6307
rect 10827 6276 11161 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 11149 6273 11161 6276
rect 11195 6273 11207 6307
rect 12406 6304 12434 6344
rect 12526 6332 12532 6344
rect 12584 6332 12590 6384
rect 12636 6372 12664 6412
rect 13262 6400 13268 6412
rect 13320 6400 13326 6452
rect 13173 6375 13231 6381
rect 13173 6372 13185 6375
rect 12636 6344 13185 6372
rect 13173 6341 13185 6344
rect 13219 6341 13231 6375
rect 13173 6335 13231 6341
rect 13078 6304 13084 6316
rect 11149 6267 11207 6273
rect 11256 6276 12112 6304
rect 12406 6276 13084 6304
rect 8294 6236 8300 6248
rect 7300 6208 7880 6236
rect 8255 6208 8300 6236
rect 7300 6180 7328 6208
rect 8294 6196 8300 6208
rect 8352 6196 8358 6248
rect 8481 6239 8539 6245
rect 8481 6205 8493 6239
rect 8527 6236 8539 6239
rect 8570 6236 8576 6248
rect 8527 6208 8576 6236
rect 8527 6205 8539 6208
rect 8481 6199 8539 6205
rect 8570 6196 8576 6208
rect 8628 6196 8634 6248
rect 9217 6239 9275 6245
rect 9217 6236 9229 6239
rect 8772 6208 9229 6236
rect 5626 6128 5632 6180
rect 5684 6168 5690 6180
rect 6730 6168 6736 6180
rect 5684 6140 6736 6168
rect 5684 6128 5690 6140
rect 6730 6128 6736 6140
rect 6788 6168 6794 6180
rect 6917 6171 6975 6177
rect 6917 6168 6929 6171
rect 6788 6140 6929 6168
rect 6788 6128 6794 6140
rect 6917 6137 6929 6140
rect 6963 6137 6975 6171
rect 7098 6168 7104 6180
rect 7059 6140 7104 6168
rect 6917 6131 6975 6137
rect 7098 6128 7104 6140
rect 7156 6128 7162 6180
rect 7282 6128 7288 6180
rect 7340 6128 7346 6180
rect 7650 6168 7656 6180
rect 7611 6140 7656 6168
rect 7650 6128 7656 6140
rect 7708 6128 7714 6180
rect 8018 6128 8024 6180
rect 8076 6168 8082 6180
rect 8772 6168 8800 6208
rect 9217 6205 9229 6208
rect 9263 6205 9275 6239
rect 9217 6199 9275 6205
rect 9490 6196 9496 6248
rect 9548 6236 9554 6248
rect 10870 6236 10876 6248
rect 9548 6208 10876 6236
rect 9548 6196 9554 6208
rect 10870 6196 10876 6208
rect 10928 6196 10934 6248
rect 8076 6140 8800 6168
rect 9129 6171 9187 6177
rect 8076 6128 8082 6140
rect 9129 6137 9141 6171
rect 9175 6168 9187 6171
rect 9674 6168 9680 6180
rect 9175 6140 9680 6168
rect 9175 6137 9187 6140
rect 9129 6131 9187 6137
rect 9674 6128 9680 6140
rect 9732 6128 9738 6180
rect 10226 6128 10232 6180
rect 10284 6168 10290 6180
rect 11256 6168 11284 6276
rect 11333 6239 11391 6245
rect 11333 6205 11345 6239
rect 11379 6205 11391 6239
rect 11974 6236 11980 6248
rect 11935 6208 11980 6236
rect 11333 6199 11391 6205
rect 10284 6140 11284 6168
rect 11348 6168 11376 6199
rect 11974 6196 11980 6208
rect 12032 6196 12038 6248
rect 12084 6245 12112 6276
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 12069 6239 12127 6245
rect 12069 6205 12081 6239
rect 12115 6205 12127 6239
rect 13354 6236 13360 6248
rect 13315 6208 13360 6236
rect 12069 6199 12127 6205
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 11517 6171 11575 6177
rect 11517 6168 11529 6171
rect 11348 6140 11529 6168
rect 10284 6128 10290 6140
rect 11517 6137 11529 6140
rect 11563 6137 11575 6171
rect 11517 6131 11575 6137
rect 12713 6171 12771 6177
rect 12713 6137 12725 6171
rect 12759 6168 12771 6171
rect 12894 6168 12900 6180
rect 12759 6140 12900 6168
rect 12759 6137 12771 6140
rect 12713 6131 12771 6137
rect 12894 6128 12900 6140
rect 12952 6128 12958 6180
rect 4028 6072 5120 6100
rect 4028 6060 4034 6072
rect 5442 6060 5448 6112
rect 5500 6100 5506 6112
rect 6457 6103 6515 6109
rect 6457 6100 6469 6103
rect 5500 6072 6469 6100
rect 5500 6060 5506 6072
rect 6457 6069 6469 6072
rect 6503 6069 6515 6103
rect 6457 6063 6515 6069
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 9490 6100 9496 6112
rect 8352 6072 9496 6100
rect 8352 6060 8358 6072
rect 9490 6060 9496 6072
rect 9548 6060 9554 6112
rect 10042 6100 10048 6112
rect 10003 6072 10048 6100
rect 10042 6060 10048 6072
rect 10100 6060 10106 6112
rect 10321 6103 10379 6109
rect 10321 6069 10333 6103
rect 10367 6100 10379 6103
rect 10870 6100 10876 6112
rect 10367 6072 10876 6100
rect 10367 6069 10379 6072
rect 10321 6063 10379 6069
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 10965 6103 11023 6109
rect 10965 6069 10977 6103
rect 11011 6100 11023 6103
rect 11882 6100 11888 6112
rect 11011 6072 11888 6100
rect 11011 6069 11023 6072
rect 10965 6063 11023 6069
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 12805 6103 12863 6109
rect 12805 6069 12817 6103
rect 12851 6100 12863 6103
rect 14001 6103 14059 6109
rect 14001 6100 14013 6103
rect 12851 6072 14013 6100
rect 12851 6069 12863 6072
rect 12805 6063 12863 6069
rect 14001 6069 14013 6072
rect 14047 6069 14059 6103
rect 14001 6063 14059 6069
rect 1104 6010 13892 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 12214 6010
rect 12266 5958 12278 6010
rect 12330 5958 12342 6010
rect 12394 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 13892 6010
rect 1104 5936 13892 5958
rect 2222 5896 2228 5908
rect 2183 5868 2228 5896
rect 2222 5856 2228 5868
rect 2280 5856 2286 5908
rect 3881 5899 3939 5905
rect 3881 5865 3893 5899
rect 3927 5865 3939 5899
rect 3881 5859 3939 5865
rect 4249 5899 4307 5905
rect 4249 5865 4261 5899
rect 4295 5896 4307 5899
rect 4706 5896 4712 5908
rect 4295 5868 4712 5896
rect 4295 5865 4307 5868
rect 4249 5859 4307 5865
rect 3896 5760 3924 5859
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 5074 5896 5080 5908
rect 4816 5868 5080 5896
rect 4430 5788 4436 5840
rect 4488 5828 4494 5840
rect 4525 5831 4583 5837
rect 4525 5828 4537 5831
rect 4488 5800 4537 5828
rect 4488 5788 4494 5800
rect 4525 5797 4537 5800
rect 4571 5828 4583 5831
rect 4816 5828 4844 5868
rect 5074 5856 5080 5868
rect 5132 5856 5138 5908
rect 6086 5896 6092 5908
rect 6047 5868 6092 5896
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 6270 5856 6276 5908
rect 6328 5896 6334 5908
rect 6733 5899 6791 5905
rect 6733 5896 6745 5899
rect 6328 5868 6745 5896
rect 6328 5856 6334 5868
rect 6733 5865 6745 5868
rect 6779 5865 6791 5899
rect 6733 5859 6791 5865
rect 6917 5899 6975 5905
rect 6917 5865 6929 5899
rect 6963 5896 6975 5899
rect 7193 5899 7251 5905
rect 7193 5896 7205 5899
rect 6963 5868 7205 5896
rect 6963 5865 6975 5868
rect 6917 5859 6975 5865
rect 7193 5865 7205 5868
rect 7239 5896 7251 5899
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 7239 5868 7849 5896
rect 7239 5865 7251 5868
rect 7193 5859 7251 5865
rect 7837 5865 7849 5868
rect 7883 5896 7895 5899
rect 7926 5896 7932 5908
rect 7883 5868 7932 5896
rect 7883 5865 7895 5868
rect 7837 5859 7895 5865
rect 7926 5856 7932 5868
rect 7984 5856 7990 5908
rect 8018 5856 8024 5908
rect 8076 5896 8082 5908
rect 8205 5899 8263 5905
rect 8076 5868 8121 5896
rect 8076 5856 8082 5868
rect 8205 5865 8217 5899
rect 8251 5865 8263 5899
rect 8205 5859 8263 5865
rect 4571 5800 4844 5828
rect 4893 5831 4951 5837
rect 4571 5797 4583 5800
rect 4525 5791 4583 5797
rect 4893 5797 4905 5831
rect 4939 5828 4951 5831
rect 5166 5828 5172 5840
rect 4939 5800 5172 5828
rect 4939 5797 4951 5800
rect 4893 5791 4951 5797
rect 5166 5788 5172 5800
rect 5224 5788 5230 5840
rect 5258 5788 5264 5840
rect 5316 5828 5322 5840
rect 5353 5831 5411 5837
rect 5353 5828 5365 5831
rect 5316 5800 5365 5828
rect 5316 5788 5322 5800
rect 5353 5797 5365 5800
rect 5399 5797 5411 5831
rect 5353 5791 5411 5797
rect 5644 5800 7144 5828
rect 3160 5732 3924 5760
rect 3160 5704 3188 5732
rect 3970 5720 3976 5772
rect 4028 5760 4034 5772
rect 4028 5732 4073 5760
rect 4028 5720 4034 5732
rect 2038 5692 2044 5704
rect 1999 5664 2044 5692
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 3142 5692 3148 5704
rect 3055 5664 3148 5692
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5692 3663 5695
rect 3694 5692 3700 5704
rect 3651 5664 3700 5692
rect 3651 5661 3663 5664
rect 3605 5655 3663 5661
rect 3694 5652 3700 5664
rect 3752 5652 3758 5704
rect 3881 5695 3939 5701
rect 3881 5661 3893 5695
rect 3927 5692 3939 5695
rect 4522 5692 4528 5704
rect 3927 5664 4528 5692
rect 3927 5661 3939 5664
rect 3881 5655 3939 5661
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 4706 5692 4712 5704
rect 4667 5664 4712 5692
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 4798 5652 4804 5704
rect 4856 5692 4862 5704
rect 4856 5664 4901 5692
rect 4856 5652 4862 5664
rect 4982 5652 4988 5704
rect 5040 5692 5046 5704
rect 5442 5692 5448 5704
rect 5500 5701 5506 5704
rect 5500 5695 5543 5701
rect 5040 5664 5085 5692
rect 5184 5664 5448 5692
rect 5040 5652 5046 5664
rect 3513 5627 3571 5633
rect 3513 5593 3525 5627
rect 3559 5624 3571 5627
rect 4614 5624 4620 5636
rect 3559 5596 4620 5624
rect 3559 5593 3571 5596
rect 3513 5587 3571 5593
rect 4614 5584 4620 5596
rect 4672 5624 4678 5636
rect 4816 5624 4844 5652
rect 5184 5624 5212 5664
rect 5442 5652 5448 5664
rect 5531 5661 5543 5695
rect 5500 5655 5543 5661
rect 5500 5652 5506 5655
rect 4672 5596 5212 5624
rect 4672 5584 4678 5596
rect 5350 5584 5356 5636
rect 5408 5624 5414 5636
rect 5644 5633 5672 5800
rect 6086 5720 6092 5772
rect 6144 5760 6150 5772
rect 7116 5760 7144 5800
rect 7282 5788 7288 5840
rect 7340 5828 7346 5840
rect 7469 5831 7527 5837
rect 7469 5828 7481 5831
rect 7340 5800 7481 5828
rect 7340 5788 7346 5800
rect 7469 5797 7481 5800
rect 7515 5797 7527 5831
rect 8220 5828 8248 5859
rect 8294 5856 8300 5908
rect 8352 5896 8358 5908
rect 9585 5899 9643 5905
rect 9585 5896 9597 5899
rect 8352 5868 9597 5896
rect 8352 5856 8358 5868
rect 9585 5865 9597 5868
rect 9631 5865 9643 5899
rect 10502 5896 10508 5908
rect 10463 5868 10508 5896
rect 9585 5859 9643 5865
rect 10502 5856 10508 5868
rect 10560 5856 10566 5908
rect 10686 5896 10692 5908
rect 10647 5868 10692 5896
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 11698 5856 11704 5908
rect 11756 5896 11762 5908
rect 12253 5899 12311 5905
rect 12253 5896 12265 5899
rect 11756 5868 12265 5896
rect 11756 5856 11762 5868
rect 12253 5865 12265 5868
rect 12299 5865 12311 5899
rect 12253 5859 12311 5865
rect 13262 5856 13268 5908
rect 13320 5896 13326 5908
rect 13449 5899 13507 5905
rect 13449 5896 13461 5899
rect 13320 5868 13461 5896
rect 13320 5856 13326 5868
rect 13449 5865 13461 5868
rect 13495 5865 13507 5899
rect 13449 5859 13507 5865
rect 7469 5791 7527 5797
rect 7668 5800 8248 5828
rect 9309 5831 9367 5837
rect 7668 5772 7696 5800
rect 9309 5797 9321 5831
rect 9355 5828 9367 5831
rect 9674 5828 9680 5840
rect 9355 5800 9680 5828
rect 9355 5797 9367 5800
rect 9309 5791 9367 5797
rect 9674 5788 9680 5800
rect 9732 5828 9738 5840
rect 10226 5828 10232 5840
rect 9732 5800 10232 5828
rect 9732 5788 9738 5800
rect 10226 5788 10232 5800
rect 10284 5828 10290 5840
rect 11146 5828 11152 5840
rect 10284 5800 11152 5828
rect 10284 5788 10290 5800
rect 11146 5788 11152 5800
rect 11204 5788 11210 5840
rect 12437 5831 12495 5837
rect 12437 5797 12449 5831
rect 12483 5828 12495 5831
rect 13354 5828 13360 5840
rect 12483 5800 13360 5828
rect 12483 5797 12495 5800
rect 12437 5791 12495 5797
rect 13354 5788 13360 5800
rect 13412 5788 13418 5840
rect 7650 5760 7656 5772
rect 6144 5732 6684 5760
rect 6144 5720 6150 5732
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5692 5963 5695
rect 6365 5695 6423 5701
rect 6365 5692 6377 5695
rect 5951 5664 6377 5692
rect 5951 5661 5963 5664
rect 5905 5655 5963 5661
rect 6365 5661 6377 5664
rect 6411 5692 6423 5695
rect 6454 5692 6460 5704
rect 6411 5664 6460 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 6656 5701 6684 5732
rect 7116 5732 7656 5760
rect 7116 5701 7144 5732
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 7745 5763 7803 5769
rect 7745 5729 7757 5763
rect 7791 5760 7803 5763
rect 8389 5763 8447 5769
rect 7791 5732 8156 5760
rect 7791 5729 7803 5732
rect 7745 5723 7803 5729
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5661 6607 5695
rect 6549 5655 6607 5661
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5661 6699 5695
rect 6641 5655 6699 5661
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5661 7159 5695
rect 7101 5655 7159 5661
rect 5629 5627 5687 5633
rect 5629 5624 5641 5627
rect 5408 5596 5641 5624
rect 5408 5584 5414 5596
rect 5629 5593 5641 5596
rect 5675 5593 5687 5627
rect 5629 5587 5687 5593
rect 5721 5627 5779 5633
rect 5721 5593 5733 5627
rect 5767 5593 5779 5627
rect 5721 5587 5779 5593
rect 5997 5627 6055 5633
rect 5997 5593 6009 5627
rect 6043 5624 6055 5627
rect 6178 5624 6184 5636
rect 6043 5596 6184 5624
rect 6043 5593 6055 5596
rect 5997 5587 6055 5593
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 3237 5559 3295 5565
rect 3237 5556 3249 5559
rect 2924 5528 3249 5556
rect 2924 5516 2930 5528
rect 3237 5525 3249 5528
rect 3283 5525 3295 5559
rect 5736 5556 5764 5587
rect 6178 5584 6184 5596
rect 6236 5584 6242 5636
rect 6564 5624 6592 5655
rect 7834 5652 7840 5704
rect 7892 5692 7898 5704
rect 7929 5695 7987 5701
rect 7929 5692 7941 5695
rect 7892 5664 7941 5692
rect 7892 5652 7898 5664
rect 7929 5661 7941 5664
rect 7975 5661 7987 5695
rect 8128 5692 8156 5732
rect 8389 5729 8401 5763
rect 8435 5760 8447 5763
rect 8754 5760 8760 5772
rect 8435 5732 8760 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 8754 5720 8760 5732
rect 8812 5720 8818 5772
rect 9217 5763 9275 5769
rect 9217 5729 9229 5763
rect 9263 5760 9275 5763
rect 9582 5760 9588 5772
rect 9263 5732 9588 5760
rect 9263 5729 9275 5732
rect 9217 5723 9275 5729
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 9953 5763 10011 5769
rect 9953 5729 9965 5763
rect 9999 5760 10011 5763
rect 10778 5760 10784 5772
rect 9999 5732 10784 5760
rect 9999 5729 10011 5732
rect 9953 5723 10011 5729
rect 10778 5720 10784 5732
rect 10836 5760 10842 5772
rect 11238 5760 11244 5772
rect 10836 5732 11244 5760
rect 10836 5720 10842 5732
rect 11238 5720 11244 5732
rect 11296 5760 11302 5772
rect 11333 5763 11391 5769
rect 11333 5760 11345 5763
rect 11296 5732 11345 5760
rect 11296 5720 11302 5732
rect 11333 5729 11345 5732
rect 11379 5760 11391 5763
rect 11609 5763 11667 5769
rect 11609 5760 11621 5763
rect 11379 5732 11621 5760
rect 11379 5729 11391 5732
rect 11333 5723 11391 5729
rect 11609 5729 11621 5732
rect 11655 5729 11667 5763
rect 11609 5723 11667 5729
rect 11793 5763 11851 5769
rect 11793 5729 11805 5763
rect 11839 5760 11851 5763
rect 12066 5760 12072 5772
rect 11839 5732 12072 5760
rect 11839 5729 11851 5732
rect 11793 5723 11851 5729
rect 12066 5720 12072 5732
rect 12124 5720 12130 5772
rect 8481 5695 8539 5701
rect 8481 5692 8493 5695
rect 8128 5664 8493 5692
rect 7929 5655 7987 5661
rect 8481 5661 8493 5664
rect 8527 5692 8539 5695
rect 8662 5692 8668 5704
rect 8527 5664 8668 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 6917 5627 6975 5633
rect 6917 5624 6929 5627
rect 6564 5596 6929 5624
rect 6564 5556 6592 5596
rect 6917 5593 6929 5596
rect 6963 5593 6975 5627
rect 6917 5587 6975 5593
rect 8110 5584 8116 5636
rect 8168 5624 8174 5636
rect 8205 5627 8263 5633
rect 8205 5624 8217 5627
rect 8168 5596 8217 5624
rect 8168 5584 8174 5596
rect 8205 5593 8217 5596
rect 8251 5593 8263 5627
rect 8205 5587 8263 5593
rect 8386 5584 8392 5636
rect 8444 5584 8450 5636
rect 8496 5624 8524 5655
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 8938 5692 8944 5704
rect 8899 5664 8944 5692
rect 8938 5652 8944 5664
rect 8996 5652 9002 5704
rect 9125 5695 9183 5701
rect 9125 5661 9137 5695
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 9030 5624 9036 5636
rect 8496 5596 9036 5624
rect 9030 5584 9036 5596
rect 9088 5584 9094 5636
rect 5736 5528 6592 5556
rect 3237 5519 3295 5525
rect 7190 5516 7196 5568
rect 7248 5556 7254 5568
rect 7466 5556 7472 5568
rect 7248 5528 7472 5556
rect 7248 5516 7254 5528
rect 7466 5516 7472 5528
rect 7524 5556 7530 5568
rect 8404 5556 8432 5584
rect 7524 5528 8432 5556
rect 8665 5559 8723 5565
rect 7524 5516 7530 5528
rect 8665 5525 8677 5559
rect 8711 5556 8723 5559
rect 9140 5556 9168 5655
rect 9306 5652 9312 5704
rect 9364 5692 9370 5704
rect 9401 5695 9459 5701
rect 9401 5692 9413 5695
rect 9364 5664 9413 5692
rect 9364 5652 9370 5664
rect 9401 5661 9413 5664
rect 9447 5692 9459 5695
rect 11054 5692 11060 5704
rect 9447 5664 11060 5692
rect 9447 5661 9459 5664
rect 9401 5655 9459 5661
rect 11054 5652 11060 5664
rect 11112 5652 11118 5704
rect 11882 5692 11888 5704
rect 11843 5664 11888 5692
rect 11882 5652 11888 5664
rect 11940 5652 11946 5704
rect 12526 5692 12532 5704
rect 12487 5664 12532 5692
rect 12526 5652 12532 5664
rect 12584 5652 12590 5704
rect 10870 5584 10876 5636
rect 10928 5624 10934 5636
rect 11149 5627 11207 5633
rect 11149 5624 11161 5627
rect 10928 5596 11161 5624
rect 10928 5584 10934 5596
rect 11149 5593 11161 5596
rect 11195 5593 11207 5627
rect 12986 5624 12992 5636
rect 12947 5596 12992 5624
rect 11149 5587 11207 5593
rect 12986 5584 12992 5596
rect 13044 5584 13050 5636
rect 13081 5627 13139 5633
rect 13081 5593 13093 5627
rect 13127 5624 13139 5627
rect 13265 5627 13323 5633
rect 13265 5624 13277 5627
rect 13127 5596 13277 5624
rect 13127 5593 13139 5596
rect 13081 5587 13139 5593
rect 13265 5593 13277 5596
rect 13311 5593 13323 5627
rect 13265 5587 13323 5593
rect 10042 5556 10048 5568
rect 8711 5528 9168 5556
rect 10003 5528 10048 5556
rect 8711 5525 8723 5528
rect 8665 5519 8723 5525
rect 10042 5516 10048 5528
rect 10100 5516 10106 5568
rect 10134 5516 10140 5568
rect 10192 5556 10198 5568
rect 10192 5528 10237 5556
rect 10192 5516 10198 5528
rect 10778 5516 10784 5568
rect 10836 5556 10842 5568
rect 11057 5559 11115 5565
rect 11057 5556 11069 5559
rect 10836 5528 11069 5556
rect 10836 5516 10842 5528
rect 11057 5525 11069 5528
rect 11103 5525 11115 5559
rect 13170 5556 13176 5568
rect 13131 5528 13176 5556
rect 11057 5519 11115 5525
rect 13170 5516 13176 5528
rect 13228 5516 13234 5568
rect 1104 5466 13892 5488
rect 1104 5414 8214 5466
rect 8266 5414 8278 5466
rect 8330 5414 8342 5466
rect 8394 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 13892 5466
rect 1104 5392 13892 5414
rect 3142 5352 3148 5364
rect 3103 5324 3148 5352
rect 3142 5312 3148 5324
rect 3200 5312 3206 5364
rect 4724 5324 7328 5352
rect 2222 5244 2228 5296
rect 2280 5244 2286 5296
rect 3510 5244 3516 5296
rect 3568 5284 3574 5296
rect 3568 5256 4476 5284
rect 3568 5244 3574 5256
rect 4448 5228 4476 5256
rect 4724 5228 4752 5324
rect 7300 5296 7328 5324
rect 8662 5312 8668 5364
rect 8720 5352 8726 5364
rect 8941 5355 8999 5361
rect 8941 5352 8953 5355
rect 8720 5324 8953 5352
rect 8720 5312 8726 5324
rect 8941 5321 8953 5324
rect 8987 5321 8999 5355
rect 10134 5352 10140 5364
rect 8941 5315 8999 5321
rect 9600 5324 10140 5352
rect 5626 5284 5632 5296
rect 5539 5256 5632 5284
rect 5626 5244 5632 5256
rect 5684 5284 5690 5296
rect 6178 5284 6184 5296
rect 5684 5256 6184 5284
rect 5684 5244 5690 5256
rect 6178 5244 6184 5256
rect 6236 5244 6242 5296
rect 6546 5244 6552 5296
rect 6604 5284 6610 5296
rect 6822 5284 6828 5296
rect 6604 5256 6828 5284
rect 6604 5244 6610 5256
rect 6822 5244 6828 5256
rect 6880 5284 6886 5296
rect 7282 5284 7288 5296
rect 6880 5256 7144 5284
rect 7195 5256 7288 5284
rect 6880 5244 6886 5256
rect 2958 5176 2964 5228
rect 3016 5216 3022 5228
rect 3786 5216 3792 5228
rect 3016 5188 3792 5216
rect 3016 5176 3022 5188
rect 3786 5176 3792 5188
rect 3844 5176 3850 5228
rect 3878 5176 3884 5228
rect 3936 5216 3942 5228
rect 3936 5188 3981 5216
rect 3936 5176 3942 5188
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 4157 5219 4215 5225
rect 4157 5216 4169 5219
rect 4120 5188 4169 5216
rect 4120 5176 4126 5188
rect 4157 5185 4169 5188
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5185 4307 5219
rect 4430 5216 4436 5228
rect 4391 5188 4436 5216
rect 4249 5179 4307 5185
rect 1394 5148 1400 5160
rect 1355 5120 1400 5148
rect 1394 5108 1400 5120
rect 1452 5108 1458 5160
rect 1673 5151 1731 5157
rect 1673 5117 1685 5151
rect 1719 5148 1731 5151
rect 2406 5148 2412 5160
rect 1719 5120 2412 5148
rect 1719 5117 1731 5120
rect 1673 5111 1731 5117
rect 2406 5108 2412 5120
rect 2464 5108 2470 5160
rect 4264 5080 4292 5179
rect 4430 5176 4436 5188
rect 4488 5176 4494 5228
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5185 4583 5219
rect 4525 5179 4583 5185
rect 4618 5219 4676 5225
rect 4618 5185 4630 5219
rect 4664 5216 4676 5219
rect 4706 5216 4712 5228
rect 4664 5188 4712 5216
rect 4664 5185 4676 5188
rect 4618 5179 4676 5185
rect 4540 5148 4568 5179
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 4890 5176 4896 5228
rect 4948 5176 4954 5228
rect 5258 5216 5264 5228
rect 5171 5188 5264 5216
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5216 5503 5219
rect 5813 5219 5871 5225
rect 5813 5216 5825 5219
rect 5491 5188 5825 5216
rect 5491 5185 5503 5188
rect 5445 5179 5503 5185
rect 5813 5185 5825 5188
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 5997 5219 6055 5225
rect 5997 5185 6009 5219
rect 6043 5216 6055 5219
rect 6089 5219 6147 5225
rect 6089 5216 6101 5219
rect 6043 5188 6101 5216
rect 6043 5185 6055 5188
rect 5997 5179 6055 5185
rect 6089 5185 6101 5188
rect 6135 5216 6147 5219
rect 6641 5219 6699 5225
rect 6641 5216 6653 5219
rect 6135 5188 6653 5216
rect 6135 5185 6147 5188
rect 6089 5179 6147 5185
rect 6641 5185 6653 5188
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 4908 5148 4936 5176
rect 4540 5120 4936 5148
rect 4614 5080 4620 5092
rect 4264 5052 4620 5080
rect 4614 5040 4620 5052
rect 4672 5040 4678 5092
rect 3605 5015 3663 5021
rect 3605 4981 3617 5015
rect 3651 5012 3663 5015
rect 3694 5012 3700 5024
rect 3651 4984 3700 5012
rect 3651 4981 3663 4984
rect 3605 4975 3663 4981
rect 3694 4972 3700 4984
rect 3752 4972 3758 5024
rect 3786 4972 3792 5024
rect 3844 5012 3850 5024
rect 4065 5015 4123 5021
rect 4065 5012 4077 5015
rect 3844 4984 4077 5012
rect 3844 4972 3850 4984
rect 4065 4981 4077 4984
rect 4111 5012 4123 5015
rect 4724 5012 4752 5120
rect 4893 5083 4951 5089
rect 4893 5049 4905 5083
rect 4939 5049 4951 5083
rect 5276 5080 5304 5176
rect 5534 5148 5540 5160
rect 5495 5120 5540 5148
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 5828 5148 5856 5179
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 7116 5225 7144 5256
rect 7282 5244 7288 5256
rect 7340 5244 7346 5296
rect 7653 5287 7711 5293
rect 7653 5253 7665 5287
rect 7699 5284 7711 5287
rect 7834 5284 7840 5296
rect 7699 5256 7840 5284
rect 7699 5253 7711 5256
rect 7653 5247 7711 5253
rect 7834 5244 7840 5256
rect 7892 5244 7898 5296
rect 8570 5284 8576 5296
rect 7944 5256 8576 5284
rect 7101 5219 7159 5225
rect 6788 5188 6833 5216
rect 6788 5176 6794 5188
rect 7101 5185 7113 5219
rect 7147 5185 7159 5219
rect 7101 5179 7159 5185
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 7745 5219 7803 5225
rect 7745 5185 7757 5219
rect 7791 5216 7803 5219
rect 7944 5216 7972 5256
rect 8570 5244 8576 5256
rect 8628 5284 8634 5296
rect 9306 5284 9312 5296
rect 8628 5256 9312 5284
rect 8628 5244 8634 5256
rect 9306 5244 9312 5256
rect 9364 5244 9370 5296
rect 7791 5188 7972 5216
rect 8205 5219 8263 5225
rect 7791 5185 7803 5188
rect 7745 5179 7803 5185
rect 8205 5185 8217 5219
rect 8251 5185 8263 5219
rect 8205 5179 8263 5185
rect 8665 5219 8723 5225
rect 8665 5185 8677 5219
rect 8711 5216 8723 5219
rect 8938 5216 8944 5228
rect 8711 5188 8944 5216
rect 8711 5185 8723 5188
rect 8665 5179 8723 5185
rect 6825 5151 6883 5157
rect 5828 5120 6132 5148
rect 6104 5080 6132 5120
rect 6825 5117 6837 5151
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 6178 5080 6184 5092
rect 5276 5052 5856 5080
rect 6104 5052 6184 5080
rect 4893 5043 4951 5049
rect 4111 4984 4752 5012
rect 4908 5012 4936 5043
rect 5718 5012 5724 5024
rect 4908 4984 5724 5012
rect 4111 4981 4123 4984
rect 4065 4975 4123 4981
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 5828 5012 5856 5052
rect 6178 5040 6184 5052
rect 6236 5080 6242 5092
rect 6840 5080 6868 5111
rect 6914 5108 6920 5160
rect 6972 5148 6978 5160
rect 7484 5148 7512 5179
rect 7837 5151 7895 5157
rect 7837 5148 7849 5151
rect 6972 5120 7017 5148
rect 7484 5120 7849 5148
rect 6972 5108 6978 5120
rect 7837 5117 7849 5120
rect 7883 5148 7895 5151
rect 8220 5148 8248 5179
rect 8938 5176 8944 5188
rect 8996 5216 9002 5228
rect 9217 5219 9275 5225
rect 9217 5216 9229 5219
rect 8996 5188 9229 5216
rect 8996 5176 9002 5188
rect 9217 5185 9229 5188
rect 9263 5185 9275 5219
rect 9217 5179 9275 5185
rect 9493 5219 9551 5225
rect 9493 5185 9505 5219
rect 9539 5216 9551 5219
rect 9600 5216 9628 5324
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 10962 5352 10968 5364
rect 10923 5324 10968 5352
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 11974 5352 11980 5364
rect 11900 5324 11980 5352
rect 11514 5284 11520 5296
rect 10336 5256 11100 5284
rect 11475 5256 11520 5284
rect 10336 5225 10364 5256
rect 11072 5228 11100 5256
rect 11514 5244 11520 5256
rect 11572 5244 11578 5296
rect 11900 5293 11928 5324
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 11885 5287 11943 5293
rect 11885 5253 11897 5287
rect 11931 5253 11943 5287
rect 11885 5247 11943 5253
rect 9539 5188 9628 5216
rect 9953 5219 10011 5225
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 9953 5185 9965 5219
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 10321 5219 10379 5225
rect 10321 5185 10333 5219
rect 10367 5185 10379 5219
rect 10502 5216 10508 5228
rect 10463 5188 10508 5216
rect 10321 5179 10379 5185
rect 9582 5148 9588 5160
rect 7883 5120 9588 5148
rect 7883 5117 7895 5120
rect 7837 5111 7895 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 9968 5148 9996 5179
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5216 10655 5219
rect 10686 5216 10692 5228
rect 10643 5188 10692 5216
rect 10643 5185 10655 5188
rect 10597 5179 10655 5185
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 10778 5209 10836 5215
rect 10778 5175 10790 5209
rect 10824 5175 10836 5209
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 11333 5219 11391 5225
rect 11333 5216 11345 5219
rect 11112 5188 11345 5216
rect 11112 5176 11118 5188
rect 11333 5185 11345 5188
rect 11379 5185 11391 5219
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 11333 5179 11391 5185
rect 11440 5188 11713 5216
rect 10778 5169 10836 5175
rect 9968 5120 10732 5148
rect 10704 5092 10732 5120
rect 10796 5092 10824 5169
rect 11440 5160 11468 5188
rect 11701 5185 11713 5188
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 11241 5151 11299 5157
rect 11241 5117 11253 5151
rect 11287 5148 11299 5151
rect 11422 5148 11428 5160
rect 11287 5120 11428 5148
rect 11287 5117 11299 5120
rect 11241 5111 11299 5117
rect 11422 5108 11428 5120
rect 11480 5108 11486 5160
rect 6236 5052 6868 5080
rect 6236 5040 6242 5052
rect 7558 5040 7564 5092
rect 7616 5080 7622 5092
rect 8110 5080 8116 5092
rect 7616 5052 8116 5080
rect 7616 5040 7622 5052
rect 8110 5040 8116 5052
rect 8168 5080 8174 5092
rect 8481 5083 8539 5089
rect 8481 5080 8493 5083
rect 8168 5052 8493 5080
rect 8168 5040 8174 5052
rect 8481 5049 8493 5052
rect 8527 5049 8539 5083
rect 8481 5043 8539 5049
rect 8573 5083 8631 5089
rect 8573 5049 8585 5083
rect 8619 5080 8631 5083
rect 9677 5083 9735 5089
rect 9677 5080 9689 5083
rect 8619 5052 9689 5080
rect 8619 5049 8631 5052
rect 8573 5043 8631 5049
rect 9677 5049 9689 5052
rect 9723 5080 9735 5083
rect 10226 5080 10232 5092
rect 9723 5052 10232 5080
rect 9723 5049 9735 5052
rect 9677 5043 9735 5049
rect 6089 5015 6147 5021
rect 6089 5012 6101 5015
rect 5828 4984 6101 5012
rect 6089 4981 6101 4984
rect 6135 4981 6147 5015
rect 6454 5012 6460 5024
rect 6415 4984 6460 5012
rect 6089 4975 6147 4981
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 8386 5012 8392 5024
rect 8347 4984 8392 5012
rect 8386 4972 8392 4984
rect 8444 4972 8450 5024
rect 8496 5012 8524 5043
rect 10226 5040 10232 5052
rect 10284 5040 10290 5092
rect 10410 5080 10416 5092
rect 10371 5052 10416 5080
rect 10410 5040 10416 5052
rect 10468 5040 10474 5092
rect 10686 5040 10692 5092
rect 10744 5040 10750 5092
rect 10778 5040 10784 5092
rect 10836 5040 10842 5092
rect 11900 5080 11928 5247
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 12526 5216 12532 5228
rect 12023 5188 12532 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 12894 5216 12900 5228
rect 12855 5188 12900 5216
rect 12894 5176 12900 5188
rect 12952 5176 12958 5228
rect 10888 5052 11928 5080
rect 9585 5015 9643 5021
rect 9585 5012 9597 5015
rect 8496 4984 9597 5012
rect 9585 4981 9597 4984
rect 9631 4981 9643 5015
rect 9585 4975 9643 4981
rect 9769 5015 9827 5021
rect 9769 4981 9781 5015
rect 9815 5012 9827 5015
rect 9858 5012 9864 5024
rect 9815 4984 9864 5012
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 10134 4972 10140 5024
rect 10192 5012 10198 5024
rect 10888 5012 10916 5052
rect 12986 5040 12992 5092
rect 13044 5080 13050 5092
rect 13265 5083 13323 5089
rect 13265 5080 13277 5083
rect 13044 5052 13277 5080
rect 13044 5040 13050 5052
rect 13265 5049 13277 5052
rect 13311 5049 13323 5083
rect 13265 5043 13323 5049
rect 10192 4984 10916 5012
rect 10192 4972 10198 4984
rect 11054 4972 11060 5024
rect 11112 5012 11118 5024
rect 11149 5015 11207 5021
rect 11149 5012 11161 5015
rect 11112 4984 11161 5012
rect 11112 4972 11118 4984
rect 11149 4981 11161 4984
rect 11195 4981 11207 5015
rect 11149 4975 11207 4981
rect 1104 4922 13892 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 12214 4922
rect 12266 4870 12278 4922
rect 12330 4870 12342 4922
rect 12394 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 13892 4922
rect 1104 4848 13892 4870
rect 2222 4808 2228 4820
rect 2183 4780 2228 4808
rect 2222 4768 2228 4780
rect 2280 4768 2286 4820
rect 2406 4768 2412 4820
rect 2464 4808 2470 4820
rect 2501 4811 2559 4817
rect 2501 4808 2513 4811
rect 2464 4780 2513 4808
rect 2464 4768 2470 4780
rect 2501 4777 2513 4780
rect 2547 4777 2559 4811
rect 2501 4771 2559 4777
rect 2961 4811 3019 4817
rect 2961 4777 2973 4811
rect 3007 4808 3019 4811
rect 3510 4808 3516 4820
rect 3007 4780 3516 4808
rect 3007 4777 3019 4780
rect 2961 4771 3019 4777
rect 3510 4768 3516 4780
rect 3568 4768 3574 4820
rect 4525 4811 4583 4817
rect 4525 4777 4537 4811
rect 4571 4808 4583 4811
rect 4614 4808 4620 4820
rect 4571 4780 4620 4808
rect 4571 4777 4583 4780
rect 4525 4771 4583 4777
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 6178 4808 6184 4820
rect 6139 4780 6184 4808
rect 6178 4768 6184 4780
rect 6236 4768 6242 4820
rect 7282 4768 7288 4820
rect 7340 4808 7346 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7340 4780 7849 4808
rect 7340 4768 7346 4780
rect 7837 4777 7849 4780
rect 7883 4808 7895 4811
rect 9858 4808 9864 4820
rect 7883 4780 9864 4808
rect 7883 4777 7895 4780
rect 7837 4771 7895 4777
rect 9858 4768 9864 4780
rect 9916 4808 9922 4820
rect 10502 4808 10508 4820
rect 9916 4780 10508 4808
rect 9916 4768 9922 4780
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 10778 4808 10784 4820
rect 10739 4780 10784 4808
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 13354 4808 13360 4820
rect 13315 4780 13360 4808
rect 13354 4768 13360 4780
rect 13412 4768 13418 4820
rect 5997 4743 6055 4749
rect 5997 4740 6009 4743
rect 3988 4712 6009 4740
rect 2866 4672 2872 4684
rect 2700 4644 2872 4672
rect 2038 4604 2044 4616
rect 1951 4576 2044 4604
rect 2038 4564 2044 4576
rect 2096 4604 2102 4616
rect 2498 4604 2504 4616
rect 2096 4576 2504 4604
rect 2096 4564 2102 4576
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 2700 4613 2728 4644
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 3053 4675 3111 4681
rect 3053 4641 3065 4675
rect 3099 4672 3111 4675
rect 3142 4672 3148 4684
rect 3099 4644 3148 4672
rect 3099 4641 3111 4644
rect 3053 4635 3111 4641
rect 3142 4632 3148 4644
rect 3200 4632 3206 4684
rect 3694 4672 3700 4684
rect 3436 4644 3700 4672
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4573 2743 4607
rect 2685 4567 2743 4573
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4604 2835 4607
rect 2958 4604 2964 4616
rect 2823 4576 2964 4604
rect 2823 4573 2835 4576
rect 2777 4567 2835 4573
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 3436 4613 3464 4644
rect 3694 4632 3700 4644
rect 3752 4672 3758 4684
rect 3988 4681 4016 4712
rect 5997 4709 6009 4712
rect 6043 4709 6055 4743
rect 8754 4740 8760 4752
rect 8715 4712 8760 4740
rect 5997 4703 6055 4709
rect 8754 4700 8760 4712
rect 8812 4740 8818 4752
rect 9677 4743 9735 4749
rect 8812 4712 9628 4740
rect 8812 4700 8818 4712
rect 3973 4675 4031 4681
rect 3973 4672 3985 4675
rect 3752 4644 3985 4672
rect 3752 4632 3758 4644
rect 3973 4641 3985 4644
rect 4019 4641 4031 4675
rect 3973 4635 4031 4641
rect 4430 4632 4436 4684
rect 4488 4672 4494 4684
rect 4798 4672 4804 4684
rect 4488 4644 4804 4672
rect 4488 4632 4494 4644
rect 4798 4632 4804 4644
rect 4856 4632 4862 4684
rect 5244 4675 5302 4681
rect 5244 4641 5256 4675
rect 5290 4672 5302 4675
rect 5350 4672 5356 4684
rect 5290 4644 5356 4672
rect 5290 4641 5302 4644
rect 5244 4635 5302 4641
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 5534 4672 5540 4684
rect 5495 4644 5540 4672
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 6365 4675 6423 4681
rect 6365 4641 6377 4675
rect 6411 4672 6423 4675
rect 7009 4675 7067 4681
rect 7009 4672 7021 4675
rect 6411 4644 7021 4672
rect 6411 4641 6423 4644
rect 6365 4635 6423 4641
rect 7009 4641 7021 4644
rect 7055 4641 7067 4675
rect 8018 4672 8024 4684
rect 7009 4635 7067 4641
rect 7392 4644 8024 4672
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4573 3479 4607
rect 3421 4567 3479 4573
rect 3605 4607 3663 4613
rect 3605 4573 3617 4607
rect 3651 4604 3663 4607
rect 4062 4604 4068 4616
rect 3651 4576 4068 4604
rect 3651 4573 3663 4576
rect 3605 4567 3663 4573
rect 4062 4564 4068 4576
rect 4120 4564 4126 4616
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4604 5503 4607
rect 5626 4604 5632 4616
rect 5491 4576 5632 4604
rect 5491 4573 5503 4576
rect 5445 4567 5503 4573
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 5723 4576 6469 4604
rect 3234 4536 3240 4548
rect 3195 4508 3240 4536
rect 3234 4496 3240 4508
rect 3292 4496 3298 4548
rect 4430 4536 4436 4548
rect 4080 4508 4436 4536
rect 4080 4477 4108 4508
rect 4430 4496 4436 4508
rect 4488 4496 4494 4548
rect 4798 4536 4804 4548
rect 4759 4508 4804 4536
rect 4798 4496 4804 4508
rect 4856 4496 4862 4548
rect 4982 4536 4988 4548
rect 4943 4508 4988 4536
rect 4982 4496 4988 4508
rect 5040 4496 5046 4548
rect 5074 4496 5080 4548
rect 5132 4536 5138 4548
rect 5329 4539 5387 4545
rect 5329 4536 5341 4539
rect 5132 4508 5341 4536
rect 5132 4496 5138 4508
rect 5329 4505 5341 4508
rect 5375 4505 5387 4539
rect 5329 4499 5387 4505
rect 5534 4496 5540 4548
rect 5592 4536 5598 4548
rect 5723 4536 5751 4576
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 6553 4607 6611 4613
rect 6553 4573 6565 4607
rect 6599 4573 6611 4607
rect 6553 4567 6611 4573
rect 6641 4607 6699 4613
rect 6641 4573 6653 4607
rect 6687 4573 6699 4607
rect 6822 4604 6828 4616
rect 6783 4576 6828 4604
rect 6641 4567 6699 4573
rect 5592 4508 5751 4536
rect 5997 4539 6055 4545
rect 5592 4496 5598 4508
rect 5997 4505 6009 4539
rect 6043 4536 6055 4539
rect 6564 4536 6592 4567
rect 6043 4508 6592 4536
rect 6656 4536 6684 4567
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 7190 4604 7196 4616
rect 7151 4576 7196 4604
rect 7190 4564 7196 4576
rect 7248 4564 7254 4616
rect 7392 4613 7420 4644
rect 8018 4632 8024 4644
rect 8076 4632 8082 4684
rect 8938 4632 8944 4684
rect 8996 4672 9002 4684
rect 9033 4675 9091 4681
rect 9033 4672 9045 4675
rect 8996 4644 9045 4672
rect 8996 4632 9002 4644
rect 9033 4641 9045 4644
rect 9079 4641 9091 4675
rect 9033 4635 9091 4641
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4573 7435 4607
rect 7377 4567 7435 4573
rect 7466 4564 7472 4616
rect 7524 4604 7530 4616
rect 7745 4607 7803 4613
rect 7524 4576 7569 4604
rect 7524 4564 7530 4576
rect 7745 4573 7757 4607
rect 7791 4604 7803 4607
rect 8386 4604 8392 4616
rect 7791 4576 8392 4604
rect 7791 4573 7803 4576
rect 7745 4567 7803 4573
rect 7208 4536 7236 4564
rect 7760 4536 7788 4567
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 8570 4604 8576 4616
rect 8531 4576 8576 4604
rect 8570 4564 8576 4576
rect 8628 4564 8634 4616
rect 9306 4604 9312 4616
rect 9267 4576 9312 4604
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 9600 4604 9628 4712
rect 9677 4709 9689 4743
rect 9723 4740 9735 4743
rect 11517 4743 11575 4749
rect 9723 4712 11100 4740
rect 9723 4709 9735 4712
rect 9677 4703 9735 4709
rect 10410 4672 10416 4684
rect 10323 4644 10416 4672
rect 10410 4632 10416 4644
rect 10468 4672 10474 4684
rect 11072 4681 11100 4712
rect 11517 4709 11529 4743
rect 11563 4740 11575 4743
rect 11563 4712 12480 4740
rect 11563 4709 11575 4712
rect 11517 4703 11575 4709
rect 11057 4675 11115 4681
rect 10468 4644 10732 4672
rect 10468 4632 10474 4644
rect 9950 4604 9956 4616
rect 9600 4576 9956 4604
rect 9950 4564 9956 4576
rect 10008 4564 10014 4616
rect 10134 4604 10140 4616
rect 10095 4576 10140 4604
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 10226 4564 10232 4616
rect 10284 4604 10290 4616
rect 10321 4607 10379 4613
rect 10321 4604 10333 4607
rect 10284 4576 10333 4604
rect 10284 4564 10290 4576
rect 10321 4573 10333 4576
rect 10367 4573 10379 4607
rect 10502 4604 10508 4616
rect 10463 4576 10508 4604
rect 10321 4567 10379 4573
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4573 10655 4607
rect 10704 4604 10732 4644
rect 11057 4641 11069 4675
rect 11103 4672 11115 4675
rect 12452 4672 12480 4712
rect 13170 4700 13176 4752
rect 13228 4700 13234 4752
rect 13188 4672 13216 4700
rect 11103 4644 11744 4672
rect 11103 4641 11115 4644
rect 11057 4635 11115 4641
rect 11514 4604 11520 4616
rect 10704 4576 11520 4604
rect 10597 4567 10655 4573
rect 6656 4508 7236 4536
rect 7300 4508 7788 4536
rect 6043 4505 6055 4508
rect 5997 4499 6055 4505
rect 4065 4471 4123 4477
rect 4065 4437 4077 4471
rect 4111 4437 4123 4471
rect 4065 4431 4123 4437
rect 4157 4471 4215 4477
rect 4157 4437 4169 4471
rect 4203 4468 4215 4471
rect 4522 4468 4528 4480
rect 4203 4440 4528 4468
rect 4203 4437 4215 4440
rect 4157 4431 4215 4437
rect 4522 4428 4528 4440
rect 4580 4468 4586 4480
rect 7300 4468 7328 4508
rect 7834 4496 7840 4548
rect 7892 4536 7898 4548
rect 7892 4508 9904 4536
rect 7892 4496 7898 4508
rect 7558 4468 7564 4480
rect 4580 4440 7328 4468
rect 7519 4440 7564 4468
rect 4580 4428 4586 4440
rect 7558 4428 7564 4440
rect 7616 4428 7622 4480
rect 8662 4428 8668 4480
rect 8720 4468 8726 4480
rect 9876 4477 9904 4508
rect 10410 4496 10416 4548
rect 10468 4536 10474 4548
rect 10612 4536 10640 4567
rect 11514 4564 11520 4576
rect 11572 4564 11578 4616
rect 11716 4613 11744 4644
rect 12452 4644 13216 4672
rect 12452 4613 12480 4644
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 12437 4607 12495 4613
rect 12437 4573 12449 4607
rect 12483 4573 12495 4607
rect 12437 4567 12495 4573
rect 12621 4607 12679 4613
rect 12621 4573 12633 4607
rect 12667 4604 12679 4607
rect 12894 4604 12900 4616
rect 12667 4576 12900 4604
rect 12667 4573 12679 4576
rect 12621 4567 12679 4573
rect 12894 4564 12900 4576
rect 12952 4564 12958 4616
rect 12986 4564 12992 4616
rect 13044 4604 13050 4616
rect 13173 4607 13231 4613
rect 13173 4604 13185 4607
rect 13044 4576 13185 4604
rect 13044 4564 13050 4576
rect 13173 4573 13185 4576
rect 13219 4573 13231 4607
rect 13173 4567 13231 4573
rect 10686 4536 10692 4548
rect 10468 4508 10692 4536
rect 10468 4496 10474 4508
rect 10686 4496 10692 4508
rect 10744 4496 10750 4548
rect 11609 4539 11667 4545
rect 11609 4505 11621 4539
rect 11655 4536 11667 4539
rect 11655 4508 12434 4536
rect 11655 4505 11667 4508
rect 11609 4499 11667 4505
rect 9217 4471 9275 4477
rect 9217 4468 9229 4471
rect 8720 4440 9229 4468
rect 8720 4428 8726 4440
rect 9217 4437 9229 4440
rect 9263 4437 9275 4471
rect 9217 4431 9275 4437
rect 9861 4471 9919 4477
rect 9861 4437 9873 4471
rect 9907 4468 9919 4471
rect 10042 4468 10048 4480
rect 9907 4440 10048 4468
rect 9907 4437 9919 4440
rect 9861 4431 9919 4437
rect 10042 4428 10048 4440
rect 10100 4428 10106 4480
rect 12406 4468 12434 4508
rect 12713 4471 12771 4477
rect 12713 4468 12725 4471
rect 12406 4440 12725 4468
rect 12713 4437 12725 4440
rect 12759 4437 12771 4471
rect 12713 4431 12771 4437
rect 13081 4471 13139 4477
rect 13081 4437 13093 4471
rect 13127 4468 13139 4471
rect 13262 4468 13268 4480
rect 13127 4440 13268 4468
rect 13127 4437 13139 4440
rect 13081 4431 13139 4437
rect 13262 4428 13268 4440
rect 13320 4428 13326 4480
rect 1104 4378 13892 4400
rect 1104 4326 8214 4378
rect 8266 4326 8278 4378
rect 8330 4326 8342 4378
rect 8394 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 13892 4378
rect 1104 4304 13892 4326
rect 3510 4264 3516 4276
rect 3471 4236 3516 4264
rect 3510 4224 3516 4236
rect 3568 4224 3574 4276
rect 4982 4264 4988 4276
rect 3896 4236 4988 4264
rect 2406 4156 2412 4208
rect 2464 4156 2470 4208
rect 2958 4156 2964 4208
rect 3016 4196 3022 4208
rect 3896 4205 3924 4236
rect 4982 4224 4988 4236
rect 5040 4224 5046 4276
rect 6454 4264 6460 4276
rect 5460 4236 6460 4264
rect 3881 4199 3939 4205
rect 3881 4196 3893 4199
rect 3016 4168 3893 4196
rect 3016 4156 3022 4168
rect 3881 4165 3893 4168
rect 3927 4165 3939 4199
rect 4522 4196 4528 4208
rect 3881 4159 3939 4165
rect 4264 4168 4528 4196
rect 3234 4088 3240 4140
rect 3292 4128 3298 4140
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 3292 4100 3341 4128
rect 3292 4088 3298 4100
rect 3329 4097 3341 4100
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 3651 4131 3709 4137
rect 3651 4097 3663 4131
rect 3697 4128 3709 4131
rect 4264 4128 4292 4168
rect 4522 4156 4528 4168
rect 4580 4156 4586 4208
rect 4617 4199 4675 4205
rect 4617 4165 4629 4199
rect 4663 4196 4675 4199
rect 4706 4196 4712 4208
rect 4663 4168 4712 4196
rect 4663 4165 4675 4168
rect 4617 4159 4675 4165
rect 4706 4156 4712 4168
rect 4764 4156 4770 4208
rect 4430 4137 4436 4140
rect 4428 4128 4436 4137
rect 3697 4100 4292 4128
rect 4391 4100 4436 4128
rect 3697 4097 3709 4100
rect 3651 4091 3709 4097
rect 1394 4060 1400 4072
rect 1355 4032 1400 4060
rect 1394 4020 1400 4032
rect 1452 4020 1458 4072
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4060 1731 4063
rect 3418 4060 3424 4072
rect 1719 4032 2774 4060
rect 3379 4032 3424 4060
rect 1719 4029 1731 4032
rect 1673 4023 1731 4029
rect 2746 3992 2774 4032
rect 3418 4020 3424 4032
rect 3476 4020 3482 4072
rect 3881 3995 3939 4001
rect 3881 3992 3893 3995
rect 2746 3964 3893 3992
rect 3881 3961 3893 3964
rect 3927 3961 3939 3995
rect 3881 3955 3939 3961
rect 3145 3927 3203 3933
rect 3145 3893 3157 3927
rect 3191 3924 3203 3927
rect 3988 3924 4016 4100
rect 4428 4091 4436 4100
rect 4430 4088 4436 4091
rect 4488 4088 4494 4140
rect 4801 4131 4859 4137
rect 4801 4097 4813 4131
rect 4847 4128 4859 4131
rect 4890 4128 4896 4140
rect 4847 4100 4896 4128
rect 4847 4097 4859 4100
rect 4801 4091 4859 4097
rect 4816 3992 4844 4091
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5000 4128 5028 4224
rect 5460 4205 5488 4236
rect 5445 4199 5503 4205
rect 5445 4165 5457 4199
rect 5491 4165 5503 4199
rect 5445 4159 5503 4165
rect 5537 4199 5595 4205
rect 5537 4165 5549 4199
rect 5583 4196 5595 4199
rect 6089 4199 6147 4205
rect 6089 4196 6101 4199
rect 5583 4168 6101 4196
rect 5583 4165 5595 4168
rect 5537 4159 5595 4165
rect 6089 4165 6101 4168
rect 6135 4165 6147 4199
rect 6089 4159 6147 4165
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 5000 4100 5181 4128
rect 5169 4097 5181 4100
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 5317 4131 5375 4137
rect 5317 4097 5329 4131
rect 5363 4128 5375 4131
rect 5675 4131 5733 4137
rect 5363 4097 5396 4128
rect 5317 4091 5396 4097
rect 5675 4097 5687 4131
rect 5721 4128 5733 4131
rect 5902 4128 5908 4140
rect 5721 4100 5908 4128
rect 5721 4097 5733 4100
rect 5675 4091 5733 4097
rect 5368 4060 5396 4091
rect 5902 4088 5908 4100
rect 5960 4088 5966 4140
rect 6181 4131 6239 4137
rect 6181 4097 6193 4131
rect 6227 4128 6239 4131
rect 6288 4128 6316 4236
rect 6454 4224 6460 4236
rect 6512 4224 6518 4276
rect 6914 4224 6920 4276
rect 6972 4264 6978 4276
rect 11149 4267 11207 4273
rect 11149 4264 11161 4267
rect 6972 4236 11161 4264
rect 6972 4224 6978 4236
rect 11149 4233 11161 4236
rect 11195 4264 11207 4267
rect 11790 4264 11796 4276
rect 11195 4236 11796 4264
rect 11195 4233 11207 4236
rect 11149 4227 11207 4233
rect 11790 4224 11796 4236
rect 11848 4224 11854 4276
rect 8018 4156 8024 4208
rect 8076 4196 8082 4208
rect 9306 4196 9312 4208
rect 8076 4168 9312 4196
rect 8076 4156 8082 4168
rect 9306 4156 9312 4168
rect 9364 4196 9370 4208
rect 9364 4168 9996 4196
rect 9364 4156 9370 4168
rect 9968 4140 9996 4168
rect 10134 4156 10140 4208
rect 10192 4196 10198 4208
rect 10505 4199 10563 4205
rect 10192 4168 10456 4196
rect 10192 4156 10198 4168
rect 6227 4100 6316 4128
rect 6227 4097 6239 4100
rect 6181 4091 6239 4097
rect 6362 4088 6368 4140
rect 6420 4128 6426 4140
rect 6641 4131 6699 4137
rect 6420 4100 6465 4128
rect 6420 4088 6426 4100
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 7006 4128 7012 4140
rect 6687 4100 7012 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 7006 4088 7012 4100
rect 7064 4128 7070 4140
rect 7374 4128 7380 4140
rect 7064 4100 7380 4128
rect 7064 4088 7070 4100
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 7834 4128 7840 4140
rect 7795 4100 7840 4128
rect 7834 4088 7840 4100
rect 7892 4088 7898 4140
rect 9214 4128 9220 4140
rect 9175 4100 9220 4128
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 9401 4131 9459 4137
rect 9401 4097 9413 4131
rect 9447 4097 9459 4131
rect 9950 4128 9956 4140
rect 9863 4100 9956 4128
rect 9401 4091 9459 4097
rect 6457 4063 6515 4069
rect 6457 4060 6469 4063
rect 5368 4032 6469 4060
rect 6457 4029 6469 4032
rect 6503 4029 6515 4063
rect 6457 4023 6515 4029
rect 8205 4063 8263 4069
rect 8205 4029 8217 4063
rect 8251 4060 8263 4063
rect 8294 4060 8300 4072
rect 8251 4032 8300 4060
rect 8251 4029 8263 4032
rect 8205 4023 8263 4029
rect 8294 4020 8300 4032
rect 8352 4060 8358 4072
rect 9122 4060 9128 4072
rect 8352 4032 9128 4060
rect 8352 4020 8358 4032
rect 9122 4020 9128 4032
rect 9180 4020 9186 4072
rect 6822 3992 6828 4004
rect 4816 3964 6828 3992
rect 6822 3952 6828 3964
rect 6880 3952 6886 4004
rect 8846 3952 8852 4004
rect 8904 3992 8910 4004
rect 9416 3992 9444 4091
rect 9950 4088 9956 4100
rect 10008 4088 10014 4140
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 10100 4100 10145 4128
rect 10100 4088 10106 4100
rect 10226 4088 10232 4140
rect 10284 4128 10290 4140
rect 10428 4137 10456 4168
rect 10505 4165 10517 4199
rect 10551 4165 10563 4199
rect 10686 4196 10692 4208
rect 10647 4168 10692 4196
rect 10505 4159 10563 4165
rect 10413 4131 10471 4137
rect 10284 4100 10377 4128
rect 10284 4088 10290 4100
rect 10413 4097 10425 4131
rect 10459 4097 10471 4131
rect 10413 4091 10471 4097
rect 10244 4060 10272 4088
rect 10520 4060 10548 4159
rect 10686 4156 10692 4168
rect 10744 4196 10750 4208
rect 11054 4196 11060 4208
rect 10744 4168 11060 4196
rect 10744 4156 10750 4168
rect 11054 4156 11060 4168
rect 11112 4156 11118 4208
rect 11514 4156 11520 4208
rect 11572 4156 11578 4208
rect 11241 4131 11299 4137
rect 11241 4097 11253 4131
rect 11287 4128 11299 4131
rect 11532 4128 11560 4156
rect 11287 4100 11560 4128
rect 12161 4131 12219 4137
rect 11287 4097 11299 4100
rect 11241 4091 11299 4097
rect 12161 4097 12173 4131
rect 12207 4128 12219 4131
rect 13262 4128 13268 4140
rect 12207 4100 13124 4128
rect 13223 4100 13268 4128
rect 12207 4097 12219 4100
rect 12161 4091 12219 4097
rect 10244 4032 10548 4060
rect 10428 4004 10456 4032
rect 8904 3964 9444 3992
rect 9585 3995 9643 4001
rect 8904 3952 8910 3964
rect 9585 3961 9597 3995
rect 9631 3992 9643 3995
rect 10137 3995 10195 4001
rect 10137 3992 10149 3995
rect 9631 3964 10149 3992
rect 9631 3961 9643 3964
rect 9585 3955 9643 3961
rect 10137 3961 10149 3964
rect 10183 3961 10195 3995
rect 10137 3955 10195 3961
rect 3191 3896 4016 3924
rect 3191 3893 3203 3896
rect 3145 3887 3203 3893
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 4249 3927 4307 3933
rect 4249 3924 4261 3927
rect 4120 3896 4261 3924
rect 4120 3884 4126 3896
rect 4249 3893 4261 3896
rect 4295 3924 4307 3927
rect 5534 3924 5540 3936
rect 4295 3896 5540 3924
rect 4295 3893 4307 3896
rect 4249 3887 4307 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 5810 3924 5816 3936
rect 5771 3896 5816 3924
rect 5810 3884 5816 3896
rect 5868 3884 5874 3936
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 8570 3924 8576 3936
rect 7524 3896 8576 3924
rect 7524 3884 7530 3896
rect 8570 3884 8576 3896
rect 8628 3884 8634 3936
rect 8662 3884 8668 3936
rect 8720 3924 8726 3936
rect 8757 3927 8815 3933
rect 8757 3924 8769 3927
rect 8720 3896 8769 3924
rect 8720 3884 8726 3896
rect 8757 3893 8769 3896
rect 8803 3893 8815 3927
rect 8757 3887 8815 3893
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 9033 3927 9091 3933
rect 9033 3924 9045 3927
rect 8996 3896 9045 3924
rect 8996 3884 9002 3896
rect 9033 3893 9045 3896
rect 9079 3893 9091 3927
rect 9033 3887 9091 3893
rect 9769 3927 9827 3933
rect 9769 3893 9781 3927
rect 9815 3924 9827 3927
rect 9858 3924 9864 3936
rect 9815 3896 9864 3924
rect 9815 3893 9827 3896
rect 9769 3887 9827 3893
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 10152 3924 10180 3955
rect 10410 3952 10416 4004
rect 10468 3952 10474 4004
rect 10778 3992 10784 4004
rect 10691 3964 10784 3992
rect 10704 3933 10732 3964
rect 10778 3952 10784 3964
rect 10836 3992 10842 4004
rect 11256 3992 11284 4091
rect 11514 4020 11520 4072
rect 11572 4060 11578 4072
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 11572 4032 11621 4060
rect 11572 4020 11578 4032
rect 11609 4029 11621 4032
rect 11655 4029 11667 4063
rect 11609 4023 11667 4029
rect 11974 4020 11980 4072
rect 12032 4060 12038 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 12032 4032 12449 4060
rect 12032 4020 12038 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12986 4060 12992 4072
rect 12947 4032 12992 4060
rect 12437 4023 12495 4029
rect 12986 4020 12992 4032
rect 13044 4020 13050 4072
rect 10836 3964 11284 3992
rect 10836 3952 10842 3964
rect 11698 3952 11704 4004
rect 11756 3992 11762 4004
rect 12069 3995 12127 4001
rect 12069 3992 12081 3995
rect 11756 3964 12081 3992
rect 11756 3952 11762 3964
rect 12069 3961 12081 3964
rect 12115 3961 12127 3995
rect 12894 3992 12900 4004
rect 12855 3964 12900 3992
rect 12069 3955 12127 3961
rect 12894 3952 12900 3964
rect 12952 3952 12958 4004
rect 13096 4001 13124 4100
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 13081 3995 13139 4001
rect 13081 3961 13093 3995
rect 13127 3961 13139 3995
rect 13081 3955 13139 3961
rect 10689 3927 10747 3933
rect 10689 3924 10701 3927
rect 10152 3896 10701 3924
rect 10689 3893 10701 3896
rect 10735 3893 10747 3927
rect 10689 3887 10747 3893
rect 10873 3927 10931 3933
rect 10873 3893 10885 3927
rect 10919 3924 10931 3927
rect 11054 3924 11060 3936
rect 10919 3896 11060 3924
rect 10919 3893 10931 3896
rect 10873 3887 10931 3893
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11882 3884 11888 3936
rect 11940 3924 11946 3936
rect 12253 3927 12311 3933
rect 12253 3924 12265 3927
rect 11940 3896 12265 3924
rect 11940 3884 11946 3896
rect 12253 3893 12265 3896
rect 12299 3893 12311 3927
rect 12253 3887 12311 3893
rect 13541 3927 13599 3933
rect 13541 3893 13553 3927
rect 13587 3924 13599 3927
rect 14001 3927 14059 3933
rect 14001 3924 14013 3927
rect 13587 3896 14013 3924
rect 13587 3893 13599 3896
rect 13541 3887 13599 3893
rect 14001 3893 14013 3896
rect 14047 3893 14059 3927
rect 14001 3887 14059 3893
rect 1104 3834 13892 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 12214 3834
rect 12266 3782 12278 3834
rect 12330 3782 12342 3834
rect 12394 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 13892 3834
rect 1104 3760 13892 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 2406 3720 2412 3732
rect 2367 3692 2412 3720
rect 2406 3680 2412 3692
rect 2464 3680 2470 3732
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 3053 3723 3111 3729
rect 3053 3720 3065 3723
rect 3016 3692 3065 3720
rect 3016 3680 3022 3692
rect 3053 3689 3065 3692
rect 3099 3689 3111 3723
rect 3053 3683 3111 3689
rect 3329 3723 3387 3729
rect 3329 3689 3341 3723
rect 3375 3720 3387 3723
rect 3418 3720 3424 3732
rect 3375 3692 3424 3720
rect 3375 3689 3387 3692
rect 3329 3683 3387 3689
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 5902 3720 5908 3732
rect 5815 3692 5908 3720
rect 5902 3680 5908 3692
rect 5960 3720 5966 3732
rect 6362 3720 6368 3732
rect 5960 3692 6368 3720
rect 5960 3680 5966 3692
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 7650 3680 7656 3732
rect 7708 3720 7714 3732
rect 9398 3720 9404 3732
rect 7708 3692 8524 3720
rect 9359 3692 9404 3720
rect 7708 3680 7714 3692
rect 5166 3652 5172 3664
rect 5127 3624 5172 3652
rect 5166 3612 5172 3624
rect 5224 3612 5230 3664
rect 5994 3612 6000 3664
rect 6052 3652 6058 3664
rect 7469 3655 7527 3661
rect 6052 3624 7420 3652
rect 6052 3612 6058 3624
rect 4614 3544 4620 3596
rect 4672 3584 4678 3596
rect 6365 3587 6423 3593
rect 6365 3584 6377 3587
rect 4672 3556 6377 3584
rect 4672 3544 4678 3556
rect 6365 3553 6377 3556
rect 6411 3553 6423 3587
rect 7006 3584 7012 3596
rect 6967 3556 7012 3584
rect 6365 3547 6423 3553
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 7392 3584 7420 3624
rect 7469 3621 7481 3655
rect 7515 3652 7527 3655
rect 8294 3652 8300 3664
rect 7515 3624 8300 3652
rect 7515 3621 7527 3624
rect 7469 3615 7527 3621
rect 8294 3612 8300 3624
rect 8352 3612 8358 3664
rect 7392 3556 8294 3584
rect 1578 3476 1584 3528
rect 1636 3516 1642 3528
rect 1765 3519 1823 3525
rect 1765 3516 1777 3519
rect 1636 3488 1777 3516
rect 1636 3476 1642 3488
rect 1765 3485 1777 3488
rect 1811 3485 1823 3519
rect 1765 3479 1823 3485
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3516 2283 3519
rect 2498 3516 2504 3528
rect 2271 3488 2504 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 2498 3476 2504 3488
rect 2556 3476 2562 3528
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3516 3203 3519
rect 3510 3516 3516 3528
rect 3191 3488 3516 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 4062 3516 4068 3528
rect 3651 3488 4068 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 5074 3476 5080 3528
rect 5132 3516 5138 3528
rect 5169 3519 5227 3525
rect 5169 3516 5181 3519
rect 5132 3488 5181 3516
rect 5132 3476 5138 3488
rect 5169 3485 5181 3488
rect 5215 3485 5227 3519
rect 5169 3479 5227 3485
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3485 5411 3519
rect 5353 3479 5411 3485
rect 5537 3519 5595 3525
rect 5537 3485 5549 3519
rect 5583 3516 5595 3519
rect 5810 3516 5816 3528
rect 5583 3488 5816 3516
rect 5583 3485 5595 3488
rect 5537 3479 5595 3485
rect 3421 3451 3479 3457
rect 3421 3417 3433 3451
rect 3467 3448 3479 3451
rect 3694 3448 3700 3460
rect 3467 3420 3700 3448
rect 3467 3417 3479 3420
rect 3421 3411 3479 3417
rect 3694 3408 3700 3420
rect 3752 3408 3758 3460
rect 5368 3448 5396 3479
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 6089 3519 6147 3525
rect 6089 3485 6101 3519
rect 6135 3485 6147 3519
rect 6089 3479 6147 3485
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3485 6239 3519
rect 6181 3479 6239 3485
rect 6457 3519 6515 3525
rect 6457 3485 6469 3519
rect 6503 3516 6515 3519
rect 6638 3516 6644 3528
rect 6503 3488 6644 3516
rect 6503 3485 6515 3488
rect 6457 3479 6515 3485
rect 6104 3448 6132 3479
rect 5368 3420 6132 3448
rect 6196 3448 6224 3479
rect 6638 3476 6644 3488
rect 6696 3516 6702 3528
rect 7466 3516 7472 3528
rect 6696 3488 7472 3516
rect 6696 3476 6702 3488
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 7834 3516 7840 3528
rect 7795 3488 7840 3516
rect 7834 3476 7840 3488
rect 7892 3476 7898 3528
rect 8266 3516 8294 3556
rect 8386 3516 8392 3528
rect 8266 3488 8392 3516
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 6822 3448 6828 3460
rect 6196 3420 6828 3448
rect 6104 3380 6132 3420
rect 6822 3408 6828 3420
rect 6880 3408 6886 3460
rect 7561 3451 7619 3457
rect 7561 3417 7573 3451
rect 7607 3448 7619 3451
rect 8021 3451 8079 3457
rect 8021 3448 8033 3451
rect 7607 3420 8033 3448
rect 7607 3417 7619 3420
rect 7561 3411 7619 3417
rect 8021 3417 8033 3420
rect 8067 3417 8079 3451
rect 8021 3411 8079 3417
rect 8496 3448 8524 3692
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 9493 3655 9551 3661
rect 9493 3652 9505 3655
rect 9324 3624 9505 3652
rect 9324 3584 9352 3624
rect 9493 3621 9505 3624
rect 9539 3621 9551 3655
rect 9493 3615 9551 3621
rect 9585 3655 9643 3661
rect 9585 3621 9597 3655
rect 9631 3652 9643 3655
rect 9950 3652 9956 3664
rect 9631 3624 9956 3652
rect 9631 3621 9643 3624
rect 9585 3615 9643 3621
rect 9950 3612 9956 3624
rect 10008 3612 10014 3664
rect 10502 3612 10508 3664
rect 10560 3652 10566 3664
rect 10597 3655 10655 3661
rect 10597 3652 10609 3655
rect 10560 3624 10609 3652
rect 10560 3612 10566 3624
rect 10597 3621 10609 3624
rect 10643 3652 10655 3655
rect 10962 3652 10968 3664
rect 10643 3624 10968 3652
rect 10643 3621 10655 3624
rect 10597 3615 10655 3621
rect 10962 3612 10968 3624
rect 11020 3612 11026 3664
rect 12894 3612 12900 3664
rect 12952 3652 12958 3664
rect 13265 3655 13323 3661
rect 13265 3652 13277 3655
rect 12952 3624 13277 3652
rect 12952 3612 12958 3624
rect 13265 3621 13277 3624
rect 13311 3621 13323 3655
rect 13265 3615 13323 3621
rect 8772 3556 9352 3584
rect 9600 3556 10456 3584
rect 8772 3528 8800 3556
rect 8570 3476 8576 3528
rect 8628 3516 8634 3528
rect 8754 3516 8760 3528
rect 8628 3488 8760 3516
rect 8628 3476 8634 3488
rect 8754 3476 8760 3488
rect 8812 3476 8818 3528
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 9309 3519 9367 3525
rect 9309 3516 9321 3519
rect 9088 3488 9321 3516
rect 9088 3476 9094 3488
rect 9309 3485 9321 3488
rect 9355 3516 9367 3519
rect 9600 3516 9628 3556
rect 10428 3525 10456 3556
rect 9355 3488 9628 3516
rect 9719 3522 9777 3525
rect 9719 3519 9772 3522
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9719 3485 9731 3519
rect 9765 3485 9772 3519
rect 9719 3479 9772 3485
rect 9766 3470 9772 3479
rect 9824 3470 9830 3522
rect 10413 3519 10471 3525
rect 10413 3485 10425 3519
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3485 10563 3519
rect 10505 3479 10563 3485
rect 10689 3519 10747 3525
rect 10689 3485 10701 3519
rect 10735 3485 10747 3519
rect 10689 3479 10747 3485
rect 10965 3519 11023 3525
rect 10965 3485 10977 3519
rect 11011 3516 11023 3519
rect 11514 3516 11520 3528
rect 11011 3488 11520 3516
rect 11011 3485 11023 3488
rect 10965 3479 11023 3485
rect 10520 3448 10548 3479
rect 8496 3420 9444 3448
rect 7466 3380 7472 3392
rect 6104 3352 7472 3380
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 7650 3380 7656 3392
rect 7611 3352 7656 3380
rect 7650 3340 7656 3352
rect 7708 3340 7714 3392
rect 7926 3380 7932 3392
rect 7887 3352 7932 3380
rect 7926 3340 7932 3352
rect 7984 3340 7990 3392
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 8496 3389 8524 3420
rect 9416 3392 9444 3420
rect 9876 3420 10548 3448
rect 10704 3448 10732 3479
rect 11514 3476 11520 3488
rect 11572 3476 11578 3528
rect 11974 3516 11980 3528
rect 11935 3488 11980 3516
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 12897 3519 12955 3525
rect 12897 3485 12909 3519
rect 12943 3516 12955 3519
rect 13262 3516 13268 3528
rect 12943 3488 13268 3516
rect 12943 3485 12955 3488
rect 12897 3479 12955 3485
rect 11054 3448 11060 3460
rect 10704 3420 11060 3448
rect 8297 3383 8355 3389
rect 8297 3380 8309 3383
rect 8168 3352 8309 3380
rect 8168 3340 8174 3352
rect 8297 3349 8309 3352
rect 8343 3349 8355 3383
rect 8297 3343 8355 3349
rect 8481 3383 8539 3389
rect 8481 3349 8493 3383
rect 8527 3349 8539 3383
rect 8481 3343 8539 3349
rect 8573 3383 8631 3389
rect 8573 3349 8585 3383
rect 8619 3380 8631 3383
rect 8846 3380 8852 3392
rect 8619 3352 8852 3380
rect 8619 3349 8631 3352
rect 8573 3343 8631 3349
rect 8846 3340 8852 3352
rect 8904 3340 8910 3392
rect 8938 3340 8944 3392
rect 8996 3380 9002 3392
rect 8996 3352 9041 3380
rect 8996 3340 9002 3352
rect 9398 3340 9404 3392
rect 9456 3380 9462 3392
rect 9876 3380 9904 3420
rect 11054 3408 11060 3420
rect 11112 3448 11118 3460
rect 11422 3448 11428 3460
rect 11112 3420 11428 3448
rect 11112 3408 11118 3420
rect 11422 3408 11428 3420
rect 11480 3408 11486 3460
rect 11698 3448 11704 3460
rect 11659 3420 11704 3448
rect 11698 3408 11704 3420
rect 11756 3408 11762 3460
rect 11885 3451 11943 3457
rect 11885 3417 11897 3451
rect 11931 3448 11943 3451
rect 12912 3448 12940 3479
rect 13262 3476 13268 3488
rect 13320 3476 13326 3528
rect 11931 3420 12940 3448
rect 11931 3417 11943 3420
rect 11885 3411 11943 3417
rect 9456 3352 9904 3380
rect 9953 3383 10011 3389
rect 9456 3340 9462 3352
rect 9953 3349 9965 3383
rect 9999 3380 10011 3383
rect 10042 3380 10048 3392
rect 9999 3352 10048 3380
rect 9999 3349 10011 3352
rect 9953 3343 10011 3349
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 10226 3380 10232 3392
rect 10187 3352 10232 3380
rect 10226 3340 10232 3352
rect 10284 3340 10290 3392
rect 1104 3290 13892 3312
rect 1104 3238 8214 3290
rect 8266 3238 8278 3290
rect 8330 3238 8342 3290
rect 8394 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 13892 3290
rect 1104 3216 13892 3238
rect 2869 3179 2927 3185
rect 2869 3145 2881 3179
rect 2915 3176 2927 3179
rect 3326 3176 3332 3188
rect 2915 3148 3332 3176
rect 2915 3145 2927 3148
rect 2869 3139 2927 3145
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 4798 3176 4804 3188
rect 3896 3148 4804 3176
rect 3896 3117 3924 3148
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 5350 3176 5356 3188
rect 5311 3148 5356 3176
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 7006 3176 7012 3188
rect 6840 3148 7012 3176
rect 3513 3111 3571 3117
rect 3513 3108 3525 3111
rect 3022 3080 3525 3108
rect 2498 3040 2504 3052
rect 2459 3012 2504 3040
rect 2498 3000 2504 3012
rect 2556 3000 2562 3052
rect 2866 3000 2872 3052
rect 2924 3040 2930 3052
rect 3022 3049 3050 3080
rect 3513 3077 3525 3080
rect 3559 3077 3571 3111
rect 3513 3071 3571 3077
rect 3881 3111 3939 3117
rect 3881 3077 3893 3111
rect 3927 3077 3939 3111
rect 3881 3071 3939 3077
rect 4614 3068 4620 3120
rect 4672 3068 4678 3120
rect 3007 3043 3065 3049
rect 3007 3040 3019 3043
rect 2924 3012 3019 3040
rect 2924 3000 2930 3012
rect 3007 3009 3019 3012
rect 3053 3009 3065 3043
rect 3007 3003 3065 3009
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3009 3203 3043
rect 5810 3040 5816 3052
rect 5771 3012 5816 3040
rect 3145 3003 3203 3009
rect 3160 2972 3188 3003
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 6840 3049 6868 3148
rect 7006 3136 7012 3148
rect 7064 3176 7070 3188
rect 8021 3179 8079 3185
rect 8021 3176 8033 3179
rect 7064 3148 8033 3176
rect 7064 3136 7070 3148
rect 8021 3145 8033 3148
rect 8067 3145 8079 3179
rect 8021 3139 8079 3145
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8389 3179 8447 3185
rect 8389 3176 8401 3179
rect 8168 3148 8401 3176
rect 8168 3136 8174 3148
rect 8389 3145 8401 3148
rect 8435 3145 8447 3179
rect 8389 3139 8447 3145
rect 8481 3179 8539 3185
rect 8481 3145 8493 3179
rect 8527 3176 8539 3179
rect 9582 3176 9588 3188
rect 8527 3148 9588 3176
rect 8527 3145 8539 3148
rect 8481 3139 8539 3145
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 9861 3179 9919 3185
rect 9861 3145 9873 3179
rect 9907 3176 9919 3179
rect 10226 3176 10232 3188
rect 9907 3148 10232 3176
rect 9907 3145 9919 3148
rect 9861 3139 9919 3145
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 11241 3179 11299 3185
rect 11241 3145 11253 3179
rect 11287 3176 11299 3179
rect 11885 3179 11943 3185
rect 11885 3176 11897 3179
rect 11287 3148 11897 3176
rect 11287 3145 11299 3148
rect 11241 3139 11299 3145
rect 11885 3145 11897 3148
rect 11931 3145 11943 3179
rect 11885 3139 11943 3145
rect 11974 3136 11980 3188
rect 12032 3176 12038 3188
rect 12529 3179 12587 3185
rect 12529 3176 12541 3179
rect 12032 3148 12541 3176
rect 12032 3136 12038 3148
rect 12529 3145 12541 3148
rect 12575 3145 12587 3179
rect 12529 3139 12587 3145
rect 12986 3136 12992 3188
rect 13044 3176 13050 3188
rect 13449 3179 13507 3185
rect 13449 3176 13461 3179
rect 13044 3148 13461 3176
rect 13044 3136 13050 3148
rect 13449 3145 13461 3148
rect 13495 3145 13507 3179
rect 13449 3139 13507 3145
rect 7466 3068 7472 3120
rect 7524 3108 7530 3120
rect 7561 3111 7619 3117
rect 7561 3108 7573 3111
rect 7524 3080 7573 3108
rect 7524 3068 7530 3080
rect 7561 3077 7573 3080
rect 7607 3108 7619 3111
rect 7926 3108 7932 3120
rect 7607 3080 7932 3108
rect 7607 3077 7619 3080
rect 7561 3071 7619 3077
rect 7926 3068 7932 3080
rect 7984 3068 7990 3120
rect 9033 3111 9091 3117
rect 9033 3077 9045 3111
rect 9079 3108 9091 3111
rect 9079 3080 11192 3108
rect 9079 3077 9091 3080
rect 9033 3071 9091 3077
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3040 7803 3043
rect 7834 3040 7840 3052
rect 7791 3012 7840 3040
rect 7791 3009 7803 3012
rect 7745 3003 7803 3009
rect 7834 3000 7840 3012
rect 7892 3040 7898 3052
rect 8110 3040 8116 3052
rect 7892 3012 8116 3040
rect 7892 3000 7898 3012
rect 8110 3000 8116 3012
rect 8168 3000 8174 3052
rect 9214 3040 9220 3052
rect 9175 3012 9220 3040
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 9398 3000 9404 3052
rect 9456 3040 9462 3052
rect 9456 3012 10364 3040
rect 9456 3000 9462 3012
rect 3418 2972 3424 2984
rect 3160 2944 3424 2972
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 3605 2975 3663 2981
rect 3605 2941 3617 2975
rect 3651 2972 3663 2975
rect 5258 2972 5264 2984
rect 3651 2944 5264 2972
rect 3651 2941 3663 2944
rect 3605 2935 3663 2941
rect 1578 2864 1584 2916
rect 1636 2904 1642 2916
rect 3620 2904 3648 2935
rect 5258 2932 5264 2944
rect 5316 2932 5322 2984
rect 7929 2975 7987 2981
rect 7929 2941 7941 2975
rect 7975 2972 7987 2975
rect 8573 2975 8631 2981
rect 8573 2972 8585 2975
rect 7975 2944 8585 2972
rect 7975 2941 7987 2944
rect 7929 2935 7987 2941
rect 8573 2941 8585 2944
rect 8619 2972 8631 2975
rect 8938 2972 8944 2984
rect 8619 2944 8944 2972
rect 8619 2941 8631 2944
rect 8573 2935 8631 2941
rect 8938 2932 8944 2944
rect 8996 2972 9002 2984
rect 9585 2975 9643 2981
rect 9585 2972 9597 2975
rect 8996 2944 9597 2972
rect 8996 2932 9002 2944
rect 9585 2941 9597 2944
rect 9631 2972 9643 2975
rect 9674 2972 9680 2984
rect 9631 2944 9680 2972
rect 9631 2941 9643 2944
rect 9585 2935 9643 2941
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 9769 2975 9827 2981
rect 9769 2941 9781 2975
rect 9815 2941 9827 2975
rect 10336 2972 10364 3012
rect 10410 3000 10416 3052
rect 10468 3040 10474 3052
rect 10597 3043 10655 3049
rect 10597 3040 10609 3043
rect 10468 3012 10609 3040
rect 10468 3000 10474 3012
rect 10597 3009 10609 3012
rect 10643 3009 10655 3043
rect 10597 3003 10655 3009
rect 10686 3000 10692 3052
rect 10744 3040 10750 3052
rect 10873 3043 10931 3049
rect 10744 3012 10789 3040
rect 10744 3000 10750 3012
rect 10873 3009 10885 3043
rect 10919 3009 10931 3043
rect 11054 3040 11060 3052
rect 11015 3012 11060 3040
rect 10873 3003 10931 3009
rect 10888 2972 10916 3003
rect 11054 3000 11060 3012
rect 11112 3000 11118 3052
rect 11164 3040 11192 3080
rect 11698 3068 11704 3120
rect 11756 3108 11762 3120
rect 13357 3111 13415 3117
rect 13357 3108 13369 3111
rect 11756 3080 13369 3108
rect 11756 3068 11762 3080
rect 13357 3077 13369 3080
rect 13403 3077 13415 3111
rect 13357 3071 13415 3077
rect 12897 3043 12955 3049
rect 12897 3040 12909 3043
rect 11164 3012 12909 3040
rect 12897 3009 12909 3012
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 12989 3043 13047 3049
rect 12989 3009 13001 3043
rect 13035 3040 13047 3043
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 13035 3012 14013 3040
rect 13035 3009 13047 3012
rect 12989 3003 13047 3009
rect 14001 3009 14013 3012
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 11882 2972 11888 2984
rect 10336 2944 10548 2972
rect 9769 2935 9827 2941
rect 1636 2876 3648 2904
rect 1636 2864 1642 2876
rect 4982 2864 4988 2916
rect 5040 2904 5046 2916
rect 8849 2907 8907 2913
rect 8849 2904 8861 2907
rect 5040 2876 8861 2904
rect 5040 2864 5046 2876
rect 8849 2873 8861 2876
rect 8895 2904 8907 2907
rect 9784 2904 9812 2935
rect 10520 2916 10548 2944
rect 10704 2944 10916 2972
rect 11164 2944 11888 2972
rect 8895 2876 9812 2904
rect 8895 2873 8907 2876
rect 8849 2867 8907 2873
rect 9950 2864 9956 2916
rect 10008 2904 10014 2916
rect 10413 2907 10471 2913
rect 10413 2904 10425 2907
rect 10008 2876 10425 2904
rect 10008 2864 10014 2876
rect 10413 2873 10425 2876
rect 10459 2873 10471 2907
rect 10413 2867 10471 2873
rect 10502 2864 10508 2916
rect 10560 2904 10566 2916
rect 10704 2904 10732 2944
rect 10560 2876 10732 2904
rect 10781 2907 10839 2913
rect 10560 2864 10566 2876
rect 10781 2873 10793 2907
rect 10827 2904 10839 2907
rect 10962 2904 10968 2916
rect 10827 2876 10968 2904
rect 10827 2873 10839 2876
rect 10781 2867 10839 2873
rect 10962 2864 10968 2876
rect 11020 2864 11026 2916
rect 11054 2864 11060 2916
rect 11112 2904 11118 2916
rect 11164 2904 11192 2944
rect 11882 2932 11888 2944
rect 11940 2972 11946 2984
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11940 2944 11989 2972
rect 11940 2932 11946 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 12066 2932 12072 2984
rect 12124 2972 12130 2984
rect 13081 2975 13139 2981
rect 13081 2972 13093 2975
rect 12124 2944 13093 2972
rect 12124 2932 12130 2944
rect 13081 2941 13093 2944
rect 13127 2941 13139 2975
rect 13081 2935 13139 2941
rect 11514 2904 11520 2916
rect 11112 2876 11192 2904
rect 11475 2876 11520 2904
rect 11112 2864 11118 2876
rect 11514 2864 11520 2876
rect 11572 2864 11578 2916
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 2685 2839 2743 2845
rect 2685 2836 2697 2839
rect 2648 2808 2697 2836
rect 2648 2796 2654 2808
rect 2685 2805 2697 2808
rect 2731 2805 2743 2839
rect 2685 2799 2743 2805
rect 5902 2796 5908 2848
rect 5960 2836 5966 2848
rect 5997 2839 6055 2845
rect 5997 2836 6009 2839
rect 5960 2808 6009 2836
rect 5960 2796 5966 2808
rect 5997 2805 6009 2808
rect 6043 2805 6055 2839
rect 5997 2799 6055 2805
rect 6178 2796 6184 2848
rect 6236 2836 6242 2848
rect 6365 2839 6423 2845
rect 6365 2836 6377 2839
rect 6236 2808 6377 2836
rect 6236 2796 6242 2808
rect 6365 2805 6377 2808
rect 6411 2836 6423 2839
rect 7929 2839 7987 2845
rect 7929 2836 7941 2839
rect 6411 2808 7941 2836
rect 6411 2805 6423 2808
rect 6365 2799 6423 2805
rect 7929 2805 7941 2808
rect 7975 2805 7987 2839
rect 7929 2799 7987 2805
rect 10229 2839 10287 2845
rect 10229 2805 10241 2839
rect 10275 2836 10287 2839
rect 10594 2836 10600 2848
rect 10275 2808 10600 2836
rect 10275 2805 10287 2808
rect 10229 2799 10287 2805
rect 10594 2796 10600 2808
rect 10652 2796 10658 2848
rect 12066 2796 12072 2848
rect 12124 2836 12130 2848
rect 12437 2839 12495 2845
rect 12437 2836 12449 2839
rect 12124 2808 12449 2836
rect 12124 2796 12130 2808
rect 12437 2805 12449 2808
rect 12483 2805 12495 2839
rect 12437 2799 12495 2805
rect 1104 2746 13892 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 12214 2746
rect 12266 2694 12278 2746
rect 12330 2694 12342 2746
rect 12394 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 13892 2746
rect 1104 2672 13892 2694
rect 3329 2635 3387 2641
rect 3329 2601 3341 2635
rect 3375 2632 3387 2635
rect 3418 2632 3424 2644
rect 3375 2604 3424 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 4614 2632 4620 2644
rect 4575 2604 4620 2632
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 6638 2632 6644 2644
rect 6599 2604 6644 2632
rect 6638 2592 6644 2604
rect 6696 2592 6702 2644
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 9582 2632 9588 2644
rect 9171 2604 9588 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 10502 2632 10508 2644
rect 10463 2604 10508 2632
rect 10502 2592 10508 2604
rect 10560 2592 10566 2644
rect 11238 2592 11244 2644
rect 11296 2632 11302 2644
rect 11793 2635 11851 2641
rect 11793 2632 11805 2635
rect 11296 2604 11805 2632
rect 11296 2592 11302 2604
rect 11793 2601 11805 2604
rect 11839 2601 11851 2635
rect 11793 2595 11851 2601
rect 7466 2564 7472 2576
rect 7427 2536 7472 2564
rect 7466 2524 7472 2536
rect 7524 2524 7530 2576
rect 7650 2564 7656 2576
rect 7576 2536 7656 2564
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 1857 2499 1915 2505
rect 1857 2465 1869 2499
rect 1903 2496 1915 2499
rect 2866 2496 2872 2508
rect 1903 2468 2872 2496
rect 1903 2465 1915 2468
rect 1857 2459 1915 2465
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 5166 2496 5172 2508
rect 5127 2468 5172 2496
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 7006 2496 7012 2508
rect 6967 2468 7012 2496
rect 7006 2456 7012 2468
rect 7064 2456 7070 2508
rect 7576 2505 7604 2536
rect 7650 2524 7656 2536
rect 7708 2524 7714 2576
rect 8110 2564 8116 2576
rect 8071 2536 8116 2564
rect 8110 2524 8116 2536
rect 8168 2524 8174 2576
rect 9490 2524 9496 2576
rect 9548 2564 9554 2576
rect 10870 2564 10876 2576
rect 9548 2536 10876 2564
rect 9548 2524 9554 2536
rect 10870 2524 10876 2536
rect 10928 2524 10934 2576
rect 13449 2567 13507 2573
rect 13449 2564 13461 2567
rect 11716 2536 13461 2564
rect 7561 2499 7619 2505
rect 7561 2465 7573 2499
rect 7607 2465 7619 2499
rect 7561 2459 7619 2465
rect 8757 2499 8815 2505
rect 8757 2465 8769 2499
rect 8803 2496 8815 2499
rect 9674 2496 9680 2508
rect 8803 2468 9680 2496
rect 8803 2465 8815 2468
rect 8757 2459 8815 2465
rect 9674 2456 9680 2468
rect 9732 2496 9738 2508
rect 10229 2499 10287 2505
rect 10229 2496 10241 2499
rect 9732 2468 10241 2496
rect 9732 2456 9738 2468
rect 10229 2465 10241 2468
rect 10275 2496 10287 2499
rect 10594 2496 10600 2508
rect 10275 2468 10600 2496
rect 10275 2465 10287 2468
rect 10229 2459 10287 2465
rect 10594 2456 10600 2468
rect 10652 2496 10658 2508
rect 10965 2499 11023 2505
rect 10965 2496 10977 2499
rect 10652 2468 10977 2496
rect 10652 2456 10658 2468
rect 10965 2465 10977 2468
rect 11011 2496 11023 2499
rect 11238 2496 11244 2508
rect 11011 2468 11244 2496
rect 11011 2465 11023 2468
rect 10965 2459 11023 2465
rect 11238 2456 11244 2468
rect 11296 2456 11302 2508
rect 11716 2505 11744 2536
rect 13449 2533 13461 2536
rect 13495 2533 13507 2567
rect 13449 2527 13507 2533
rect 11701 2499 11759 2505
rect 11701 2465 11713 2499
rect 11747 2465 11759 2499
rect 11701 2459 11759 2465
rect 11793 2499 11851 2505
rect 11793 2465 11805 2499
rect 11839 2496 11851 2499
rect 11974 2496 11980 2508
rect 11839 2468 11980 2496
rect 11839 2465 11851 2468
rect 11793 2459 11851 2465
rect 11974 2456 11980 2468
rect 12032 2456 12038 2508
rect 4157 2431 4215 2437
rect 4157 2397 4169 2431
rect 4203 2428 4215 2431
rect 4433 2431 4491 2437
rect 4433 2428 4445 2431
rect 4203 2400 4445 2428
rect 4203 2397 4215 2400
rect 4157 2391 4215 2397
rect 4433 2397 4445 2400
rect 4479 2428 4491 2431
rect 4893 2431 4951 2437
rect 4479 2400 4752 2428
rect 4479 2397 4491 2400
rect 4433 2391 4491 2397
rect 2590 2320 2596 2372
rect 2648 2320 2654 2372
rect 4341 2295 4399 2301
rect 4341 2261 4353 2295
rect 4387 2292 4399 2295
rect 4614 2292 4620 2304
rect 4387 2264 4620 2292
rect 4387 2261 4399 2264
rect 4341 2255 4399 2261
rect 4614 2252 4620 2264
rect 4672 2252 4678 2304
rect 4724 2292 4752 2400
rect 4893 2397 4905 2431
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2428 7711 2431
rect 7742 2428 7748 2440
rect 7699 2400 7748 2428
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 4908 2360 4936 2391
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2428 8079 2431
rect 8938 2428 8944 2440
rect 8067 2400 8944 2428
rect 8067 2397 8079 2400
rect 8021 2391 8079 2397
rect 8938 2388 8944 2400
rect 8996 2388 9002 2440
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 11054 2428 11060 2440
rect 10091 2400 11060 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 11149 2431 11207 2437
rect 11149 2397 11161 2431
rect 11195 2428 11207 2431
rect 11330 2428 11336 2440
rect 11195 2400 11336 2428
rect 11195 2397 11207 2400
rect 11149 2391 11207 2397
rect 11330 2388 11336 2400
rect 11388 2388 11394 2440
rect 11422 2388 11428 2440
rect 11480 2428 11486 2440
rect 12253 2431 12311 2437
rect 12253 2428 12265 2431
rect 11480 2400 12265 2428
rect 11480 2388 11486 2400
rect 12253 2397 12265 2400
rect 12299 2397 12311 2431
rect 12713 2431 12771 2437
rect 12713 2428 12725 2431
rect 12253 2391 12311 2397
rect 12636 2400 12725 2428
rect 5258 2360 5264 2372
rect 4908 2332 5264 2360
rect 5258 2320 5264 2332
rect 5316 2320 5322 2372
rect 5902 2320 5908 2372
rect 5960 2320 5966 2372
rect 8297 2363 8355 2369
rect 8297 2360 8309 2363
rect 8036 2332 8309 2360
rect 5810 2292 5816 2304
rect 4724 2264 5816 2292
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 8036 2301 8064 2332
rect 8297 2329 8309 2332
rect 8343 2360 8355 2363
rect 8570 2360 8576 2372
rect 8343 2332 8576 2360
rect 8343 2329 8355 2332
rect 8297 2323 8355 2329
rect 8570 2320 8576 2332
rect 8628 2320 8634 2372
rect 9306 2360 9312 2372
rect 9267 2332 9312 2360
rect 9306 2320 9312 2332
rect 9364 2320 9370 2372
rect 9493 2363 9551 2369
rect 9493 2329 9505 2363
rect 9539 2360 9551 2363
rect 9858 2360 9864 2372
rect 9539 2332 9864 2360
rect 9539 2329 9551 2332
rect 9493 2323 9551 2329
rect 9858 2320 9864 2332
rect 9916 2320 9922 2372
rect 10597 2363 10655 2369
rect 10597 2329 10609 2363
rect 10643 2329 10655 2363
rect 10778 2360 10784 2372
rect 10739 2332 10784 2360
rect 10597 2323 10655 2329
rect 6825 2295 6883 2301
rect 6825 2292 6837 2295
rect 6512 2264 6837 2292
rect 6512 2252 6518 2264
rect 6825 2261 6837 2264
rect 6871 2261 6883 2295
rect 6825 2255 6883 2261
rect 8021 2295 8079 2301
rect 8021 2261 8033 2295
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 9582 2252 9588 2304
rect 9640 2292 9646 2304
rect 9640 2264 9685 2292
rect 9640 2252 9646 2264
rect 9766 2252 9772 2304
rect 9824 2292 9830 2304
rect 9953 2295 10011 2301
rect 9953 2292 9965 2295
rect 9824 2264 9965 2292
rect 9824 2252 9830 2264
rect 9953 2261 9965 2264
rect 9999 2261 10011 2295
rect 10612 2292 10640 2323
rect 10778 2320 10784 2332
rect 10836 2320 10842 2372
rect 11606 2360 11612 2372
rect 11567 2332 11612 2360
rect 11606 2320 11612 2332
rect 11664 2320 11670 2372
rect 12636 2304 12664 2400
rect 12713 2397 12725 2400
rect 12759 2397 12771 2431
rect 12713 2391 12771 2397
rect 13078 2320 13084 2372
rect 13136 2360 13142 2372
rect 13173 2363 13231 2369
rect 13173 2360 13185 2363
rect 13136 2332 13185 2360
rect 13136 2320 13142 2332
rect 13173 2329 13185 2332
rect 13219 2329 13231 2363
rect 13173 2323 13231 2329
rect 11146 2292 11152 2304
rect 10612 2264 11152 2292
rect 9953 2255 10011 2261
rect 11146 2252 11152 2264
rect 11204 2252 11210 2304
rect 12066 2252 12072 2304
rect 12124 2292 12130 2304
rect 12161 2295 12219 2301
rect 12161 2292 12173 2295
rect 12124 2264 12173 2292
rect 12124 2252 12130 2264
rect 12161 2261 12173 2264
rect 12207 2261 12219 2295
rect 12618 2292 12624 2304
rect 12579 2264 12624 2292
rect 12161 2255 12219 2261
rect 12618 2252 12624 2264
rect 12676 2252 12682 2304
rect 13188 2292 13216 2323
rect 13262 2320 13268 2372
rect 13320 2360 13326 2372
rect 13320 2332 13365 2360
rect 13320 2320 13326 2332
rect 13357 2295 13415 2301
rect 13357 2292 13369 2295
rect 13188 2264 13369 2292
rect 13357 2261 13369 2264
rect 13403 2261 13415 2295
rect 13357 2255 13415 2261
rect 1104 2202 13892 2224
rect 1104 2150 8214 2202
rect 8266 2150 8278 2202
rect 8330 2150 8342 2202
rect 8394 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 13892 2202
rect 1104 2128 13892 2150
rect 5537 2091 5595 2097
rect 5537 2057 5549 2091
rect 5583 2088 5595 2091
rect 5718 2088 5724 2100
rect 5583 2060 5724 2088
rect 5583 2057 5595 2060
rect 5537 2051 5595 2057
rect 5718 2048 5724 2060
rect 5776 2048 5782 2100
rect 7742 2088 7748 2100
rect 6840 2060 7748 2088
rect 1578 2020 1584 2032
rect 1412 1992 1584 2020
rect 1412 1961 1440 1992
rect 1578 1980 1584 1992
rect 1636 1980 1642 2032
rect 2222 1980 2228 2032
rect 2280 1980 2286 2032
rect 3418 1980 3424 2032
rect 3476 2020 3482 2032
rect 6840 2029 6868 2060
rect 7742 2048 7748 2060
rect 7800 2048 7806 2100
rect 8938 2088 8944 2100
rect 8899 2060 8944 2088
rect 8938 2048 8944 2060
rect 8996 2048 9002 2100
rect 10042 2048 10048 2100
rect 10100 2088 10106 2100
rect 10965 2091 11023 2097
rect 10965 2088 10977 2091
rect 10100 2060 10977 2088
rect 10100 2048 10106 2060
rect 10965 2057 10977 2060
rect 11011 2057 11023 2091
rect 11330 2088 11336 2100
rect 11291 2060 11336 2088
rect 10965 2051 11023 2057
rect 11330 2048 11336 2060
rect 11388 2048 11394 2100
rect 6181 2023 6239 2029
rect 3476 1992 3726 2020
rect 3476 1980 3482 1992
rect 6181 1989 6193 2023
rect 6227 2020 6239 2023
rect 6825 2023 6883 2029
rect 6227 1992 6684 2020
rect 6227 1989 6239 1992
rect 6181 1983 6239 1989
rect 1397 1955 1455 1961
rect 1397 1921 1409 1955
rect 1443 1921 1455 1955
rect 1397 1915 1455 1921
rect 5169 1955 5227 1961
rect 5169 1921 5181 1955
rect 5215 1952 5227 1955
rect 5258 1952 5264 1964
rect 5215 1924 5264 1952
rect 5215 1921 5227 1924
rect 5169 1915 5227 1921
rect 5258 1912 5264 1924
rect 5316 1912 5322 1964
rect 5442 1912 5448 1964
rect 5500 1961 5506 1964
rect 5500 1955 5533 1961
rect 5521 1952 5533 1955
rect 5994 1952 6000 1964
rect 5521 1924 6000 1952
rect 5521 1921 5533 1924
rect 5500 1915 5533 1921
rect 5500 1912 5506 1915
rect 5994 1912 6000 1924
rect 6052 1912 6058 1964
rect 6454 1912 6460 1964
rect 6512 1952 6518 1964
rect 6656 1961 6684 1992
rect 6825 1989 6837 2023
rect 6871 1989 6883 2023
rect 6825 1983 6883 1989
rect 7116 1992 9812 2020
rect 6641 1955 6699 1961
rect 6512 1924 6605 1952
rect 6512 1912 6518 1924
rect 6641 1921 6653 1955
rect 6687 1952 6699 1955
rect 7116 1952 7144 1992
rect 6687 1924 7144 1952
rect 7193 1955 7251 1961
rect 6687 1921 6699 1924
rect 6641 1915 6699 1921
rect 7193 1921 7205 1955
rect 7239 1921 7251 1955
rect 7193 1915 7251 1921
rect 7285 1955 7343 1961
rect 7285 1921 7297 1955
rect 7331 1952 7343 1955
rect 7558 1952 7564 1964
rect 7331 1924 7564 1952
rect 7331 1921 7343 1924
rect 7285 1915 7343 1921
rect 1673 1887 1731 1893
rect 1673 1853 1685 1887
rect 1719 1884 1731 1887
rect 3050 1884 3056 1896
rect 1719 1856 3056 1884
rect 1719 1853 1731 1856
rect 1673 1847 1731 1853
rect 3050 1844 3056 1856
rect 3108 1844 3114 1896
rect 3145 1887 3203 1893
rect 3145 1853 3157 1887
rect 3191 1884 3203 1887
rect 4893 1887 4951 1893
rect 4893 1884 4905 1887
rect 3191 1856 4905 1884
rect 3191 1853 3203 1856
rect 3145 1847 3203 1853
rect 4893 1853 4905 1856
rect 4939 1853 4951 1887
rect 6472 1884 6500 1912
rect 4893 1847 4951 1853
rect 5230 1856 6500 1884
rect 7208 1884 7236 1915
rect 7558 1912 7564 1924
rect 7616 1912 7622 1964
rect 8757 1955 8815 1961
rect 8757 1921 8769 1955
rect 8803 1921 8815 1955
rect 8757 1915 8815 1921
rect 9309 1955 9367 1961
rect 9309 1921 9321 1955
rect 9355 1952 9367 1955
rect 9582 1952 9588 1964
rect 9355 1924 9588 1952
rect 9355 1921 9367 1924
rect 9309 1915 9367 1921
rect 8772 1884 8800 1915
rect 9582 1912 9588 1924
rect 9640 1912 9646 1964
rect 9784 1952 9812 1992
rect 9858 1980 9864 2032
rect 9916 2020 9922 2032
rect 9953 2023 10011 2029
rect 9953 2020 9965 2023
rect 9916 1992 9965 2020
rect 9916 1980 9922 1992
rect 9953 1989 9965 1992
rect 9999 1989 10011 2023
rect 10318 2020 10324 2032
rect 9953 1983 10011 1989
rect 10060 1992 10324 2020
rect 10060 1952 10088 1992
rect 10318 1980 10324 1992
rect 10376 1980 10382 2032
rect 9784 1924 10088 1952
rect 10229 1955 10287 1961
rect 10229 1921 10241 1955
rect 10275 1952 10287 1955
rect 10505 1955 10563 1961
rect 10505 1952 10517 1955
rect 10275 1924 10517 1952
rect 10275 1921 10287 1924
rect 10229 1915 10287 1921
rect 10505 1921 10517 1924
rect 10551 1921 10563 1955
rect 11348 1952 11376 2048
rect 12894 1980 12900 2032
rect 12952 2020 12958 2032
rect 13265 2023 13323 2029
rect 13265 2020 13277 2023
rect 12952 1992 13277 2020
rect 12952 1980 12958 1992
rect 13265 1989 13277 1992
rect 13311 1989 13323 2023
rect 13265 1983 13323 1989
rect 11517 1955 11575 1961
rect 11517 1952 11529 1955
rect 11348 1924 11529 1952
rect 10505 1915 10563 1921
rect 11517 1921 11529 1924
rect 11563 1921 11575 1955
rect 11517 1915 11575 1921
rect 12989 1955 13047 1961
rect 12989 1921 13001 1955
rect 13035 1921 13047 1955
rect 12989 1915 13047 1921
rect 10244 1884 10272 1915
rect 7208 1856 8616 1884
rect 8772 1856 10272 1884
rect 2866 1776 2872 1828
rect 2924 1816 2930 1828
rect 3421 1819 3479 1825
rect 3421 1816 3433 1819
rect 2924 1788 3433 1816
rect 2924 1776 2930 1788
rect 3421 1785 3433 1788
rect 3467 1785 3479 1819
rect 3421 1779 3479 1785
rect 934 1708 940 1760
rect 992 1748 998 1760
rect 5230 1748 5258 1856
rect 8588 1828 8616 1856
rect 5718 1776 5724 1828
rect 5776 1816 5782 1828
rect 5905 1819 5963 1825
rect 5905 1816 5917 1819
rect 5776 1788 5917 1816
rect 5776 1776 5782 1788
rect 5905 1785 5917 1788
rect 5951 1785 5963 1819
rect 8570 1816 8576 1828
rect 8531 1788 8576 1816
rect 5905 1779 5963 1785
rect 8570 1776 8576 1788
rect 8628 1776 8634 1828
rect 10520 1816 10548 1915
rect 10594 1844 10600 1896
rect 10652 1884 10658 1896
rect 10689 1887 10747 1893
rect 10689 1884 10701 1887
rect 10652 1856 10701 1884
rect 10652 1844 10658 1856
rect 10689 1853 10701 1856
rect 10735 1853 10747 1887
rect 10870 1884 10876 1896
rect 10831 1856 10876 1884
rect 10689 1847 10747 1853
rect 10870 1844 10876 1856
rect 10928 1844 10934 1896
rect 13004 1884 13032 1915
rect 13354 1884 13360 1896
rect 13004 1856 13360 1884
rect 13354 1844 13360 1856
rect 13412 1884 13418 1896
rect 13449 1887 13507 1893
rect 13449 1884 13461 1887
rect 13412 1856 13461 1884
rect 13412 1844 13418 1856
rect 13449 1853 13461 1856
rect 13495 1853 13507 1887
rect 13449 1847 13507 1853
rect 11606 1816 11612 1828
rect 10520 1788 11612 1816
rect 11606 1776 11612 1788
rect 11664 1816 11670 1828
rect 12805 1819 12863 1825
rect 12805 1816 12817 1819
rect 11664 1788 12817 1816
rect 11664 1776 11670 1788
rect 12805 1785 12817 1788
rect 12851 1785 12863 1819
rect 12805 1779 12863 1785
rect 5350 1748 5356 1760
rect 992 1720 5258 1748
rect 5311 1720 5356 1748
rect 992 1708 998 1720
rect 5350 1708 5356 1720
rect 5408 1708 5414 1760
rect 7006 1748 7012 1760
rect 6967 1720 7012 1748
rect 7006 1708 7012 1720
rect 7064 1708 7070 1760
rect 10318 1748 10324 1760
rect 10279 1720 10324 1748
rect 10318 1708 10324 1720
rect 10376 1708 10382 1760
rect 1104 1658 13892 1680
rect 1104 1606 4214 1658
rect 4266 1606 4278 1658
rect 4330 1606 4342 1658
rect 4394 1606 4406 1658
rect 4458 1606 4470 1658
rect 4522 1606 12214 1658
rect 12266 1606 12278 1658
rect 12330 1606 12342 1658
rect 12394 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 13892 1658
rect 1104 1584 13892 1606
rect 2222 1544 2228 1556
rect 2183 1516 2228 1544
rect 2222 1504 2228 1516
rect 2280 1504 2286 1556
rect 3418 1544 3424 1556
rect 3379 1516 3424 1544
rect 3418 1504 3424 1516
rect 3476 1504 3482 1556
rect 5810 1544 5816 1556
rect 4172 1516 5816 1544
rect 2041 1343 2099 1349
rect 2041 1309 2053 1343
rect 2087 1340 2099 1343
rect 2498 1340 2504 1352
rect 2087 1312 2504 1340
rect 2087 1309 2099 1312
rect 2041 1303 2099 1309
rect 2498 1300 2504 1312
rect 2556 1340 2562 1352
rect 3237 1343 3295 1349
rect 3237 1340 3249 1343
rect 2556 1312 3249 1340
rect 2556 1300 2562 1312
rect 3237 1309 3249 1312
rect 3283 1340 3295 1343
rect 4172 1340 4200 1516
rect 5810 1504 5816 1516
rect 5868 1504 5874 1556
rect 6546 1504 6552 1556
rect 6604 1544 6610 1556
rect 9490 1544 9496 1556
rect 6604 1516 9496 1544
rect 6604 1504 6610 1516
rect 9490 1504 9496 1516
rect 9548 1504 9554 1556
rect 10505 1547 10563 1553
rect 10505 1544 10517 1547
rect 9646 1516 10517 1544
rect 7558 1476 7564 1488
rect 7519 1448 7564 1476
rect 7558 1436 7564 1448
rect 7616 1436 7622 1488
rect 8570 1476 8576 1488
rect 8531 1448 8576 1476
rect 8570 1436 8576 1448
rect 8628 1436 8634 1488
rect 5350 1408 5356 1420
rect 5311 1380 5356 1408
rect 5350 1368 5356 1380
rect 5408 1368 5414 1420
rect 5810 1408 5816 1420
rect 5771 1380 5816 1408
rect 5810 1368 5816 1380
rect 5868 1368 5874 1420
rect 8665 1411 8723 1417
rect 6012 1380 7788 1408
rect 6012 1349 6040 1380
rect 7760 1352 7788 1380
rect 8665 1377 8677 1411
rect 8711 1408 8723 1411
rect 9306 1408 9312 1420
rect 8711 1380 9312 1408
rect 8711 1377 8723 1380
rect 8665 1371 8723 1377
rect 9306 1368 9312 1380
rect 9364 1368 9370 1420
rect 9493 1411 9551 1417
rect 9493 1377 9505 1411
rect 9539 1408 9551 1411
rect 9646 1408 9674 1516
rect 10505 1513 10517 1516
rect 10551 1544 10563 1547
rect 10594 1544 10600 1556
rect 10551 1516 10600 1544
rect 10551 1513 10563 1516
rect 10505 1507 10563 1513
rect 10594 1504 10600 1516
rect 10652 1544 10658 1556
rect 10781 1547 10839 1553
rect 10781 1544 10793 1547
rect 10652 1516 10793 1544
rect 10652 1504 10658 1516
rect 10781 1513 10793 1516
rect 10827 1544 10839 1547
rect 11793 1547 11851 1553
rect 11793 1544 11805 1547
rect 10827 1516 11805 1544
rect 10827 1513 10839 1516
rect 10781 1507 10839 1513
rect 11793 1513 11805 1516
rect 11839 1544 11851 1547
rect 12161 1547 12219 1553
rect 12161 1544 12173 1547
rect 11839 1516 12173 1544
rect 11839 1513 11851 1516
rect 11793 1507 11851 1513
rect 12161 1513 12173 1516
rect 12207 1513 12219 1547
rect 12161 1507 12219 1513
rect 13262 1504 13268 1556
rect 13320 1544 13326 1556
rect 13357 1547 13415 1553
rect 13357 1544 13369 1547
rect 13320 1516 13369 1544
rect 13320 1504 13326 1516
rect 13357 1513 13369 1516
rect 13403 1513 13415 1547
rect 13357 1507 13415 1513
rect 9858 1436 9864 1488
rect 9916 1476 9922 1488
rect 10229 1479 10287 1485
rect 10229 1476 10241 1479
rect 9916 1448 10241 1476
rect 9916 1436 9922 1448
rect 10229 1445 10241 1448
rect 10275 1445 10287 1479
rect 10229 1439 10287 1445
rect 10318 1408 10324 1420
rect 9539 1380 9674 1408
rect 10279 1380 10324 1408
rect 9539 1377 9551 1380
rect 9493 1371 9551 1377
rect 10318 1368 10324 1380
rect 10376 1368 10382 1420
rect 10965 1411 11023 1417
rect 10965 1377 10977 1411
rect 11011 1408 11023 1411
rect 11054 1408 11060 1420
rect 11011 1380 11060 1408
rect 11011 1377 11023 1380
rect 10965 1371 11023 1377
rect 11054 1368 11060 1380
rect 11112 1408 11118 1420
rect 13998 1408 14004 1420
rect 11112 1380 14004 1408
rect 11112 1368 11118 1380
rect 13998 1368 14004 1380
rect 14056 1368 14062 1420
rect 3283 1312 4200 1340
rect 5629 1343 5687 1349
rect 3283 1309 3295 1312
rect 3237 1303 3295 1309
rect 5629 1309 5641 1343
rect 5675 1309 5687 1343
rect 5629 1303 5687 1309
rect 5997 1343 6055 1349
rect 5997 1309 6009 1343
rect 6043 1309 6055 1343
rect 6178 1340 6184 1352
rect 6139 1312 6184 1340
rect 5997 1303 6055 1309
rect 2774 1232 2780 1284
rect 2832 1272 2838 1284
rect 3050 1272 3056 1284
rect 2832 1244 3056 1272
rect 2832 1232 2838 1244
rect 3050 1232 3056 1244
rect 3108 1272 3114 1284
rect 3513 1275 3571 1281
rect 3513 1272 3525 1275
rect 3108 1244 3525 1272
rect 3108 1232 3114 1244
rect 3513 1241 3525 1244
rect 3559 1241 3571 1275
rect 3513 1235 3571 1241
rect 4614 1232 4620 1284
rect 4672 1232 4678 1284
rect 5258 1232 5264 1284
rect 5316 1272 5322 1284
rect 5644 1272 5672 1303
rect 6178 1300 6184 1312
rect 6236 1300 6242 1352
rect 7006 1340 7012 1352
rect 6967 1312 7012 1340
rect 7006 1300 7012 1312
rect 7064 1300 7070 1352
rect 7742 1340 7748 1352
rect 7703 1312 7748 1340
rect 7742 1300 7748 1312
rect 7800 1300 7806 1352
rect 7929 1343 7987 1349
rect 7929 1309 7941 1343
rect 7975 1340 7987 1343
rect 8113 1343 8171 1349
rect 8113 1340 8125 1343
rect 7975 1312 8125 1340
rect 7975 1309 7987 1312
rect 7929 1303 7987 1309
rect 8113 1309 8125 1312
rect 8159 1340 8171 1343
rect 8159 1312 8984 1340
rect 8159 1309 8171 1312
rect 8113 1303 8171 1309
rect 6457 1275 6515 1281
rect 6457 1272 6469 1275
rect 5316 1244 6469 1272
rect 5316 1232 5322 1244
rect 6457 1241 6469 1244
rect 6503 1241 6515 1275
rect 6457 1235 6515 1241
rect 3881 1207 3939 1213
rect 3881 1173 3893 1207
rect 3927 1204 3939 1207
rect 5442 1204 5448 1216
rect 3927 1176 5448 1204
rect 3927 1173 3939 1176
rect 3881 1167 3939 1173
rect 5442 1164 5448 1176
rect 5500 1164 5506 1216
rect 8956 1213 8984 1312
rect 9582 1300 9588 1352
rect 9640 1340 9646 1352
rect 9769 1343 9827 1349
rect 9769 1340 9781 1343
rect 9640 1312 9781 1340
rect 9640 1300 9646 1312
rect 9769 1309 9781 1312
rect 9815 1309 9827 1343
rect 10686 1340 10692 1352
rect 9769 1303 9827 1309
rect 10060 1312 10692 1340
rect 9309 1275 9367 1281
rect 9309 1241 9321 1275
rect 9355 1272 9367 1275
rect 9950 1272 9956 1284
rect 9355 1244 9956 1272
rect 9355 1241 9367 1244
rect 9309 1235 9367 1241
rect 9950 1232 9956 1244
rect 10008 1232 10014 1284
rect 8941 1207 8999 1213
rect 8941 1173 8953 1207
rect 8987 1173 8999 1207
rect 8941 1167 8999 1173
rect 9401 1207 9459 1213
rect 9401 1173 9413 1207
rect 9447 1204 9459 1207
rect 10060 1204 10088 1312
rect 10686 1300 10692 1312
rect 10744 1300 10750 1352
rect 10870 1300 10876 1352
rect 10928 1340 10934 1352
rect 11698 1340 11704 1352
rect 10928 1312 11704 1340
rect 10928 1300 10934 1312
rect 11698 1300 11704 1312
rect 11756 1300 11762 1352
rect 12345 1343 12403 1349
rect 12345 1309 12357 1343
rect 12391 1340 12403 1343
rect 12618 1340 12624 1352
rect 12391 1312 12624 1340
rect 12391 1309 12403 1312
rect 12345 1303 12403 1309
rect 12618 1300 12624 1312
rect 12676 1300 12682 1352
rect 13078 1340 13084 1352
rect 13039 1312 13084 1340
rect 13078 1300 13084 1312
rect 13136 1300 13142 1352
rect 13265 1343 13323 1349
rect 13265 1309 13277 1343
rect 13311 1340 13323 1343
rect 13354 1340 13360 1352
rect 13311 1312 13360 1340
rect 13311 1309 13323 1312
rect 13265 1303 13323 1309
rect 13354 1300 13360 1312
rect 13412 1340 13418 1352
rect 13541 1343 13599 1349
rect 13541 1340 13553 1343
rect 13412 1312 13553 1340
rect 13412 1300 13418 1312
rect 13541 1309 13553 1312
rect 13587 1309 13599 1343
rect 13541 1303 13599 1309
rect 9447 1176 10088 1204
rect 9447 1173 9459 1176
rect 9401 1167 9459 1173
rect 1104 1114 13892 1136
rect 1104 1062 8214 1114
rect 8266 1062 8278 1114
rect 8330 1062 8342 1114
rect 8394 1062 8406 1114
rect 8458 1062 8470 1114
rect 8522 1062 13892 1114
rect 1104 1040 13892 1062
rect 13906 484 13912 536
rect 13964 524 13970 536
rect 14001 527 14059 533
rect 14001 524 14013 527
rect 13964 496 14013 524
rect 13964 484 13970 496
rect 14001 493 14013 496
rect 14047 493 14059 527
rect 14001 487 14059 493
<< via1 >>
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 12214 13574 12266 13626
rect 12278 13574 12330 13626
rect 12342 13574 12394 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 3148 13515 3200 13524
rect 3148 13481 3157 13515
rect 3157 13481 3191 13515
rect 3191 13481 3200 13515
rect 3148 13472 3200 13481
rect 8208 13472 8260 13524
rect 6736 13404 6788 13456
rect 7932 13336 7984 13388
rect 2044 13268 2096 13320
rect 2688 13268 2740 13320
rect 3332 13268 3384 13320
rect 6092 13268 6144 13320
rect 6920 13268 6972 13320
rect 7380 13311 7432 13320
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 7748 13311 7800 13320
rect 7748 13277 7757 13311
rect 7757 13277 7791 13311
rect 7791 13277 7800 13311
rect 7748 13268 7800 13277
rect 7840 13311 7892 13320
rect 7840 13277 7849 13311
rect 7849 13277 7883 13311
rect 7883 13277 7892 13311
rect 7840 13268 7892 13277
rect 8576 13268 8628 13320
rect 9404 13336 9456 13388
rect 9772 13472 9824 13524
rect 10876 13515 10928 13524
rect 10876 13481 10885 13515
rect 10885 13481 10919 13515
rect 10919 13481 10928 13515
rect 10876 13472 10928 13481
rect 9588 13404 9640 13456
rect 11152 13268 11204 13320
rect 12072 13311 12124 13320
rect 12072 13277 12081 13311
rect 12081 13277 12115 13311
rect 12115 13277 12124 13311
rect 12072 13268 12124 13277
rect 12624 13268 12676 13320
rect 8760 13200 8812 13252
rect 13176 13243 13228 13252
rect 13176 13209 13185 13243
rect 13185 13209 13219 13243
rect 13219 13209 13228 13243
rect 13176 13200 13228 13209
rect 13268 13243 13320 13252
rect 13268 13209 13277 13243
rect 13277 13209 13311 13243
rect 13311 13209 13320 13243
rect 13268 13200 13320 13209
rect 2596 13175 2648 13184
rect 2596 13141 2605 13175
rect 2605 13141 2639 13175
rect 2639 13141 2648 13175
rect 2596 13132 2648 13141
rect 3608 13132 3660 13184
rect 4620 13175 4672 13184
rect 4620 13141 4629 13175
rect 4629 13141 4663 13175
rect 4663 13141 4672 13175
rect 4620 13132 4672 13141
rect 7748 13132 7800 13184
rect 8024 13132 8076 13184
rect 9312 13175 9364 13184
rect 9312 13141 9321 13175
rect 9321 13141 9355 13175
rect 9355 13141 9364 13175
rect 10692 13175 10744 13184
rect 9312 13132 9364 13141
rect 10692 13141 10701 13175
rect 10701 13141 10735 13175
rect 10735 13141 10744 13175
rect 10692 13132 10744 13141
rect 11704 13175 11756 13184
rect 11704 13141 11713 13175
rect 11713 13141 11747 13175
rect 11747 13141 11756 13175
rect 11704 13132 11756 13141
rect 11980 13175 12032 13184
rect 11980 13141 11989 13175
rect 11989 13141 12023 13175
rect 12023 13141 12032 13175
rect 11980 13132 12032 13141
rect 13452 13175 13504 13184
rect 13452 13141 13461 13175
rect 13461 13141 13495 13175
rect 13495 13141 13504 13175
rect 13452 13132 13504 13141
rect 8214 13030 8266 13082
rect 8278 13030 8330 13082
rect 8342 13030 8394 13082
rect 8406 13030 8458 13082
rect 8470 13030 8522 13082
rect 2596 12860 2648 12912
rect 1860 12767 1912 12776
rect 1860 12733 1869 12767
rect 1869 12733 1903 12767
rect 1903 12733 1912 12767
rect 1860 12724 1912 12733
rect 3976 12860 4028 12912
rect 4620 12860 4672 12912
rect 7380 12928 7432 12980
rect 8116 12928 8168 12980
rect 9404 12971 9456 12980
rect 9404 12937 9413 12971
rect 9413 12937 9447 12971
rect 9447 12937 9456 12971
rect 9404 12928 9456 12937
rect 13268 12928 13320 12980
rect 6920 12860 6972 12912
rect 7104 12860 7156 12912
rect 3516 12724 3568 12776
rect 3976 12724 4028 12776
rect 4896 12724 4948 12776
rect 5632 12792 5684 12844
rect 5724 12724 5776 12776
rect 8024 12724 8076 12776
rect 9772 12860 9824 12912
rect 11152 12903 11204 12912
rect 11152 12869 11161 12903
rect 11161 12869 11195 12903
rect 11195 12869 11204 12903
rect 11152 12860 11204 12869
rect 8852 12792 8904 12844
rect 9588 12835 9640 12844
rect 9588 12801 9597 12835
rect 9597 12801 9631 12835
rect 9631 12801 9640 12835
rect 9588 12792 9640 12801
rect 10508 12835 10560 12844
rect 10508 12801 10517 12835
rect 10517 12801 10551 12835
rect 10551 12801 10560 12835
rect 10508 12792 10560 12801
rect 11704 12792 11756 12844
rect 13360 12792 13412 12844
rect 11704 12656 11756 12708
rect 13268 12656 13320 12708
rect 3516 12588 3568 12640
rect 5356 12631 5408 12640
rect 5356 12597 5365 12631
rect 5365 12597 5399 12631
rect 5399 12597 5408 12631
rect 5356 12588 5408 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 12214 12486 12266 12538
rect 12278 12486 12330 12538
rect 12342 12486 12394 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 2688 12316 2740 12368
rect 2964 12316 3016 12368
rect 7104 12384 7156 12436
rect 8576 12384 8628 12436
rect 9680 12384 9732 12436
rect 9864 12384 9916 12436
rect 11980 12316 12032 12368
rect 12072 12316 12124 12368
rect 13268 12316 13320 12368
rect 2872 12248 2924 12300
rect 2688 12180 2740 12232
rect 4528 12248 4580 12300
rect 7748 12291 7800 12300
rect 7748 12257 7757 12291
rect 7757 12257 7791 12291
rect 7791 12257 7800 12291
rect 7748 12248 7800 12257
rect 7932 12291 7984 12300
rect 7932 12257 7941 12291
rect 7941 12257 7975 12291
rect 7975 12257 7984 12291
rect 7932 12248 7984 12257
rect 1492 12155 1544 12164
rect 1492 12121 1501 12155
rect 1501 12121 1535 12155
rect 1535 12121 1544 12155
rect 1492 12112 1544 12121
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 3424 12180 3476 12232
rect 4068 12180 4120 12232
rect 3240 12112 3292 12164
rect 3516 12112 3568 12164
rect 6092 12180 6144 12232
rect 7380 12180 7432 12232
rect 8760 12248 8812 12300
rect 9036 12291 9088 12300
rect 9036 12257 9045 12291
rect 9045 12257 9079 12291
rect 9079 12257 9088 12291
rect 9036 12248 9088 12257
rect 11704 12291 11756 12300
rect 4436 12155 4488 12164
rect 3792 12044 3844 12096
rect 4436 12121 4445 12155
rect 4445 12121 4479 12155
rect 4479 12121 4488 12155
rect 4436 12112 4488 12121
rect 5724 12044 5776 12096
rect 5908 12087 5960 12096
rect 5908 12053 5917 12087
rect 5917 12053 5951 12087
rect 5951 12053 5960 12087
rect 5908 12044 5960 12053
rect 6920 12112 6972 12164
rect 7012 12044 7064 12096
rect 8024 12044 8076 12096
rect 8576 12112 8628 12164
rect 9588 12223 9640 12232
rect 9588 12189 9597 12223
rect 9597 12189 9631 12223
rect 9631 12189 9640 12223
rect 9588 12180 9640 12189
rect 9956 12180 10008 12232
rect 10692 12180 10744 12232
rect 9680 12112 9732 12164
rect 10508 12112 10560 12164
rect 8668 12044 8720 12096
rect 10876 12155 10928 12164
rect 10876 12121 10885 12155
rect 10885 12121 10919 12155
rect 10919 12121 10928 12155
rect 11704 12257 11713 12291
rect 11713 12257 11747 12291
rect 11747 12257 11756 12291
rect 11704 12248 11756 12257
rect 13452 12248 13504 12300
rect 11428 12223 11480 12232
rect 11428 12189 11437 12223
rect 11437 12189 11471 12223
rect 11471 12189 11480 12223
rect 11428 12180 11480 12189
rect 12624 12180 12676 12232
rect 13176 12223 13228 12232
rect 13176 12189 13185 12223
rect 13185 12189 13219 12223
rect 13219 12189 13228 12223
rect 13176 12180 13228 12189
rect 10876 12112 10928 12121
rect 10968 12044 11020 12096
rect 11612 12087 11664 12096
rect 11612 12053 11621 12087
rect 11621 12053 11655 12087
rect 11655 12053 11664 12087
rect 11612 12044 11664 12053
rect 13360 12112 13412 12164
rect 8214 11942 8266 11994
rect 8278 11942 8330 11994
rect 8342 11942 8394 11994
rect 8406 11942 8458 11994
rect 8470 11942 8522 11994
rect 1860 11840 1912 11892
rect 3608 11883 3660 11892
rect 3608 11849 3617 11883
rect 3617 11849 3651 11883
rect 3651 11849 3660 11883
rect 3608 11840 3660 11849
rect 2780 11704 2832 11756
rect 3056 11772 3108 11824
rect 2964 11704 3016 11756
rect 3332 11636 3384 11688
rect 4620 11815 4672 11824
rect 4620 11781 4629 11815
rect 4629 11781 4663 11815
rect 4663 11781 4672 11815
rect 5908 11840 5960 11892
rect 4620 11772 4672 11781
rect 3884 11747 3936 11756
rect 3884 11713 3893 11747
rect 3893 11713 3927 11747
rect 3927 11713 3936 11747
rect 3884 11704 3936 11713
rect 4344 11747 4396 11756
rect 4344 11713 4393 11747
rect 4393 11713 4396 11747
rect 4804 11747 4856 11756
rect 4344 11704 4396 11713
rect 4804 11713 4813 11747
rect 4813 11713 4847 11747
rect 4847 11713 4856 11747
rect 4804 11704 4856 11713
rect 5356 11704 5408 11756
rect 6000 11704 6052 11756
rect 4436 11568 4488 11620
rect 5172 11568 5224 11620
rect 4988 11543 5040 11552
rect 4988 11509 4997 11543
rect 4997 11509 5031 11543
rect 5031 11509 5040 11543
rect 4988 11500 5040 11509
rect 5264 11543 5316 11552
rect 5264 11509 5273 11543
rect 5273 11509 5307 11543
rect 5307 11509 5316 11543
rect 5264 11500 5316 11509
rect 8116 11772 8168 11824
rect 7012 11747 7064 11756
rect 7012 11713 7021 11747
rect 7021 11713 7055 11747
rect 7055 11713 7064 11747
rect 7012 11704 7064 11713
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 8484 11704 8536 11756
rect 9036 11772 9088 11824
rect 9680 11772 9732 11824
rect 10692 11840 10744 11892
rect 10968 11883 11020 11892
rect 7932 11568 7984 11620
rect 8024 11568 8076 11620
rect 7840 11543 7892 11552
rect 7840 11509 7849 11543
rect 7849 11509 7883 11543
rect 7883 11509 7892 11543
rect 7840 11500 7892 11509
rect 8208 11500 8260 11552
rect 9588 11704 9640 11756
rect 9772 11704 9824 11756
rect 10140 11704 10192 11756
rect 10508 11704 10560 11756
rect 10968 11849 10977 11883
rect 10977 11849 11011 11883
rect 11011 11849 11020 11883
rect 10968 11840 11020 11849
rect 13268 11815 13320 11824
rect 13268 11781 13277 11815
rect 13277 11781 13311 11815
rect 13311 11781 13320 11815
rect 13268 11772 13320 11781
rect 10876 11704 10928 11756
rect 11060 11747 11112 11756
rect 11060 11713 11069 11747
rect 11069 11713 11103 11747
rect 11103 11713 11112 11747
rect 11060 11704 11112 11713
rect 13452 11747 13504 11756
rect 8668 11568 8720 11620
rect 9864 11679 9916 11688
rect 9864 11645 9873 11679
rect 9873 11645 9907 11679
rect 9907 11645 9916 11679
rect 9864 11636 9916 11645
rect 13452 11713 13461 11747
rect 13461 11713 13495 11747
rect 13495 11713 13504 11747
rect 13452 11704 13504 11713
rect 11888 11636 11940 11688
rect 10784 11568 10836 11620
rect 12808 11611 12860 11620
rect 12808 11577 12817 11611
rect 12817 11577 12851 11611
rect 12851 11577 12860 11611
rect 12808 11568 12860 11577
rect 9956 11500 10008 11552
rect 10968 11500 11020 11552
rect 11428 11500 11480 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 12214 11398 12266 11450
rect 12278 11398 12330 11450
rect 12342 11398 12394 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 3148 11296 3200 11348
rect 2596 11160 2648 11212
rect 3332 11228 3384 11280
rect 3976 11296 4028 11348
rect 6920 11296 6972 11348
rect 7012 11296 7064 11348
rect 7380 11296 7432 11348
rect 7932 11296 7984 11348
rect 5448 11228 5500 11280
rect 3332 11135 3384 11144
rect 3332 11101 3341 11135
rect 3341 11101 3375 11135
rect 3375 11101 3384 11135
rect 3792 11135 3844 11144
rect 3332 11092 3384 11101
rect 3792 11101 3801 11135
rect 3801 11101 3835 11135
rect 3835 11101 3844 11135
rect 3792 11092 3844 11101
rect 3884 11092 3936 11144
rect 4068 11092 4120 11144
rect 4344 11160 4396 11212
rect 5264 11160 5316 11212
rect 4620 11092 4672 11144
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 4896 11092 4948 11144
rect 5632 11092 5684 11144
rect 2228 11024 2280 11076
rect 2964 11067 3016 11076
rect 2964 11033 2973 11067
rect 2973 11033 3007 11067
rect 3007 11033 3016 11067
rect 2964 11024 3016 11033
rect 5172 11067 5224 11076
rect 5172 11033 5181 11067
rect 5181 11033 5215 11067
rect 5215 11033 5224 11067
rect 5172 11024 5224 11033
rect 5908 11160 5960 11212
rect 7840 11228 7892 11280
rect 756 10956 808 11008
rect 2780 10956 2832 11008
rect 3332 10956 3384 11008
rect 4252 10956 4304 11008
rect 4896 10956 4948 11008
rect 6000 11067 6052 11076
rect 6000 11033 6009 11067
rect 6009 11033 6043 11067
rect 6043 11033 6052 11067
rect 7104 11160 7156 11212
rect 8208 11160 8260 11212
rect 6552 11092 6604 11144
rect 7012 11092 7064 11144
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8116 11092 8168 11101
rect 9864 11296 9916 11348
rect 11060 11228 11112 11280
rect 12440 11228 12492 11280
rect 12808 11228 12860 11280
rect 6000 11024 6052 11033
rect 6644 10956 6696 11008
rect 6920 11024 6972 11076
rect 8760 11092 8812 11144
rect 9680 11160 9732 11212
rect 11888 11203 11940 11212
rect 11888 11169 11897 11203
rect 11897 11169 11931 11203
rect 11931 11169 11940 11203
rect 11888 11160 11940 11169
rect 9772 11092 9824 11144
rect 9680 11024 9732 11076
rect 7012 10956 7064 11008
rect 8576 10956 8628 11008
rect 10600 10956 10652 11008
rect 10692 10956 10744 11008
rect 12716 11092 12768 11144
rect 13452 11135 13504 11144
rect 13452 11101 13461 11135
rect 13461 11101 13495 11135
rect 13495 11101 13504 11135
rect 13452 11092 13504 11101
rect 12808 11024 12860 11076
rect 13176 11067 13228 11076
rect 13176 11033 13185 11067
rect 13185 11033 13219 11067
rect 13219 11033 13228 11067
rect 13176 11024 13228 11033
rect 8214 10854 8266 10906
rect 8278 10854 8330 10906
rect 8342 10854 8394 10906
rect 8406 10854 8458 10906
rect 8470 10854 8522 10906
rect 2228 10795 2280 10804
rect 2228 10761 2237 10795
rect 2237 10761 2271 10795
rect 2271 10761 2280 10795
rect 2228 10752 2280 10761
rect 2964 10752 3016 10804
rect 4068 10795 4120 10804
rect 2596 10727 2648 10736
rect 2596 10693 2605 10727
rect 2605 10693 2639 10727
rect 2639 10693 2648 10727
rect 2596 10684 2648 10693
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 2412 10659 2464 10668
rect 2412 10625 2421 10659
rect 2421 10625 2455 10659
rect 2455 10625 2464 10659
rect 2412 10616 2464 10625
rect 2872 10659 2924 10668
rect 2872 10625 2875 10659
rect 2875 10625 2924 10659
rect 1492 10548 1544 10600
rect 2872 10616 2924 10625
rect 3148 10616 3200 10668
rect 3332 10616 3384 10668
rect 3609 10659 3661 10668
rect 3792 10684 3844 10736
rect 4068 10761 4077 10795
rect 4077 10761 4111 10795
rect 4111 10761 4120 10795
rect 4068 10752 4120 10761
rect 4252 10752 4304 10804
rect 3976 10684 4028 10736
rect 4988 10752 5040 10804
rect 7840 10752 7892 10804
rect 8760 10752 8812 10804
rect 9128 10752 9180 10804
rect 10324 10795 10376 10804
rect 10324 10761 10333 10795
rect 10333 10761 10367 10795
rect 10367 10761 10376 10795
rect 10324 10752 10376 10761
rect 3609 10625 3622 10659
rect 3622 10625 3656 10659
rect 3656 10625 3661 10659
rect 3609 10616 3661 10625
rect 3056 10548 3108 10600
rect 3792 10548 3844 10600
rect 4528 10616 4580 10668
rect 4896 10659 4948 10668
rect 4896 10625 4905 10659
rect 4905 10625 4939 10659
rect 4939 10625 4948 10659
rect 4896 10616 4948 10625
rect 5264 10616 5316 10668
rect 5816 10616 5868 10668
rect 4344 10548 4396 10600
rect 6552 10616 6604 10668
rect 6920 10659 6972 10668
rect 6920 10625 6929 10659
rect 6929 10625 6963 10659
rect 6963 10625 6972 10659
rect 6920 10616 6972 10625
rect 7196 10684 7248 10736
rect 10140 10727 10192 10736
rect 7472 10616 7524 10668
rect 7656 10659 7708 10668
rect 7656 10625 7665 10659
rect 7665 10625 7699 10659
rect 7699 10625 7708 10659
rect 7656 10616 7708 10625
rect 7840 10659 7892 10668
rect 7840 10625 7849 10659
rect 7849 10625 7883 10659
rect 7883 10625 7892 10659
rect 7840 10616 7892 10625
rect 8024 10659 8076 10668
rect 8024 10625 8033 10659
rect 8033 10625 8067 10659
rect 8067 10625 8076 10659
rect 8024 10616 8076 10625
rect 8392 10659 8444 10668
rect 8392 10625 8401 10659
rect 8401 10625 8435 10659
rect 8435 10625 8444 10659
rect 8392 10616 8444 10625
rect 9036 10616 9088 10668
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 10140 10693 10149 10727
rect 10149 10693 10183 10727
rect 10183 10693 10192 10727
rect 10140 10684 10192 10693
rect 11060 10727 11112 10736
rect 11060 10693 11069 10727
rect 11069 10693 11103 10727
rect 11103 10693 11112 10727
rect 11060 10684 11112 10693
rect 12440 10727 12492 10736
rect 12440 10693 12449 10727
rect 12449 10693 12483 10727
rect 12483 10693 12492 10727
rect 12440 10684 12492 10693
rect 13176 10727 13228 10736
rect 13176 10693 13185 10727
rect 13185 10693 13219 10727
rect 13219 10693 13228 10727
rect 13176 10684 13228 10693
rect 9128 10616 9180 10625
rect 9220 10548 9272 10600
rect 9772 10659 9824 10668
rect 9772 10625 9781 10659
rect 9781 10625 9815 10659
rect 9815 10625 9824 10659
rect 9772 10616 9824 10625
rect 9956 10659 10008 10668
rect 9956 10625 9965 10659
rect 9965 10625 9999 10659
rect 9999 10625 10008 10659
rect 10600 10659 10652 10668
rect 9956 10616 10008 10625
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 10692 10616 10744 10668
rect 11612 10616 11664 10668
rect 13452 10616 13504 10668
rect 2320 10480 2372 10532
rect 2964 10455 3016 10464
rect 2964 10421 2973 10455
rect 2973 10421 3007 10455
rect 3007 10421 3016 10455
rect 2964 10412 3016 10421
rect 3608 10412 3660 10464
rect 5172 10412 5224 10464
rect 5540 10412 5592 10464
rect 6368 10412 6420 10464
rect 12716 10591 12768 10600
rect 12716 10557 12725 10591
rect 12725 10557 12759 10591
rect 12759 10557 12768 10591
rect 12716 10548 12768 10557
rect 12624 10523 12676 10532
rect 12624 10489 12633 10523
rect 12633 10489 12667 10523
rect 12667 10489 12676 10523
rect 12624 10480 12676 10489
rect 7012 10412 7064 10464
rect 7932 10455 7984 10464
rect 7932 10421 7941 10455
rect 7941 10421 7975 10455
rect 7975 10421 7984 10455
rect 7932 10412 7984 10421
rect 8392 10412 8444 10464
rect 10508 10455 10560 10464
rect 10508 10421 10517 10455
rect 10517 10421 10551 10455
rect 10551 10421 10560 10455
rect 10508 10412 10560 10421
rect 11796 10412 11848 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 12214 10310 12266 10362
rect 12278 10310 12330 10362
rect 12342 10310 12394 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 1492 10251 1544 10260
rect 1492 10217 1501 10251
rect 1501 10217 1535 10251
rect 1535 10217 1544 10251
rect 1492 10208 1544 10217
rect 2780 10208 2832 10260
rect 6920 10251 6972 10260
rect 3884 10140 3936 10192
rect 4068 10183 4120 10192
rect 4068 10149 4077 10183
rect 4077 10149 4111 10183
rect 4111 10149 4120 10183
rect 4068 10140 4120 10149
rect 2964 10115 3016 10124
rect 2964 10081 2973 10115
rect 2973 10081 3007 10115
rect 3007 10081 3016 10115
rect 2964 10072 3016 10081
rect 3424 10072 3476 10124
rect 4620 10140 4672 10192
rect 6920 10217 6929 10251
rect 6929 10217 6963 10251
rect 6963 10217 6972 10251
rect 6920 10208 6972 10217
rect 7656 10208 7708 10260
rect 7748 10208 7800 10260
rect 8208 10208 8260 10260
rect 8944 10208 8996 10260
rect 9036 10208 9088 10260
rect 7472 10140 7524 10192
rect 3608 10004 3660 10056
rect 3976 10004 4028 10056
rect 4896 10072 4948 10124
rect 5448 10115 5500 10124
rect 5448 10081 5457 10115
rect 5457 10081 5491 10115
rect 5491 10081 5500 10115
rect 5448 10072 5500 10081
rect 6644 10072 6696 10124
rect 7380 10072 7432 10124
rect 8576 10140 8628 10192
rect 9220 10140 9272 10192
rect 8760 10072 8812 10124
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 7288 10004 7340 10056
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 8392 10004 8444 10056
rect 10508 10208 10560 10260
rect 12808 10208 12860 10260
rect 2228 9936 2280 9988
rect 5724 9936 5776 9988
rect 5908 9936 5960 9988
rect 7012 9936 7064 9988
rect 10048 10140 10100 10192
rect 11796 10115 11848 10124
rect 11796 10081 11805 10115
rect 11805 10081 11839 10115
rect 11839 10081 11848 10115
rect 11796 10072 11848 10081
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 12440 10047 12492 10056
rect 12440 10013 12449 10047
rect 12449 10013 12483 10047
rect 12483 10013 12492 10047
rect 12440 10004 12492 10013
rect 13176 10004 13228 10056
rect 3516 9868 3568 9920
rect 7196 9868 7248 9920
rect 7472 9868 7524 9920
rect 10692 9936 10744 9988
rect 11612 9936 11664 9988
rect 12900 9979 12952 9988
rect 12900 9945 12909 9979
rect 12909 9945 12943 9979
rect 12943 9945 12952 9979
rect 12900 9936 12952 9945
rect 9680 9868 9732 9920
rect 13360 9911 13412 9920
rect 13360 9877 13369 9911
rect 13369 9877 13403 9911
rect 13403 9877 13412 9911
rect 13360 9868 13412 9877
rect 8214 9766 8266 9818
rect 8278 9766 8330 9818
rect 8342 9766 8394 9818
rect 8406 9766 8458 9818
rect 8470 9766 8522 9818
rect 2228 9664 2280 9716
rect 2872 9596 2924 9648
rect 2044 9528 2096 9580
rect 3240 9596 3292 9648
rect 3148 9571 3200 9580
rect 3148 9537 3156 9571
rect 3156 9537 3190 9571
rect 3190 9537 3200 9571
rect 3148 9528 3200 9537
rect 3976 9664 4028 9716
rect 5540 9707 5592 9716
rect 5540 9673 5549 9707
rect 5549 9673 5583 9707
rect 5583 9673 5592 9707
rect 5540 9664 5592 9673
rect 7196 9664 7248 9716
rect 4804 9596 4856 9648
rect 6644 9596 6696 9648
rect 3608 9528 3660 9580
rect 6000 9571 6052 9580
rect 6000 9537 6009 9571
rect 6009 9537 6043 9571
rect 6043 9537 6052 9571
rect 6000 9528 6052 9537
rect 7288 9596 7340 9648
rect 14188 9664 14240 9716
rect 8392 9596 8444 9648
rect 13360 9596 13412 9648
rect 3424 9460 3476 9512
rect 5356 9460 5408 9512
rect 7012 9528 7064 9580
rect 7196 9571 7248 9580
rect 7196 9537 7205 9571
rect 7205 9537 7239 9571
rect 7239 9537 7248 9571
rect 7196 9528 7248 9537
rect 6552 9503 6604 9512
rect 6552 9469 6561 9503
rect 6561 9469 6595 9503
rect 6595 9469 6604 9503
rect 6552 9460 6604 9469
rect 6644 9460 6696 9512
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 8024 9528 8076 9580
rect 8944 9528 8996 9580
rect 8484 9503 8536 9512
rect 8484 9469 8493 9503
rect 8493 9469 8527 9503
rect 8527 9469 8536 9503
rect 8484 9460 8536 9469
rect 6000 9392 6052 9444
rect 7380 9392 7432 9444
rect 10048 9571 10100 9580
rect 10048 9537 10057 9571
rect 10057 9537 10091 9571
rect 10091 9537 10100 9571
rect 10048 9528 10100 9537
rect 11520 9528 11572 9580
rect 12440 9528 12492 9580
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 13084 9528 13136 9580
rect 10600 9460 10652 9512
rect 10508 9392 10560 9444
rect 12900 9435 12952 9444
rect 12900 9401 12909 9435
rect 12909 9401 12943 9435
rect 12943 9401 12952 9435
rect 12900 9392 12952 9401
rect 4068 9324 4120 9376
rect 6460 9367 6512 9376
rect 6460 9333 6469 9367
rect 6469 9333 6503 9367
rect 6503 9333 6512 9367
rect 6460 9324 6512 9333
rect 6552 9324 6604 9376
rect 7472 9324 7524 9376
rect 9036 9367 9088 9376
rect 9036 9333 9045 9367
rect 9045 9333 9079 9367
rect 9079 9333 9088 9367
rect 9036 9324 9088 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 12214 9222 12266 9274
rect 12278 9222 12330 9274
rect 12342 9222 12394 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 4804 9120 4856 9172
rect 3148 9095 3200 9104
rect 3148 9061 3157 9095
rect 3157 9061 3191 9095
rect 3191 9061 3200 9095
rect 3148 9052 3200 9061
rect 4068 8984 4120 9036
rect 6644 9120 6696 9172
rect 7196 9120 7248 9172
rect 7472 9163 7524 9172
rect 7472 9129 7481 9163
rect 7481 9129 7515 9163
rect 7515 9129 7524 9163
rect 7472 9120 7524 9129
rect 8392 9163 8444 9172
rect 8392 9129 8401 9163
rect 8401 9129 8435 9163
rect 8435 9129 8444 9163
rect 8392 9120 8444 9129
rect 8484 9120 8536 9172
rect 9680 9120 9732 9172
rect 11520 9163 11572 9172
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 3792 8959 3844 8968
rect 3792 8925 3801 8959
rect 3801 8925 3835 8959
rect 3835 8925 3844 8959
rect 3792 8916 3844 8925
rect 4436 8959 4488 8968
rect 2412 8848 2464 8900
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 6920 9052 6972 9104
rect 5356 8984 5408 9036
rect 10692 9095 10744 9104
rect 10692 9061 10701 9095
rect 10701 9061 10735 9095
rect 10735 9061 10744 9095
rect 10692 9052 10744 9061
rect 11520 9129 11529 9163
rect 11529 9129 11563 9163
rect 11563 9129 11572 9163
rect 11520 9120 11572 9129
rect 9036 8984 9088 9036
rect 12624 9052 12676 9104
rect 10876 9027 10928 9036
rect 10876 8993 10885 9027
rect 10885 8993 10919 9027
rect 10919 8993 10928 9027
rect 10876 8984 10928 8993
rect 11244 8984 11296 9036
rect 4620 8916 4672 8968
rect 5264 8891 5316 8900
rect 5264 8857 5273 8891
rect 5273 8857 5307 8891
rect 5307 8857 5316 8891
rect 5264 8848 5316 8857
rect 6000 8848 6052 8900
rect 8576 8916 8628 8968
rect 10508 8959 10560 8968
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 10600 8916 10652 8968
rect 13360 9052 13412 9104
rect 12900 8916 12952 8968
rect 8024 8848 8076 8900
rect 13084 8891 13136 8900
rect 13084 8857 13093 8891
rect 13093 8857 13127 8891
rect 13127 8857 13136 8891
rect 13084 8848 13136 8857
rect 13176 8891 13228 8900
rect 13176 8857 13185 8891
rect 13185 8857 13219 8891
rect 13219 8857 13228 8891
rect 13176 8848 13228 8857
rect 3792 8780 3844 8832
rect 4896 8780 4948 8832
rect 6736 8823 6788 8832
rect 6736 8789 6745 8823
rect 6745 8789 6779 8823
rect 6779 8789 6788 8823
rect 6736 8780 6788 8789
rect 7472 8780 7524 8832
rect 9588 8823 9640 8832
rect 9588 8789 9597 8823
rect 9597 8789 9631 8823
rect 9631 8789 9640 8823
rect 9588 8780 9640 8789
rect 11152 8823 11204 8832
rect 11152 8789 11161 8823
rect 11161 8789 11195 8823
rect 11195 8789 11204 8823
rect 11152 8780 11204 8789
rect 8214 8678 8266 8730
rect 8278 8678 8330 8730
rect 8342 8678 8394 8730
rect 8406 8678 8458 8730
rect 8470 8678 8522 8730
rect 2412 8576 2464 8628
rect 3792 8576 3844 8628
rect 4620 8576 4672 8628
rect 5908 8576 5960 8628
rect 6000 8576 6052 8628
rect 3424 8551 3476 8560
rect 3424 8517 3433 8551
rect 3433 8517 3467 8551
rect 3467 8517 3476 8551
rect 3424 8508 3476 8517
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 2228 8347 2280 8356
rect 2228 8313 2237 8347
rect 2237 8313 2271 8347
rect 2271 8313 2280 8347
rect 2228 8304 2280 8313
rect 3240 8440 3292 8492
rect 3700 8440 3752 8492
rect 3976 8440 4028 8492
rect 4712 8508 4764 8560
rect 6736 8508 6788 8560
rect 10048 8576 10100 8628
rect 12624 8619 12676 8628
rect 9588 8508 9640 8560
rect 4620 8483 4672 8492
rect 4620 8449 4629 8483
rect 4629 8449 4663 8483
rect 4663 8449 4672 8483
rect 4620 8440 4672 8449
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 5356 8483 5408 8492
rect 5356 8449 5359 8483
rect 5359 8449 5408 8483
rect 4436 8372 4488 8424
rect 5356 8440 5408 8449
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 7196 8440 7248 8492
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 8668 8483 8720 8492
rect 8668 8449 8677 8483
rect 8677 8449 8711 8483
rect 8711 8449 8720 8483
rect 8668 8440 8720 8449
rect 12624 8585 12633 8619
rect 12633 8585 12667 8619
rect 12667 8585 12676 8619
rect 12624 8576 12676 8585
rect 12716 8576 12768 8628
rect 12900 8508 12952 8560
rect 7748 8372 7800 8424
rect 11520 8440 11572 8492
rect 13084 8440 13136 8492
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 4804 8347 4856 8356
rect 4804 8313 4813 8347
rect 4813 8313 4847 8347
rect 4847 8313 4856 8347
rect 4804 8304 4856 8313
rect 5264 8304 5316 8356
rect 8760 8347 8812 8356
rect 8760 8313 8769 8347
rect 8769 8313 8803 8347
rect 8803 8313 8812 8347
rect 8760 8304 8812 8313
rect 11796 8372 11848 8424
rect 12624 8372 12676 8424
rect 13268 8415 13320 8424
rect 13268 8381 13277 8415
rect 13277 8381 13311 8415
rect 13311 8381 13320 8415
rect 13268 8372 13320 8381
rect 4068 8236 4120 8288
rect 4620 8236 4672 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 12214 8134 12266 8186
rect 12278 8134 12330 8186
rect 12342 8134 12394 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 3424 8032 3476 8084
rect 4712 8032 4764 8084
rect 9312 8032 9364 8084
rect 5080 7964 5132 8016
rect 8760 7964 8812 8016
rect 9220 7964 9272 8016
rect 9956 8032 10008 8084
rect 13268 8032 13320 8084
rect 10048 7964 10100 8016
rect 11152 7964 11204 8016
rect 12624 7964 12676 8016
rect 4068 7939 4120 7948
rect 4068 7905 4077 7939
rect 4077 7905 4111 7939
rect 4111 7905 4120 7939
rect 4068 7896 4120 7905
rect 4160 7896 4212 7948
rect 5356 7896 5408 7948
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 9496 7896 9548 7948
rect 6460 7828 6512 7880
rect 7104 7828 7156 7880
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 7472 7828 7524 7880
rect 8668 7871 8720 7880
rect 8668 7837 8677 7871
rect 8677 7837 8711 7871
rect 8711 7837 8720 7871
rect 8668 7828 8720 7837
rect 8944 7828 8996 7880
rect 9404 7871 9456 7880
rect 9404 7837 9413 7871
rect 9413 7837 9447 7871
rect 9447 7837 9456 7871
rect 9404 7828 9456 7837
rect 1676 7803 1728 7812
rect 1676 7769 1685 7803
rect 1685 7769 1719 7803
rect 1719 7769 1728 7803
rect 1676 7760 1728 7769
rect 2228 7760 2280 7812
rect 4804 7760 4856 7812
rect 6644 7760 6696 7812
rect 9128 7760 9180 7812
rect 10692 7828 10744 7880
rect 11520 7871 11572 7880
rect 11520 7837 11529 7871
rect 11529 7837 11563 7871
rect 11563 7837 11572 7871
rect 11520 7828 11572 7837
rect 11796 7871 11848 7880
rect 11796 7837 11805 7871
rect 11805 7837 11839 7871
rect 11839 7837 11848 7871
rect 11796 7828 11848 7837
rect 13176 7871 13228 7880
rect 13176 7837 13185 7871
rect 13185 7837 13219 7871
rect 13219 7837 13228 7871
rect 13176 7828 13228 7837
rect 10048 7760 10100 7812
rect 10324 7803 10376 7812
rect 10324 7769 10333 7803
rect 10333 7769 10367 7803
rect 10367 7769 10376 7803
rect 10324 7760 10376 7769
rect 7012 7735 7064 7744
rect 7012 7701 7021 7735
rect 7021 7701 7055 7735
rect 7055 7701 7064 7735
rect 7012 7692 7064 7701
rect 7564 7735 7616 7744
rect 7564 7701 7573 7735
rect 7573 7701 7607 7735
rect 7607 7701 7616 7735
rect 7564 7692 7616 7701
rect 7656 7692 7708 7744
rect 8760 7692 8812 7744
rect 11796 7692 11848 7744
rect 8214 7590 8266 7642
rect 8278 7590 8330 7642
rect 8342 7590 8394 7642
rect 8406 7590 8458 7642
rect 8470 7590 8522 7642
rect 1676 7488 1728 7540
rect 3516 7488 3568 7540
rect 4068 7488 4120 7540
rect 4620 7488 4672 7540
rect 2320 7420 2372 7472
rect 3792 7463 3844 7472
rect 3792 7429 3801 7463
rect 3801 7429 3835 7463
rect 3835 7429 3844 7463
rect 3792 7420 3844 7429
rect 3424 7352 3476 7404
rect 3516 7395 3568 7404
rect 3516 7361 3565 7395
rect 3565 7361 3568 7395
rect 3516 7352 3568 7361
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 2412 7284 2464 7336
rect 3148 7327 3200 7336
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 3148 7284 3200 7293
rect 7932 7488 7984 7540
rect 8576 7531 8628 7540
rect 8576 7497 8585 7531
rect 8585 7497 8619 7531
rect 8619 7497 8628 7531
rect 8576 7488 8628 7497
rect 9404 7531 9456 7540
rect 9404 7497 9413 7531
rect 9413 7497 9447 7531
rect 9447 7497 9456 7531
rect 9404 7488 9456 7497
rect 10876 7488 10928 7540
rect 11888 7488 11940 7540
rect 12808 7488 12860 7540
rect 6460 7420 6512 7472
rect 7564 7420 7616 7472
rect 5080 7352 5132 7404
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 6000 7395 6052 7404
rect 6000 7361 6009 7395
rect 6009 7361 6043 7395
rect 6043 7361 6052 7395
rect 6000 7352 6052 7361
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 7472 7395 7524 7404
rect 7472 7361 7481 7395
rect 7481 7361 7515 7395
rect 7515 7361 7524 7395
rect 7472 7352 7524 7361
rect 8392 7395 8444 7404
rect 8392 7361 8401 7395
rect 8401 7361 8435 7395
rect 8435 7361 8444 7395
rect 8392 7352 8444 7361
rect 8668 7352 8720 7404
rect 9312 7420 9364 7472
rect 9588 7420 9640 7472
rect 9956 7420 10008 7472
rect 10324 7420 10376 7472
rect 4712 7327 4764 7336
rect 4712 7293 4721 7327
rect 4721 7293 4755 7327
rect 4755 7293 4764 7327
rect 4712 7284 4764 7293
rect 4896 7284 4948 7336
rect 6644 7284 6696 7336
rect 7656 7284 7708 7336
rect 9772 7352 9824 7404
rect 10048 7395 10100 7404
rect 10048 7361 10057 7395
rect 10057 7361 10091 7395
rect 10091 7361 10100 7395
rect 10048 7352 10100 7361
rect 12900 7463 12952 7472
rect 12900 7429 12909 7463
rect 12909 7429 12943 7463
rect 12943 7429 12952 7463
rect 12900 7420 12952 7429
rect 11796 7395 11848 7404
rect 9128 7284 9180 7336
rect 9312 7284 9364 7336
rect 5724 7259 5776 7268
rect 5724 7225 5733 7259
rect 5733 7225 5767 7259
rect 5767 7225 5776 7259
rect 5724 7216 5776 7225
rect 4988 7148 5040 7200
rect 5816 7148 5868 7200
rect 6368 7148 6420 7200
rect 8668 7216 8720 7268
rect 9036 7216 9088 7268
rect 9864 7216 9916 7268
rect 10232 7216 10284 7268
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 11796 7352 11848 7361
rect 11336 7191 11388 7200
rect 11336 7157 11345 7191
rect 11345 7157 11379 7191
rect 11379 7157 11388 7191
rect 11336 7148 11388 7157
rect 11612 7191 11664 7200
rect 11612 7157 11621 7191
rect 11621 7157 11655 7191
rect 11655 7157 11664 7191
rect 11612 7148 11664 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 12214 7046 12266 7098
rect 12278 7046 12330 7098
rect 12342 7046 12394 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 2320 6987 2372 6996
rect 2320 6953 2329 6987
rect 2329 6953 2363 6987
rect 2363 6953 2372 6987
rect 2320 6944 2372 6953
rect 5724 6987 5776 6996
rect 5724 6953 5754 6987
rect 5754 6953 5776 6987
rect 5724 6944 5776 6953
rect 9496 6944 9548 6996
rect 10968 6987 11020 6996
rect 10968 6953 10977 6987
rect 10977 6953 11011 6987
rect 11011 6953 11020 6987
rect 10968 6944 11020 6953
rect 12900 6944 12952 6996
rect 2412 6919 2464 6928
rect 2412 6885 2421 6919
rect 2421 6885 2455 6919
rect 2455 6885 2464 6919
rect 2412 6876 2464 6885
rect 4528 6876 4580 6928
rect 6736 6876 6788 6928
rect 3976 6808 4028 6860
rect 2044 6740 2096 6792
rect 3148 6740 3200 6792
rect 4620 6808 4672 6860
rect 4896 6808 4948 6860
rect 5172 6808 5224 6860
rect 5448 6851 5500 6860
rect 5448 6817 5457 6851
rect 5457 6817 5491 6851
rect 5491 6817 5500 6851
rect 5448 6808 5500 6817
rect 7748 6808 7800 6860
rect 5264 6740 5316 6792
rect 8392 6876 8444 6928
rect 9036 6876 9088 6928
rect 10232 6876 10284 6928
rect 8024 6851 8076 6860
rect 8024 6817 8033 6851
rect 8033 6817 8067 6851
rect 8067 6817 8076 6851
rect 8024 6808 8076 6817
rect 9404 6808 9456 6860
rect 9956 6808 10008 6860
rect 10324 6808 10376 6860
rect 10876 6876 10928 6928
rect 11520 6919 11572 6928
rect 11520 6885 11529 6919
rect 11529 6885 11563 6919
rect 11563 6885 11572 6919
rect 11520 6876 11572 6885
rect 11336 6808 11388 6860
rect 11612 6851 11664 6860
rect 11612 6817 11621 6851
rect 11621 6817 11655 6851
rect 11655 6817 11664 6851
rect 11612 6808 11664 6817
rect 3884 6647 3936 6656
rect 3884 6613 3885 6647
rect 3885 6613 3919 6647
rect 3919 6613 3936 6647
rect 3884 6604 3936 6613
rect 3976 6604 4028 6656
rect 4068 6604 4120 6656
rect 5172 6672 5224 6724
rect 8760 6740 8812 6792
rect 5632 6672 5684 6724
rect 7012 6672 7064 6724
rect 7932 6672 7984 6724
rect 8668 6672 8720 6724
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 10692 6740 10744 6792
rect 11152 6740 11204 6792
rect 11796 6740 11848 6792
rect 12072 6740 12124 6792
rect 13360 6740 13412 6792
rect 9128 6715 9180 6724
rect 9128 6681 9137 6715
rect 9137 6681 9171 6715
rect 9171 6681 9180 6715
rect 9128 6672 9180 6681
rect 9496 6672 9548 6724
rect 9864 6672 9916 6724
rect 5724 6604 5776 6656
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 7748 6647 7800 6656
rect 7748 6613 7757 6647
rect 7757 6613 7791 6647
rect 7791 6613 7800 6647
rect 7748 6604 7800 6613
rect 8024 6604 8076 6656
rect 8576 6604 8628 6656
rect 8944 6604 8996 6656
rect 9680 6604 9732 6656
rect 10140 6604 10192 6656
rect 11980 6647 12032 6656
rect 11980 6613 11989 6647
rect 11989 6613 12023 6647
rect 12023 6613 12032 6647
rect 11980 6604 12032 6613
rect 12624 6604 12676 6656
rect 8214 6502 8266 6554
rect 8278 6502 8330 6554
rect 8342 6502 8394 6554
rect 8406 6502 8458 6554
rect 8470 6502 8522 6554
rect 2228 6332 2280 6384
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 3608 6307 3660 6316
rect 3608 6273 3617 6307
rect 3617 6273 3651 6307
rect 3651 6273 3660 6307
rect 3608 6264 3660 6273
rect 4896 6443 4948 6452
rect 4896 6409 4905 6443
rect 4905 6409 4939 6443
rect 4939 6409 4948 6443
rect 4896 6400 4948 6409
rect 5080 6400 5132 6452
rect 6000 6443 6052 6452
rect 6000 6409 6009 6443
rect 6009 6409 6043 6443
rect 6043 6409 6052 6443
rect 6000 6400 6052 6409
rect 7472 6400 7524 6452
rect 8852 6443 8904 6452
rect 8852 6409 8861 6443
rect 8861 6409 8895 6443
rect 8895 6409 8904 6443
rect 8852 6400 8904 6409
rect 8944 6400 8996 6452
rect 10324 6400 10376 6452
rect 5724 6375 5776 6384
rect 5724 6341 5733 6375
rect 5733 6341 5767 6375
rect 5767 6341 5776 6375
rect 5724 6332 5776 6341
rect 7104 6332 7156 6384
rect 7748 6332 7800 6384
rect 11980 6400 12032 6452
rect 13268 6443 13320 6452
rect 4160 6264 4212 6316
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 3792 6196 3844 6248
rect 4528 6264 4580 6316
rect 3884 6128 3936 6180
rect 4528 6128 4580 6180
rect 3976 6060 4028 6112
rect 5172 6307 5224 6316
rect 5172 6273 5181 6307
rect 5181 6273 5215 6307
rect 5215 6273 5224 6307
rect 5356 6307 5408 6316
rect 5172 6264 5224 6273
rect 5356 6273 5365 6307
rect 5365 6273 5399 6307
rect 5399 6273 5408 6307
rect 5356 6264 5408 6273
rect 5632 6307 5684 6316
rect 5632 6273 5641 6307
rect 5641 6273 5675 6307
rect 5675 6273 5684 6307
rect 5632 6264 5684 6273
rect 6092 6264 6144 6316
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 6644 6307 6696 6316
rect 6644 6273 6653 6307
rect 6653 6273 6687 6307
rect 6687 6273 6696 6307
rect 6644 6264 6696 6273
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 7196 6264 7248 6316
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 6276 6196 6328 6248
rect 8208 6307 8260 6316
rect 8208 6273 8217 6307
rect 8217 6273 8251 6307
rect 8251 6273 8260 6307
rect 8208 6264 8260 6273
rect 8392 6264 8444 6316
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 11060 6332 11112 6384
rect 12532 6375 12584 6384
rect 12532 6341 12541 6375
rect 12541 6341 12575 6375
rect 12575 6341 12584 6375
rect 12532 6332 12584 6341
rect 13268 6409 13277 6443
rect 13277 6409 13311 6443
rect 13311 6409 13320 6443
rect 13268 6400 13320 6409
rect 8300 6239 8352 6248
rect 8300 6205 8309 6239
rect 8309 6205 8343 6239
rect 8343 6205 8352 6239
rect 8300 6196 8352 6205
rect 8576 6196 8628 6248
rect 5632 6128 5684 6180
rect 6736 6128 6788 6180
rect 7104 6171 7156 6180
rect 7104 6137 7113 6171
rect 7113 6137 7147 6171
rect 7147 6137 7156 6171
rect 7104 6128 7156 6137
rect 7288 6128 7340 6180
rect 7656 6171 7708 6180
rect 7656 6137 7665 6171
rect 7665 6137 7699 6171
rect 7699 6137 7708 6171
rect 7656 6128 7708 6137
rect 8024 6128 8076 6180
rect 9496 6196 9548 6248
rect 10876 6196 10928 6248
rect 9680 6128 9732 6180
rect 10232 6128 10284 6180
rect 11980 6239 12032 6248
rect 11980 6205 11989 6239
rect 11989 6205 12023 6239
rect 12023 6205 12032 6239
rect 11980 6196 12032 6205
rect 13084 6264 13136 6316
rect 13360 6239 13412 6248
rect 13360 6205 13369 6239
rect 13369 6205 13403 6239
rect 13403 6205 13412 6239
rect 13360 6196 13412 6205
rect 12900 6128 12952 6180
rect 5448 6060 5500 6112
rect 8300 6060 8352 6112
rect 9496 6103 9548 6112
rect 9496 6069 9505 6103
rect 9505 6069 9539 6103
rect 9539 6069 9548 6103
rect 9496 6060 9548 6069
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 10048 6060 10100 6069
rect 10876 6060 10928 6112
rect 11888 6060 11940 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 12214 5958 12266 6010
rect 12278 5958 12330 6010
rect 12342 5958 12394 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 2228 5899 2280 5908
rect 2228 5865 2237 5899
rect 2237 5865 2271 5899
rect 2271 5865 2280 5899
rect 2228 5856 2280 5865
rect 4712 5856 4764 5908
rect 4436 5788 4488 5840
rect 5080 5856 5132 5908
rect 6092 5899 6144 5908
rect 6092 5865 6101 5899
rect 6101 5865 6135 5899
rect 6135 5865 6144 5899
rect 6092 5856 6144 5865
rect 6276 5856 6328 5908
rect 7932 5856 7984 5908
rect 8024 5899 8076 5908
rect 8024 5865 8033 5899
rect 8033 5865 8067 5899
rect 8067 5865 8076 5899
rect 8024 5856 8076 5865
rect 5172 5788 5224 5840
rect 5264 5788 5316 5840
rect 3976 5763 4028 5772
rect 3976 5729 3985 5763
rect 3985 5729 4019 5763
rect 4019 5729 4028 5763
rect 3976 5720 4028 5729
rect 2044 5695 2096 5704
rect 2044 5661 2053 5695
rect 2053 5661 2087 5695
rect 2087 5661 2096 5695
rect 2044 5652 2096 5661
rect 3148 5695 3200 5704
rect 3148 5661 3157 5695
rect 3157 5661 3191 5695
rect 3191 5661 3200 5695
rect 3148 5652 3200 5661
rect 3700 5652 3752 5704
rect 4528 5652 4580 5704
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 4988 5695 5040 5704
rect 4988 5661 4997 5695
rect 4997 5661 5031 5695
rect 5031 5661 5040 5695
rect 5448 5695 5500 5704
rect 4988 5652 5040 5661
rect 4620 5584 4672 5636
rect 5448 5661 5497 5695
rect 5497 5661 5500 5695
rect 5448 5652 5500 5661
rect 5356 5584 5408 5636
rect 6092 5720 6144 5772
rect 7288 5788 7340 5840
rect 8300 5856 8352 5908
rect 10508 5899 10560 5908
rect 10508 5865 10517 5899
rect 10517 5865 10551 5899
rect 10551 5865 10560 5899
rect 10508 5856 10560 5865
rect 10692 5899 10744 5908
rect 10692 5865 10701 5899
rect 10701 5865 10735 5899
rect 10735 5865 10744 5899
rect 10692 5856 10744 5865
rect 11704 5856 11756 5908
rect 13268 5856 13320 5908
rect 9680 5788 9732 5840
rect 10232 5788 10284 5840
rect 11152 5788 11204 5840
rect 13360 5788 13412 5840
rect 6460 5652 6512 5704
rect 7656 5720 7708 5772
rect 2872 5516 2924 5568
rect 6184 5584 6236 5636
rect 7840 5695 7892 5704
rect 7840 5661 7849 5695
rect 7849 5661 7883 5695
rect 7883 5661 7892 5695
rect 7840 5652 7892 5661
rect 8760 5720 8812 5772
rect 9588 5720 9640 5772
rect 10784 5720 10836 5772
rect 11244 5720 11296 5772
rect 12072 5720 12124 5772
rect 8116 5584 8168 5636
rect 8392 5584 8444 5636
rect 8668 5652 8720 5704
rect 8944 5695 8996 5704
rect 8944 5661 8953 5695
rect 8953 5661 8987 5695
rect 8987 5661 8996 5695
rect 8944 5652 8996 5661
rect 9036 5584 9088 5636
rect 7196 5516 7248 5568
rect 7472 5516 7524 5568
rect 9312 5652 9364 5704
rect 11060 5652 11112 5704
rect 11888 5695 11940 5704
rect 11888 5661 11897 5695
rect 11897 5661 11931 5695
rect 11931 5661 11940 5695
rect 11888 5652 11940 5661
rect 12532 5695 12584 5704
rect 12532 5661 12541 5695
rect 12541 5661 12575 5695
rect 12575 5661 12584 5695
rect 12532 5652 12584 5661
rect 10876 5584 10928 5636
rect 12992 5627 13044 5636
rect 12992 5593 13001 5627
rect 13001 5593 13035 5627
rect 13035 5593 13044 5627
rect 12992 5584 13044 5593
rect 10048 5559 10100 5568
rect 10048 5525 10057 5559
rect 10057 5525 10091 5559
rect 10091 5525 10100 5559
rect 10048 5516 10100 5525
rect 10140 5559 10192 5568
rect 10140 5525 10149 5559
rect 10149 5525 10183 5559
rect 10183 5525 10192 5559
rect 10140 5516 10192 5525
rect 10784 5516 10836 5568
rect 13176 5559 13228 5568
rect 13176 5525 13185 5559
rect 13185 5525 13219 5559
rect 13219 5525 13228 5559
rect 13176 5516 13228 5525
rect 8214 5414 8266 5466
rect 8278 5414 8330 5466
rect 8342 5414 8394 5466
rect 8406 5414 8458 5466
rect 8470 5414 8522 5466
rect 3148 5355 3200 5364
rect 3148 5321 3157 5355
rect 3157 5321 3191 5355
rect 3191 5321 3200 5355
rect 3148 5312 3200 5321
rect 2228 5244 2280 5296
rect 3516 5244 3568 5296
rect 8668 5312 8720 5364
rect 10140 5355 10192 5364
rect 5632 5287 5684 5296
rect 5632 5253 5641 5287
rect 5641 5253 5675 5287
rect 5675 5253 5684 5287
rect 5632 5244 5684 5253
rect 6184 5244 6236 5296
rect 6552 5244 6604 5296
rect 6828 5244 6880 5296
rect 7288 5287 7340 5296
rect 2964 5176 3016 5228
rect 3792 5219 3844 5228
rect 3792 5185 3801 5219
rect 3801 5185 3835 5219
rect 3835 5185 3844 5219
rect 3792 5176 3844 5185
rect 3884 5219 3936 5228
rect 3884 5185 3893 5219
rect 3893 5185 3927 5219
rect 3927 5185 3936 5219
rect 3884 5176 3936 5185
rect 4068 5176 4120 5228
rect 4436 5219 4488 5228
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 2412 5108 2464 5160
rect 4436 5185 4445 5219
rect 4445 5185 4479 5219
rect 4479 5185 4488 5219
rect 4436 5176 4488 5185
rect 4712 5176 4764 5228
rect 4896 5176 4948 5228
rect 5264 5219 5316 5228
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 4620 5040 4672 5092
rect 3700 4972 3752 5024
rect 3792 4972 3844 5024
rect 5540 5151 5592 5160
rect 5540 5117 5549 5151
rect 5549 5117 5583 5151
rect 5583 5117 5592 5151
rect 5540 5108 5592 5117
rect 6736 5219 6788 5228
rect 6736 5185 6745 5219
rect 6745 5185 6779 5219
rect 6779 5185 6788 5219
rect 7288 5253 7297 5287
rect 7297 5253 7331 5287
rect 7331 5253 7340 5287
rect 7288 5244 7340 5253
rect 7840 5244 7892 5296
rect 6736 5176 6788 5185
rect 8576 5244 8628 5296
rect 9312 5244 9364 5296
rect 5724 4972 5776 5024
rect 6184 5040 6236 5092
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 8944 5176 8996 5228
rect 10140 5321 10149 5355
rect 10149 5321 10183 5355
rect 10183 5321 10192 5355
rect 10140 5312 10192 5321
rect 10968 5355 11020 5364
rect 10968 5321 10977 5355
rect 10977 5321 11011 5355
rect 11011 5321 11020 5355
rect 10968 5312 11020 5321
rect 11520 5287 11572 5296
rect 11520 5253 11529 5287
rect 11529 5253 11563 5287
rect 11563 5253 11572 5287
rect 11520 5244 11572 5253
rect 11980 5312 12032 5364
rect 10508 5219 10560 5228
rect 9588 5108 9640 5160
rect 10508 5185 10517 5219
rect 10517 5185 10551 5219
rect 10551 5185 10560 5219
rect 10508 5176 10560 5185
rect 10692 5176 10744 5228
rect 11060 5176 11112 5228
rect 11428 5108 11480 5160
rect 7564 5040 7616 5092
rect 8116 5040 8168 5092
rect 6460 5015 6512 5024
rect 6460 4981 6469 5015
rect 6469 4981 6503 5015
rect 6503 4981 6512 5015
rect 6460 4972 6512 4981
rect 8392 5015 8444 5024
rect 8392 4981 8401 5015
rect 8401 4981 8435 5015
rect 8435 4981 8444 5015
rect 8392 4972 8444 4981
rect 10232 5040 10284 5092
rect 10416 5083 10468 5092
rect 10416 5049 10425 5083
rect 10425 5049 10459 5083
rect 10459 5049 10468 5083
rect 10416 5040 10468 5049
rect 10692 5040 10744 5092
rect 10784 5040 10836 5092
rect 12532 5176 12584 5228
rect 12900 5219 12952 5228
rect 12900 5185 12909 5219
rect 12909 5185 12943 5219
rect 12943 5185 12952 5219
rect 12900 5176 12952 5185
rect 9864 4972 9916 5024
rect 10140 4972 10192 5024
rect 12992 5040 13044 5092
rect 11060 4972 11112 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 12214 4870 12266 4922
rect 12278 4870 12330 4922
rect 12342 4870 12394 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 2228 4811 2280 4820
rect 2228 4777 2237 4811
rect 2237 4777 2271 4811
rect 2271 4777 2280 4811
rect 2228 4768 2280 4777
rect 2412 4768 2464 4820
rect 3516 4768 3568 4820
rect 4620 4768 4672 4820
rect 6184 4811 6236 4820
rect 6184 4777 6193 4811
rect 6193 4777 6227 4811
rect 6227 4777 6236 4811
rect 6184 4768 6236 4777
rect 7288 4768 7340 4820
rect 9864 4768 9916 4820
rect 10508 4768 10560 4820
rect 10784 4811 10836 4820
rect 10784 4777 10793 4811
rect 10793 4777 10827 4811
rect 10827 4777 10836 4811
rect 10784 4768 10836 4777
rect 13360 4811 13412 4820
rect 13360 4777 13369 4811
rect 13369 4777 13403 4811
rect 13403 4777 13412 4811
rect 13360 4768 13412 4777
rect 2044 4607 2096 4616
rect 2044 4573 2053 4607
rect 2053 4573 2087 4607
rect 2087 4573 2096 4607
rect 2044 4564 2096 4573
rect 2504 4564 2556 4616
rect 2872 4632 2924 4684
rect 3148 4632 3200 4684
rect 2964 4564 3016 4616
rect 3700 4632 3752 4684
rect 8760 4743 8812 4752
rect 8760 4709 8769 4743
rect 8769 4709 8803 4743
rect 8803 4709 8812 4743
rect 8760 4700 8812 4709
rect 4436 4632 4488 4684
rect 4804 4632 4856 4684
rect 5356 4632 5408 4684
rect 5540 4675 5592 4684
rect 5540 4641 5549 4675
rect 5549 4641 5583 4675
rect 5583 4641 5592 4675
rect 5540 4632 5592 4641
rect 4068 4564 4120 4616
rect 5632 4564 5684 4616
rect 3240 4539 3292 4548
rect 3240 4505 3249 4539
rect 3249 4505 3283 4539
rect 3283 4505 3292 4539
rect 3240 4496 3292 4505
rect 4436 4496 4488 4548
rect 4804 4539 4856 4548
rect 4804 4505 4813 4539
rect 4813 4505 4847 4539
rect 4847 4505 4856 4539
rect 4804 4496 4856 4505
rect 4988 4539 5040 4548
rect 4988 4505 4997 4539
rect 4997 4505 5031 4539
rect 5031 4505 5040 4539
rect 4988 4496 5040 4505
rect 5080 4496 5132 4548
rect 5540 4496 5592 4548
rect 6828 4607 6880 4616
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 7196 4607 7248 4616
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7196 4564 7248 4573
rect 8024 4632 8076 4684
rect 8944 4632 8996 4684
rect 7472 4607 7524 4616
rect 7472 4573 7481 4607
rect 7481 4573 7515 4607
rect 7515 4573 7524 4607
rect 7472 4564 7524 4573
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 8576 4607 8628 4616
rect 8576 4573 8585 4607
rect 8585 4573 8619 4607
rect 8619 4573 8628 4607
rect 8576 4564 8628 4573
rect 9312 4607 9364 4616
rect 9312 4573 9321 4607
rect 9321 4573 9355 4607
rect 9355 4573 9364 4607
rect 9312 4564 9364 4573
rect 10416 4675 10468 4684
rect 10416 4641 10425 4675
rect 10425 4641 10459 4675
rect 10459 4641 10468 4675
rect 10416 4632 10468 4641
rect 9956 4607 10008 4616
rect 9956 4573 9965 4607
rect 9965 4573 9999 4607
rect 9999 4573 10008 4607
rect 9956 4564 10008 4573
rect 10140 4607 10192 4616
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 10232 4564 10284 4616
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 13176 4700 13228 4752
rect 4528 4428 4580 4480
rect 7840 4496 7892 4548
rect 7564 4471 7616 4480
rect 7564 4437 7573 4471
rect 7573 4437 7607 4471
rect 7607 4437 7616 4471
rect 7564 4428 7616 4437
rect 8668 4428 8720 4480
rect 10416 4496 10468 4548
rect 11520 4564 11572 4616
rect 12900 4607 12952 4616
rect 12900 4573 12909 4607
rect 12909 4573 12943 4607
rect 12943 4573 12952 4607
rect 12900 4564 12952 4573
rect 12992 4564 13044 4616
rect 10692 4496 10744 4548
rect 10048 4428 10100 4480
rect 13268 4428 13320 4480
rect 8214 4326 8266 4378
rect 8278 4326 8330 4378
rect 8342 4326 8394 4378
rect 8406 4326 8458 4378
rect 8470 4326 8522 4378
rect 3516 4267 3568 4276
rect 3516 4233 3525 4267
rect 3525 4233 3559 4267
rect 3559 4233 3568 4267
rect 3516 4224 3568 4233
rect 2412 4156 2464 4208
rect 2964 4156 3016 4208
rect 4988 4224 5040 4276
rect 4528 4199 4580 4208
rect 3240 4088 3292 4140
rect 4528 4165 4537 4199
rect 4537 4165 4571 4199
rect 4571 4165 4580 4199
rect 4528 4156 4580 4165
rect 4712 4156 4764 4208
rect 4436 4131 4488 4140
rect 1400 4063 1452 4072
rect 1400 4029 1409 4063
rect 1409 4029 1443 4063
rect 1443 4029 1452 4063
rect 1400 4020 1452 4029
rect 3424 4063 3476 4072
rect 3424 4029 3433 4063
rect 3433 4029 3467 4063
rect 3467 4029 3476 4063
rect 3424 4020 3476 4029
rect 4436 4097 4440 4131
rect 4440 4097 4474 4131
rect 4474 4097 4488 4131
rect 4436 4088 4488 4097
rect 4896 4088 4948 4140
rect 5908 4088 5960 4140
rect 6460 4224 6512 4276
rect 6920 4224 6972 4276
rect 11796 4224 11848 4276
rect 8024 4156 8076 4208
rect 9312 4156 9364 4208
rect 10140 4156 10192 4208
rect 6368 4131 6420 4140
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 7012 4088 7064 4140
rect 7380 4088 7432 4140
rect 7840 4131 7892 4140
rect 7840 4097 7849 4131
rect 7849 4097 7883 4131
rect 7883 4097 7892 4131
rect 7840 4088 7892 4097
rect 9220 4131 9272 4140
rect 9220 4097 9229 4131
rect 9229 4097 9263 4131
rect 9263 4097 9272 4131
rect 9220 4088 9272 4097
rect 9956 4131 10008 4140
rect 8300 4020 8352 4072
rect 9128 4020 9180 4072
rect 6828 3952 6880 4004
rect 8852 3952 8904 4004
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 10048 4131 10100 4140
rect 10048 4097 10057 4131
rect 10057 4097 10091 4131
rect 10091 4097 10100 4131
rect 10048 4088 10100 4097
rect 10232 4131 10284 4140
rect 10232 4097 10241 4131
rect 10241 4097 10275 4131
rect 10275 4097 10284 4131
rect 10692 4199 10744 4208
rect 10232 4088 10284 4097
rect 10692 4165 10701 4199
rect 10701 4165 10735 4199
rect 10735 4165 10744 4199
rect 10692 4156 10744 4165
rect 11060 4156 11112 4208
rect 11520 4156 11572 4208
rect 13268 4131 13320 4140
rect 4068 3884 4120 3936
rect 5540 3884 5592 3936
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 7472 3884 7524 3936
rect 8576 3884 8628 3936
rect 8668 3884 8720 3936
rect 8944 3884 8996 3936
rect 9864 3884 9916 3936
rect 10416 3952 10468 4004
rect 10784 3952 10836 4004
rect 11520 4020 11572 4072
rect 11980 4020 12032 4072
rect 12992 4063 13044 4072
rect 12992 4029 13001 4063
rect 13001 4029 13035 4063
rect 13035 4029 13044 4063
rect 12992 4020 13044 4029
rect 11704 3952 11756 4004
rect 12900 3995 12952 4004
rect 12900 3961 12909 3995
rect 12909 3961 12943 3995
rect 12943 3961 12952 3995
rect 12900 3952 12952 3961
rect 13268 4097 13277 4131
rect 13277 4097 13311 4131
rect 13311 4097 13320 4131
rect 13268 4088 13320 4097
rect 11060 3884 11112 3936
rect 11888 3884 11940 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 12214 3782 12266 3834
rect 12278 3782 12330 3834
rect 12342 3782 12394 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 2412 3723 2464 3732
rect 2412 3689 2421 3723
rect 2421 3689 2455 3723
rect 2455 3689 2464 3723
rect 2412 3680 2464 3689
rect 2964 3680 3016 3732
rect 3424 3680 3476 3732
rect 5908 3723 5960 3732
rect 5908 3689 5917 3723
rect 5917 3689 5951 3723
rect 5951 3689 5960 3723
rect 5908 3680 5960 3689
rect 6368 3680 6420 3732
rect 7656 3680 7708 3732
rect 9404 3723 9456 3732
rect 5172 3655 5224 3664
rect 5172 3621 5181 3655
rect 5181 3621 5215 3655
rect 5215 3621 5224 3655
rect 5172 3612 5224 3621
rect 6000 3612 6052 3664
rect 4620 3544 4672 3596
rect 7012 3587 7064 3596
rect 7012 3553 7021 3587
rect 7021 3553 7055 3587
rect 7055 3553 7064 3587
rect 7012 3544 7064 3553
rect 8300 3612 8352 3664
rect 1584 3476 1636 3528
rect 2504 3476 2556 3528
rect 3516 3476 3568 3528
rect 4068 3476 4120 3528
rect 5080 3476 5132 3528
rect 3700 3408 3752 3460
rect 5816 3476 5868 3528
rect 6644 3476 6696 3528
rect 7472 3476 7524 3528
rect 7840 3519 7892 3528
rect 7840 3485 7849 3519
rect 7849 3485 7883 3519
rect 7883 3485 7892 3519
rect 7840 3476 7892 3485
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 6828 3408 6880 3460
rect 9404 3689 9413 3723
rect 9413 3689 9447 3723
rect 9447 3689 9456 3723
rect 9404 3680 9456 3689
rect 9956 3612 10008 3664
rect 10508 3612 10560 3664
rect 10968 3612 11020 3664
rect 12900 3612 12952 3664
rect 8576 3476 8628 3528
rect 8760 3519 8812 3528
rect 8760 3485 8769 3519
rect 8769 3485 8803 3519
rect 8803 3485 8812 3519
rect 8760 3476 8812 3485
rect 9036 3476 9088 3528
rect 9772 3470 9824 3522
rect 7472 3340 7524 3392
rect 7656 3383 7708 3392
rect 7656 3349 7665 3383
rect 7665 3349 7699 3383
rect 7699 3349 7708 3383
rect 7656 3340 7708 3349
rect 7932 3383 7984 3392
rect 7932 3349 7941 3383
rect 7941 3349 7975 3383
rect 7975 3349 7984 3383
rect 7932 3340 7984 3349
rect 8116 3340 8168 3392
rect 11520 3476 11572 3528
rect 11980 3519 12032 3528
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 8852 3340 8904 3392
rect 8944 3383 8996 3392
rect 8944 3349 8953 3383
rect 8953 3349 8987 3383
rect 8987 3349 8996 3383
rect 8944 3340 8996 3349
rect 9404 3340 9456 3392
rect 11060 3408 11112 3460
rect 11428 3408 11480 3460
rect 11704 3451 11756 3460
rect 11704 3417 11713 3451
rect 11713 3417 11747 3451
rect 11747 3417 11756 3451
rect 11704 3408 11756 3417
rect 13268 3476 13320 3528
rect 10048 3340 10100 3392
rect 10232 3383 10284 3392
rect 10232 3349 10241 3383
rect 10241 3349 10275 3383
rect 10275 3349 10284 3383
rect 10232 3340 10284 3349
rect 8214 3238 8266 3290
rect 8278 3238 8330 3290
rect 8342 3238 8394 3290
rect 8406 3238 8458 3290
rect 8470 3238 8522 3290
rect 3332 3136 3384 3188
rect 4804 3136 4856 3188
rect 5356 3179 5408 3188
rect 5356 3145 5365 3179
rect 5365 3145 5399 3179
rect 5399 3145 5408 3179
rect 5356 3136 5408 3145
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 2872 3000 2924 3052
rect 4620 3068 4672 3120
rect 5816 3043 5868 3052
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 5816 3000 5868 3009
rect 7012 3136 7064 3188
rect 8116 3136 8168 3188
rect 9588 3136 9640 3188
rect 10232 3136 10284 3188
rect 11980 3136 12032 3188
rect 12992 3136 13044 3188
rect 7472 3068 7524 3120
rect 7932 3068 7984 3120
rect 7840 3000 7892 3052
rect 8116 3000 8168 3052
rect 9220 3043 9272 3052
rect 9220 3009 9229 3043
rect 9229 3009 9263 3043
rect 9263 3009 9272 3043
rect 9220 3000 9272 3009
rect 9404 3043 9456 3052
rect 9404 3009 9413 3043
rect 9413 3009 9447 3043
rect 9447 3009 9456 3043
rect 9404 3000 9456 3009
rect 3424 2975 3476 2984
rect 3424 2941 3433 2975
rect 3433 2941 3467 2975
rect 3467 2941 3476 2975
rect 3424 2932 3476 2941
rect 1584 2864 1636 2916
rect 5264 2932 5316 2984
rect 8944 2932 8996 2984
rect 9680 2932 9732 2984
rect 10416 3000 10468 3052
rect 10692 3043 10744 3052
rect 10692 3009 10701 3043
rect 10701 3009 10735 3043
rect 10735 3009 10744 3043
rect 10692 3000 10744 3009
rect 11060 3043 11112 3052
rect 11060 3009 11069 3043
rect 11069 3009 11103 3043
rect 11103 3009 11112 3043
rect 11060 3000 11112 3009
rect 11704 3068 11756 3120
rect 4988 2864 5040 2916
rect 9956 2864 10008 2916
rect 10508 2864 10560 2916
rect 10968 2864 11020 2916
rect 11060 2864 11112 2916
rect 11888 2932 11940 2984
rect 12072 2975 12124 2984
rect 12072 2941 12081 2975
rect 12081 2941 12115 2975
rect 12115 2941 12124 2975
rect 12072 2932 12124 2941
rect 11520 2907 11572 2916
rect 11520 2873 11529 2907
rect 11529 2873 11563 2907
rect 11563 2873 11572 2907
rect 11520 2864 11572 2873
rect 2596 2796 2648 2848
rect 5908 2796 5960 2848
rect 6184 2796 6236 2848
rect 10600 2796 10652 2848
rect 12072 2796 12124 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 12214 2694 12266 2746
rect 12278 2694 12330 2746
rect 12342 2694 12394 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 3424 2592 3476 2644
rect 4620 2635 4672 2644
rect 4620 2601 4629 2635
rect 4629 2601 4663 2635
rect 4663 2601 4672 2635
rect 4620 2592 4672 2601
rect 6644 2635 6696 2644
rect 6644 2601 6653 2635
rect 6653 2601 6687 2635
rect 6687 2601 6696 2635
rect 6644 2592 6696 2601
rect 9588 2592 9640 2644
rect 10508 2635 10560 2644
rect 10508 2601 10517 2635
rect 10517 2601 10551 2635
rect 10551 2601 10560 2635
rect 10508 2592 10560 2601
rect 11244 2592 11296 2644
rect 7472 2567 7524 2576
rect 7472 2533 7481 2567
rect 7481 2533 7515 2567
rect 7515 2533 7524 2567
rect 7472 2524 7524 2533
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 2872 2456 2924 2508
rect 5172 2499 5224 2508
rect 5172 2465 5181 2499
rect 5181 2465 5215 2499
rect 5215 2465 5224 2499
rect 5172 2456 5224 2465
rect 7012 2499 7064 2508
rect 7012 2465 7021 2499
rect 7021 2465 7055 2499
rect 7055 2465 7064 2499
rect 7012 2456 7064 2465
rect 7656 2524 7708 2576
rect 8116 2567 8168 2576
rect 8116 2533 8125 2567
rect 8125 2533 8159 2567
rect 8159 2533 8168 2567
rect 8116 2524 8168 2533
rect 9496 2524 9548 2576
rect 10876 2524 10928 2576
rect 9680 2456 9732 2508
rect 10600 2456 10652 2508
rect 11244 2456 11296 2508
rect 11980 2499 12032 2508
rect 11980 2465 11989 2499
rect 11989 2465 12023 2499
rect 12023 2465 12032 2499
rect 11980 2456 12032 2465
rect 2596 2320 2648 2372
rect 4620 2252 4672 2304
rect 7748 2388 7800 2440
rect 8944 2388 8996 2440
rect 11060 2388 11112 2440
rect 11336 2388 11388 2440
rect 11428 2388 11480 2440
rect 5264 2320 5316 2372
rect 5908 2320 5960 2372
rect 5816 2252 5868 2304
rect 6460 2252 6512 2304
rect 8576 2320 8628 2372
rect 9312 2363 9364 2372
rect 9312 2329 9321 2363
rect 9321 2329 9355 2363
rect 9355 2329 9364 2363
rect 9312 2320 9364 2329
rect 9864 2320 9916 2372
rect 10784 2363 10836 2372
rect 9588 2295 9640 2304
rect 9588 2261 9597 2295
rect 9597 2261 9631 2295
rect 9631 2261 9640 2295
rect 9588 2252 9640 2261
rect 9772 2252 9824 2304
rect 10784 2329 10793 2363
rect 10793 2329 10827 2363
rect 10827 2329 10836 2363
rect 10784 2320 10836 2329
rect 11612 2363 11664 2372
rect 11612 2329 11621 2363
rect 11621 2329 11655 2363
rect 11655 2329 11664 2363
rect 11612 2320 11664 2329
rect 13084 2320 13136 2372
rect 11152 2252 11204 2304
rect 12072 2252 12124 2304
rect 12624 2295 12676 2304
rect 12624 2261 12633 2295
rect 12633 2261 12667 2295
rect 12667 2261 12676 2295
rect 12624 2252 12676 2261
rect 13268 2363 13320 2372
rect 13268 2329 13277 2363
rect 13277 2329 13311 2363
rect 13311 2329 13320 2363
rect 13268 2320 13320 2329
rect 8214 2150 8266 2202
rect 8278 2150 8330 2202
rect 8342 2150 8394 2202
rect 8406 2150 8458 2202
rect 8470 2150 8522 2202
rect 5724 2048 5776 2100
rect 1584 1980 1636 2032
rect 2228 1980 2280 2032
rect 3424 1980 3476 2032
rect 7748 2048 7800 2100
rect 8944 2091 8996 2100
rect 8944 2057 8953 2091
rect 8953 2057 8987 2091
rect 8987 2057 8996 2091
rect 8944 2048 8996 2057
rect 10048 2048 10100 2100
rect 11336 2091 11388 2100
rect 11336 2057 11345 2091
rect 11345 2057 11379 2091
rect 11379 2057 11388 2091
rect 11336 2048 11388 2057
rect 5264 1912 5316 1964
rect 5448 1955 5500 1964
rect 5448 1921 5487 1955
rect 5487 1921 5500 1955
rect 6000 1955 6052 1964
rect 5448 1912 5500 1921
rect 6000 1921 6009 1955
rect 6009 1921 6043 1955
rect 6043 1921 6052 1955
rect 6000 1912 6052 1921
rect 6460 1955 6512 1964
rect 6460 1921 6469 1955
rect 6469 1921 6503 1955
rect 6503 1921 6512 1955
rect 6460 1912 6512 1921
rect 3056 1844 3108 1896
rect 7564 1912 7616 1964
rect 9588 1912 9640 1964
rect 9864 1980 9916 2032
rect 10324 1980 10376 2032
rect 12900 1980 12952 2032
rect 2872 1776 2924 1828
rect 940 1708 992 1760
rect 5724 1776 5776 1828
rect 8576 1819 8628 1828
rect 8576 1785 8585 1819
rect 8585 1785 8619 1819
rect 8619 1785 8628 1819
rect 8576 1776 8628 1785
rect 10600 1844 10652 1896
rect 10876 1887 10928 1896
rect 10876 1853 10885 1887
rect 10885 1853 10919 1887
rect 10919 1853 10928 1887
rect 10876 1844 10928 1853
rect 13360 1844 13412 1896
rect 11612 1776 11664 1828
rect 5356 1751 5408 1760
rect 5356 1717 5365 1751
rect 5365 1717 5399 1751
rect 5399 1717 5408 1751
rect 5356 1708 5408 1717
rect 7012 1751 7064 1760
rect 7012 1717 7021 1751
rect 7021 1717 7055 1751
rect 7055 1717 7064 1751
rect 7012 1708 7064 1717
rect 10324 1751 10376 1760
rect 10324 1717 10333 1751
rect 10333 1717 10367 1751
rect 10367 1717 10376 1751
rect 10324 1708 10376 1717
rect 4214 1606 4266 1658
rect 4278 1606 4330 1658
rect 4342 1606 4394 1658
rect 4406 1606 4458 1658
rect 4470 1606 4522 1658
rect 12214 1606 12266 1658
rect 12278 1606 12330 1658
rect 12342 1606 12394 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 2228 1547 2280 1556
rect 2228 1513 2237 1547
rect 2237 1513 2271 1547
rect 2271 1513 2280 1547
rect 2228 1504 2280 1513
rect 3424 1547 3476 1556
rect 3424 1513 3433 1547
rect 3433 1513 3467 1547
rect 3467 1513 3476 1547
rect 3424 1504 3476 1513
rect 2504 1300 2556 1352
rect 5816 1504 5868 1556
rect 6552 1504 6604 1556
rect 9496 1504 9548 1556
rect 7564 1479 7616 1488
rect 7564 1445 7573 1479
rect 7573 1445 7607 1479
rect 7607 1445 7616 1479
rect 7564 1436 7616 1445
rect 8576 1479 8628 1488
rect 8576 1445 8585 1479
rect 8585 1445 8619 1479
rect 8619 1445 8628 1479
rect 8576 1436 8628 1445
rect 5356 1411 5408 1420
rect 5356 1377 5365 1411
rect 5365 1377 5399 1411
rect 5399 1377 5408 1411
rect 5356 1368 5408 1377
rect 5816 1411 5868 1420
rect 5816 1377 5825 1411
rect 5825 1377 5859 1411
rect 5859 1377 5868 1411
rect 5816 1368 5868 1377
rect 9312 1368 9364 1420
rect 10600 1504 10652 1556
rect 13268 1504 13320 1556
rect 9864 1436 9916 1488
rect 10324 1411 10376 1420
rect 10324 1377 10333 1411
rect 10333 1377 10367 1411
rect 10367 1377 10376 1411
rect 10324 1368 10376 1377
rect 11060 1368 11112 1420
rect 14004 1368 14056 1420
rect 6184 1343 6236 1352
rect 2780 1232 2832 1284
rect 3056 1232 3108 1284
rect 4620 1232 4672 1284
rect 5264 1232 5316 1284
rect 6184 1309 6193 1343
rect 6193 1309 6227 1343
rect 6227 1309 6236 1343
rect 6184 1300 6236 1309
rect 7012 1343 7064 1352
rect 7012 1309 7021 1343
rect 7021 1309 7055 1343
rect 7055 1309 7064 1343
rect 7012 1300 7064 1309
rect 7748 1343 7800 1352
rect 7748 1309 7757 1343
rect 7757 1309 7791 1343
rect 7791 1309 7800 1343
rect 7748 1300 7800 1309
rect 5448 1164 5500 1216
rect 9588 1300 9640 1352
rect 10692 1343 10744 1352
rect 9956 1232 10008 1284
rect 10692 1309 10701 1343
rect 10701 1309 10735 1343
rect 10735 1309 10744 1343
rect 10692 1300 10744 1309
rect 10876 1300 10928 1352
rect 11704 1343 11756 1352
rect 11704 1309 11713 1343
rect 11713 1309 11747 1343
rect 11747 1309 11756 1343
rect 11704 1300 11756 1309
rect 12624 1300 12676 1352
rect 13084 1343 13136 1352
rect 13084 1309 13093 1343
rect 13093 1309 13127 1343
rect 13127 1309 13136 1343
rect 13084 1300 13136 1309
rect 13360 1300 13412 1352
rect 8214 1062 8266 1114
rect 8278 1062 8330 1114
rect 8342 1062 8394 1114
rect 8406 1062 8458 1114
rect 8470 1062 8522 1114
rect 13912 484 13964 536
<< metal2 >>
rect 754 14200 810 15000
rect 2226 14200 2282 15000
rect 3698 14200 3754 15000
rect 5170 14200 5226 15000
rect 6734 14200 6790 15000
rect 8206 14200 8262 15000
rect 9678 14200 9734 15000
rect 10874 14512 10930 14521
rect 10874 14447 10930 14456
rect 768 11014 796 14200
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1492 12164 1544 12170
rect 1492 12106 1544 12112
rect 1504 11257 1532 12106
rect 1872 11898 1900 12718
rect 1860 11892 1912 11898
rect 1860 11834 1912 11840
rect 1490 11248 1546 11257
rect 1490 11183 1546 11192
rect 756 11008 808 11014
rect 756 10950 808 10956
rect 2056 10674 2084 13262
rect 2240 11234 2268 14200
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2596 13184 2648 13190
rect 2596 13126 2648 13132
rect 2608 12918 2636 13126
rect 2596 12912 2648 12918
rect 2596 12854 2648 12860
rect 2700 12374 2728 13262
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 2872 12300 2924 12306
rect 2792 12260 2872 12288
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2240 11206 2360 11234
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2240 10810 2268 11018
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1504 10266 1532 10542
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 2056 9586 2084 10610
rect 2332 10538 2360 11206
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2608 10985 2636 11154
rect 2594 10976 2650 10985
rect 2594 10911 2650 10920
rect 2608 10742 2636 10911
rect 2596 10736 2648 10742
rect 2700 10713 2728 12174
rect 2792 11762 2820 12260
rect 2872 12242 2924 12248
rect 2976 11762 3004 12310
rect 3160 12238 3188 13466
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3148 12232 3200 12238
rect 3068 12192 3148 12220
rect 3068 11830 3096 12192
rect 3148 12174 3200 12180
rect 3344 12220 3372 13262
rect 3608 13184 3660 13190
rect 3608 13126 3660 13132
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3528 12646 3556 12718
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3424 12232 3476 12238
rect 3344 12192 3424 12220
rect 3240 12164 3292 12170
rect 3240 12106 3292 12112
rect 3056 11824 3108 11830
rect 3056 11766 3108 11772
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 3068 11336 3096 11766
rect 3148 11348 3200 11354
rect 3068 11308 3148 11336
rect 3148 11290 3200 11296
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2596 10678 2648 10684
rect 2686 10704 2742 10713
rect 2412 10668 2464 10674
rect 2686 10639 2742 10648
rect 2412 10610 2464 10616
rect 2320 10532 2372 10538
rect 2320 10474 2372 10480
rect 2424 10441 2452 10610
rect 2410 10432 2466 10441
rect 2410 10367 2466 10376
rect 2792 10266 2820 10950
rect 2976 10810 3004 11018
rect 3054 10840 3110 10849
rect 2964 10804 3016 10810
rect 3054 10775 3110 10784
rect 2964 10746 3016 10752
rect 2870 10704 2926 10713
rect 2870 10639 2872 10648
rect 2924 10639 2926 10648
rect 2872 10610 2924 10616
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 2240 9722 2268 9930
rect 2228 9716 2280 9722
rect 2228 9658 2280 9664
rect 2884 9654 2912 10610
rect 3068 10606 3096 10775
rect 3160 10674 3188 11290
rect 3252 11132 3280 12106
rect 3344 11694 3372 12192
rect 3424 12174 3476 12180
rect 3528 12170 3556 12582
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3332 11280 3384 11286
rect 3528 11268 3556 12106
rect 3620 11898 3648 13126
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3384 11240 3556 11268
rect 3332 11222 3384 11228
rect 3332 11144 3384 11150
rect 3252 11104 3332 11132
rect 3252 10985 3280 11104
rect 3332 11086 3384 11092
rect 3332 11008 3384 11014
rect 3238 10976 3294 10985
rect 3332 10950 3384 10956
rect 3238 10911 3294 10920
rect 3344 10674 3372 10950
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3344 10520 3372 10610
rect 3160 10492 3372 10520
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2976 10130 3004 10406
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 3160 9586 3188 10492
rect 3436 10130 3464 11240
rect 3712 11200 3740 14200
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4632 12918 4660 13126
rect 3976 12912 4028 12918
rect 4620 12912 4672 12918
rect 4028 12872 4108 12900
rect 3976 12854 4028 12860
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3528 11172 3740 11200
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1412 7886 1440 8910
rect 2056 8498 2084 9522
rect 3160 9110 3188 9522
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2424 8634 2452 8842
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 3252 8498 3280 9590
rect 3436 9518 3464 10066
rect 3528 9926 3556 11172
rect 3804 11150 3832 12038
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3896 11150 3924 11698
rect 3988 11354 4016 12718
rect 4080 12238 4108 12872
rect 4620 12854 4672 12860
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4436 12164 4488 12170
rect 4436 12106 4488 12112
rect 4342 11792 4398 11801
rect 4342 11727 4344 11736
rect 4396 11727 4398 11736
rect 4344 11698 4396 11704
rect 4448 11626 4476 12106
rect 4540 11812 4568 12242
rect 4620 11824 4672 11830
rect 4540 11784 4620 11812
rect 4620 11766 4672 11772
rect 4710 11792 4766 11801
rect 4710 11727 4766 11736
rect 4804 11756 4856 11762
rect 4436 11620 4488 11626
rect 4436 11562 4488 11568
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 4724 11234 4752 11727
rect 4908 11744 4936 12718
rect 4856 11716 4936 11744
rect 4804 11698 4856 11704
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4540 11206 4752 11234
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4080 10810 4108 11086
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4264 10810 4292 10950
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 3792 10736 3844 10742
rect 3976 10736 4028 10742
rect 3844 10696 3924 10724
rect 3792 10678 3844 10684
rect 3609 10668 3661 10674
rect 3609 10610 3661 10616
rect 3620 10470 3648 10610
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3608 10464 3660 10470
rect 3804 10441 3832 10542
rect 3608 10406 3660 10412
rect 3790 10432 3846 10441
rect 3620 10062 3648 10406
rect 3790 10367 3846 10376
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3620 9586 3648 9998
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3804 8974 3832 10367
rect 3896 10198 3924 10696
rect 3976 10678 4028 10684
rect 3884 10192 3936 10198
rect 3884 10134 3936 10140
rect 3988 10062 4016 10678
rect 4356 10606 4384 11154
rect 4540 10713 4568 11206
rect 4908 11150 4936 11716
rect 5184 11626 5212 14200
rect 6748 13462 6776 14200
rect 8220 13530 8248 14200
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 7668 13382 7880 13410
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 7380 13320 7432 13326
rect 7668 13308 7696 13382
rect 7852 13326 7880 13382
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7432 13280 7696 13308
rect 7748 13320 7800 13326
rect 7380 13262 7432 13268
rect 7748 13262 7800 13268
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5368 11762 5396 12582
rect 5644 11801 5672 12786
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5736 12102 5764 12718
rect 6104 12238 6132 13262
rect 6932 12918 6960 13262
rect 7392 12986 7420 13262
rect 7760 13190 7788 13262
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7116 12442 7144 12854
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7392 12238 7420 12922
rect 7760 12306 7788 13126
rect 7944 12306 7972 13330
rect 8024 13184 8076 13190
rect 8220 13172 8248 13466
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8024 13126 8076 13132
rect 8128 13144 8248 13172
rect 8036 12782 8064 13126
rect 8128 12986 8156 13144
rect 8214 13084 8522 13104
rect 8214 13082 8220 13084
rect 8276 13082 8300 13084
rect 8356 13082 8380 13084
rect 8436 13082 8460 13084
rect 8516 13082 8522 13084
rect 8276 13030 8278 13082
rect 8458 13030 8460 13082
rect 8214 13028 8220 13030
rect 8276 13028 8300 13030
rect 8356 13028 8380 13030
rect 8436 13028 8460 13030
rect 8516 13028 8522 13030
rect 8214 13008 8522 13028
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5920 11898 5948 12038
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 5630 11792 5686 11801
rect 5356 11756 5408 11762
rect 5630 11727 5686 11736
rect 5356 11698 5408 11704
rect 5172 11620 5224 11626
rect 5172 11562 5224 11568
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4526 10704 4582 10713
rect 4526 10639 4528 10648
rect 4580 10639 4582 10648
rect 4528 10610 4580 10616
rect 4344 10600 4396 10606
rect 4540 10579 4568 10610
rect 4344 10542 4396 10548
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4632 10198 4660 11086
rect 4724 10849 4752 11086
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4710 10840 4766 10849
rect 4710 10775 4766 10784
rect 4908 10674 4936 10950
rect 5000 10810 5028 11494
rect 5276 11218 5304 11494
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3988 9722 4016 9998
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 4080 9382 4108 10134
rect 4908 10130 4936 10610
rect 5184 10470 5212 11018
rect 5276 10674 5304 11154
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5460 10130 5488 11222
rect 5644 11150 5672 11727
rect 5920 11218 5948 11834
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 6012 11082 6040 11698
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 6104 10962 6132 12174
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6932 11354 6960 12106
rect 8036 12102 8064 12718
rect 8588 12442 8616 13262
rect 8760 13252 8812 13258
rect 8760 13194 8812 13200
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8772 12306 8800 13194
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7024 11762 7052 12038
rect 8214 11996 8522 12016
rect 8214 11994 8220 11996
rect 8276 11994 8300 11996
rect 8356 11994 8380 11996
rect 8436 11994 8460 11996
rect 8516 11994 8522 11996
rect 8276 11942 8278 11994
rect 8458 11942 8460 11994
rect 8214 11940 8220 11942
rect 8276 11940 8300 11942
rect 8356 11940 8380 11942
rect 8436 11940 8460 11942
rect 8516 11940 8522 11942
rect 8214 11920 8522 11940
rect 8116 11824 8168 11830
rect 8588 11778 8616 12106
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8116 11766 8168 11772
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7024 11354 7052 11698
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7392 11354 7420 11630
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7852 11286 7880 11494
rect 7944 11354 7972 11562
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 5920 10934 6132 10962
rect 5816 10668 5868 10674
rect 5736 10628 5816 10656
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5184 9674 5212 9998
rect 5552 9722 5580 10406
rect 5736 9994 5764 10628
rect 5816 10610 5868 10616
rect 5920 9994 5948 10934
rect 6564 10674 6592 11086
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6368 10464 6420 10470
rect 6564 10452 6592 10610
rect 6420 10424 6592 10452
rect 6368 10406 6420 10412
rect 6656 10130 6684 10950
rect 6932 10674 6960 11018
rect 7024 11014 7052 11086
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6932 10266 6960 10610
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6644 10124 6696 10130
rect 7024 10112 7052 10406
rect 6644 10066 6696 10072
rect 6932 10084 7052 10112
rect 5724 9988 5776 9994
rect 5724 9930 5776 9936
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5540 9716 5592 9722
rect 4804 9648 4856 9654
rect 5184 9646 5396 9674
rect 5540 9658 5592 9664
rect 4804 9590 4856 9596
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4080 9042 4108 9318
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4816 9178 4844 9590
rect 5368 9518 5396 9646
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 5368 9042 5396 9454
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 5356 9036 5408 9042
rect 5408 8996 5488 9024
rect 5356 8978 5408 8984
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 3804 8838 3832 8910
rect 3792 8832 3844 8838
rect 3712 8780 3792 8786
rect 3712 8774 3844 8780
rect 3712 8758 3832 8774
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 7342 1440 7822
rect 1676 7812 1728 7818
rect 1676 7754 1728 7760
rect 1688 7546 1716 7754
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1412 6254 1440 7278
rect 2056 6798 2084 8434
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2240 7818 2268 8298
rect 2228 7812 2280 7818
rect 2228 7754 2280 7760
rect 2320 7472 2372 7478
rect 2320 7414 2372 7420
rect 2332 7002 2360 7414
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3252 7290 3280 8434
rect 3436 8090 3464 8502
rect 3712 8498 3740 8758
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3436 7410 3464 8026
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3528 7410 3556 7482
rect 3804 7478 3832 8570
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3988 7410 4016 8434
rect 4448 8430 4476 8910
rect 4632 8634 4660 8910
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4632 8498 4660 8570
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4080 7954 4108 8230
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4172 7834 4200 7890
rect 4080 7806 4200 7834
rect 4080 7546 4108 7806
rect 4632 7546 4660 8230
rect 4724 8090 4752 8502
rect 4908 8498 4936 8774
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4908 8378 4936 8434
rect 4804 8356 4856 8362
rect 4908 8350 5120 8378
rect 5276 8362 5304 8842
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 4804 8298 4856 8304
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4816 7818 4844 8298
rect 5092 8022 5120 8350
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 5368 7954 5396 8434
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 4804 7812 4856 7818
rect 4804 7754 4856 7760
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 3528 7290 3556 7346
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2424 6934 2452 7278
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 3160 6798 3188 7278
rect 3252 7262 3556 7290
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1412 5166 1440 6190
rect 2056 5710 2084 6734
rect 2228 6384 2280 6390
rect 2228 6326 2280 6332
rect 2240 5914 2268 6326
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1412 4078 1440 5102
rect 2056 4622 2084 5646
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2228 5296 2280 5302
rect 2228 5238 2280 5244
rect 2240 4826 2268 5238
rect 2884 5216 2912 5510
rect 3160 5370 3188 5646
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 2964 5228 3016 5234
rect 2884 5188 2964 5216
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2424 4826 2452 5102
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2884 4690 2912 5188
rect 2964 5170 3016 5176
rect 3160 4690 3188 5306
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2412 4208 2464 4214
rect 2412 4150 2464 4156
rect 1400 4072 1452 4078
rect 1400 4014 1452 4020
rect 1412 3516 1440 4014
rect 1582 3768 1638 3777
rect 2424 3738 2452 4150
rect 1582 3703 1584 3712
rect 1636 3703 1638 3712
rect 2412 3732 2464 3738
rect 1584 3674 1636 3680
rect 2412 3674 2464 3680
rect 2516 3534 2544 4558
rect 2976 4214 3004 4558
rect 3240 4548 3292 4554
rect 3240 4490 3292 4496
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 2976 3738 3004 4150
rect 3252 4146 3280 4490
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 1584 3528 1636 3534
rect 1412 3488 1584 3516
rect 1584 3470 1636 3476
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 1596 2922 1624 3470
rect 2516 3058 2544 3470
rect 3344 3194 3372 7262
rect 3988 6866 4016 7346
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4528 6928 4580 6934
rect 4528 6870 4580 6876
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3606 6488 3662 6497
rect 3606 6423 3662 6432
rect 3422 6352 3478 6361
rect 3620 6322 3648 6423
rect 3422 6287 3424 6296
rect 3476 6287 3478 6296
rect 3608 6316 3660 6322
rect 3424 6258 3476 6264
rect 3608 6258 3660 6264
rect 3792 6248 3844 6254
rect 3792 6190 3844 6196
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3516 5296 3568 5302
rect 3516 5238 3568 5244
rect 3528 4826 3556 5238
rect 3712 5114 3740 5646
rect 3804 5234 3832 6190
rect 3896 6186 3924 6598
rect 3884 6180 3936 6186
rect 3884 6122 3936 6128
rect 3896 5234 3924 6122
rect 3988 6118 4016 6598
rect 4080 6304 4108 6598
rect 4540 6322 4568 6870
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4160 6316 4212 6322
rect 4080 6276 4160 6304
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5778 4016 6054
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 4080 5234 4108 6276
rect 4160 6258 4212 6264
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4540 6186 4568 6258
rect 4528 6180 4580 6186
rect 4528 6122 4580 6128
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4436 5840 4488 5846
rect 4436 5782 4488 5788
rect 4526 5808 4582 5817
rect 4448 5234 4476 5782
rect 4526 5743 4582 5752
rect 4540 5710 4568 5743
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4632 5642 4660 6802
rect 4724 5914 4752 7278
rect 4908 6866 4936 7278
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4894 6488 4950 6497
rect 4894 6423 4896 6432
rect 4948 6423 4950 6432
rect 4896 6394 4948 6400
rect 4894 6352 4950 6361
rect 4894 6287 4950 6296
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4712 5704 4764 5710
rect 4710 5672 4712 5681
rect 4804 5704 4856 5710
rect 4764 5672 4766 5681
rect 4620 5636 4672 5642
rect 4804 5646 4856 5652
rect 4710 5607 4766 5616
rect 4620 5578 4672 5584
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 3712 5086 3832 5114
rect 3804 5030 3832 5086
rect 4620 5092 4672 5098
rect 4620 5034 4672 5040
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3528 4282 3556 4762
rect 3712 4690 3740 4966
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4632 4826 4660 5034
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 3516 4276 3568 4282
rect 3516 4218 3568 4224
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3436 3738 3464 4014
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3528 3534 3556 4218
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3712 3466 3740 4626
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4080 3942 4108 4558
rect 4448 4554 4476 4626
rect 4436 4548 4488 4554
rect 4436 4490 4488 4496
rect 4448 4146 4476 4490
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4540 4214 4568 4422
rect 4724 4214 4752 5170
rect 4816 4690 4844 5646
rect 4908 5352 4936 6287
rect 5000 5710 5028 7142
rect 5092 6458 5120 7346
rect 5170 6896 5226 6905
rect 5460 6866 5488 8996
rect 5920 8634 5948 9930
rect 6656 9654 6684 10066
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6012 9450 6040 9522
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 6564 9382 6592 9454
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 6012 8634 6040 8842
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5920 8498 5948 8570
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 6472 7886 6500 9318
rect 6656 9178 6684 9454
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6932 9110 6960 10084
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 7024 9586 7052 9930
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6748 8566 6776 8774
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 7116 7886 7144 11154
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7208 10742 7236 11086
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7852 10674 7880 10746
rect 8036 10674 8064 11562
rect 8128 11150 8156 11766
rect 8496 11762 8616 11778
rect 8484 11756 8616 11762
rect 8536 11750 8616 11756
rect 8484 11698 8536 11704
rect 8680 11626 8708 12038
rect 8668 11620 8720 11626
rect 8668 11562 8720 11568
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8220 11218 8248 11494
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8214 10908 8522 10928
rect 8214 10906 8220 10908
rect 8276 10906 8300 10908
rect 8356 10906 8380 10908
rect 8436 10906 8460 10908
rect 8516 10906 8522 10908
rect 8276 10854 8278 10906
rect 8458 10854 8460 10906
rect 8214 10852 8220 10854
rect 8276 10852 8300 10854
rect 8356 10852 8380 10854
rect 8436 10852 8460 10854
rect 8516 10852 8522 10854
rect 8214 10832 8522 10852
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7656 10668 7708 10674
rect 7840 10668 7892 10674
rect 7708 10628 7788 10656
rect 7656 10610 7708 10616
rect 7484 10198 7512 10610
rect 7760 10266 7788 10628
rect 7840 10610 7892 10616
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8404 10470 8432 10610
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7208 9722 7236 9862
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7300 9654 7328 9998
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7208 9178 7236 9522
rect 7392 9450 7420 10066
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 7484 9382 7512 9862
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7484 9178 7512 9318
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7484 8498 7512 8774
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7208 7886 7236 8434
rect 7484 7886 7512 8434
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7668 7834 7696 10202
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7760 8430 7788 9522
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 6472 7478 6500 7822
rect 6644 7812 6696 7818
rect 7668 7806 7788 7834
rect 6644 7754 6696 7760
rect 6460 7472 6512 7478
rect 6460 7414 6512 7420
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5724 7268 5776 7274
rect 5724 7210 5776 7216
rect 5736 7002 5764 7210
rect 5828 7206 5856 7346
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5170 6831 5172 6840
rect 5224 6831 5226 6840
rect 5448 6860 5500 6866
rect 5172 6802 5224 6808
rect 5500 6820 5580 6848
rect 5448 6802 5500 6808
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5092 5914 5120 6394
rect 5184 6322 5212 6666
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5276 5930 5304 6734
rect 5354 6352 5410 6361
rect 5354 6287 5356 6296
rect 5408 6287 5410 6296
rect 5356 6258 5408 6264
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 5184 5902 5304 5930
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4908 5324 5028 5352
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4528 4208 4580 4214
rect 4528 4150 4580 4156
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4448 4026 4476 4082
rect 4448 3998 4660 4026
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4080 3534 4108 3878
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4632 3602 4660 3998
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 4816 3194 4844 4490
rect 4908 4146 4936 5170
rect 5000 4554 5028 5324
rect 5092 4554 5120 5850
rect 5184 5846 5212 5902
rect 5172 5840 5224 5846
rect 5172 5782 5224 5788
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 5276 5234 5304 5782
rect 5460 5710 5488 6054
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5368 4690 5396 5578
rect 5552 5556 5580 6820
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5644 6322 5672 6666
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5736 6390 5764 6598
rect 6012 6458 6040 7346
rect 6656 7342 6684 7754
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5724 6384 5776 6390
rect 5724 6326 5776 6332
rect 6380 6322 6408 7142
rect 6656 6322 6684 7278
rect 6748 6934 6776 7346
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6748 6322 6776 6870
rect 7024 6730 7052 7686
rect 7576 7478 7604 7686
rect 7564 7472 7616 7478
rect 7564 7414 7616 7420
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7286 6896 7342 6905
rect 7286 6831 7342 6840
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 5644 6186 5672 6258
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 6104 5914 6132 6258
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 6288 5914 6316 6190
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6104 5778 6132 5850
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6460 5704 6512 5710
rect 6656 5692 6684 6258
rect 7116 6186 7144 6326
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 7104 6180 7156 6186
rect 7104 6122 7156 6128
rect 6512 5664 6684 5692
rect 6460 5646 6512 5652
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 5460 5528 5580 5556
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 5080 4548 5132 4554
rect 5080 4490 5132 4496
rect 5000 4282 5028 4490
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 5092 3534 5120 4490
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 1584 2916 1636 2922
rect 1584 2858 1636 2864
rect 1596 2514 1624 2858
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 1596 2038 1624 2450
rect 1584 2032 1636 2038
rect 1584 1974 1636 1980
rect 2228 2032 2280 2038
rect 2228 1974 2280 1980
rect 940 1760 992 1766
rect 940 1702 992 1708
rect 952 800 980 1702
rect 2240 1562 2268 1974
rect 2228 1556 2280 1562
rect 2228 1498 2280 1504
rect 2516 1358 2544 2994
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2608 2378 2636 2790
rect 2884 2514 2912 2994
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3436 2650 3464 2926
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4632 2650 4660 3062
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 5000 2774 5028 2858
rect 4908 2746 5028 2774
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 2884 1834 2912 2450
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 3424 2032 3476 2038
rect 3424 1974 3476 1980
rect 3056 1896 3108 1902
rect 3056 1838 3108 1844
rect 2872 1828 2924 1834
rect 2872 1770 2924 1776
rect 2504 1352 2556 1358
rect 2504 1294 2556 1300
rect 3068 1290 3096 1838
rect 3436 1562 3464 1974
rect 4214 1660 4522 1680
rect 4214 1658 4220 1660
rect 4276 1658 4300 1660
rect 4356 1658 4380 1660
rect 4436 1658 4460 1660
rect 4516 1658 4522 1660
rect 4276 1606 4278 1658
rect 4458 1606 4460 1658
rect 4214 1604 4220 1606
rect 4276 1604 4300 1606
rect 4356 1604 4380 1606
rect 4436 1604 4460 1606
rect 4516 1604 4522 1606
rect 4214 1584 4522 1604
rect 3424 1556 3476 1562
rect 3424 1498 3476 1504
rect 4632 1290 4660 2246
rect 2780 1284 2832 1290
rect 2780 1226 2832 1232
rect 3056 1284 3108 1290
rect 3056 1226 3108 1232
rect 4620 1284 4672 1290
rect 4620 1226 4672 1232
rect 2792 800 2820 1226
rect 4632 870 4752 898
rect 4632 800 4660 870
rect 938 0 994 800
rect 2778 0 2834 800
rect 4618 0 4674 800
rect 4724 762 4752 870
rect 4908 762 4936 2746
rect 5184 2514 5212 3606
rect 5368 3194 5396 4626
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5264 2984 5316 2990
rect 5460 2972 5488 5528
rect 6196 5302 6224 5578
rect 6564 5302 6592 5664
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 6184 5296 6236 5302
rect 6184 5238 6236 5244
rect 6552 5296 6604 5302
rect 6552 5238 6604 5244
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5552 4690 5580 5102
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5644 4622 5672 5238
rect 6748 5234 6776 6122
rect 7116 5817 7144 6122
rect 7102 5808 7158 5817
rect 7102 5743 7158 5752
rect 7208 5574 7236 6258
rect 7300 6186 7328 6831
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7288 6180 7340 6186
rect 7288 6122 7340 6128
rect 7300 5846 7328 6122
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6184 5092 6236 5098
rect 6184 5034 6236 5040
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5552 3942 5580 4490
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5316 2944 5488 2972
rect 5264 2926 5316 2932
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 5276 2378 5304 2926
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 5276 1970 5304 2314
rect 5736 2106 5764 4966
rect 6196 4826 6224 5034
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6472 4282 6500 4966
rect 6840 4622 6868 5238
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5828 3534 5856 3878
rect 5920 3738 5948 4082
rect 6380 3738 6408 4082
rect 6840 4010 6868 4558
rect 6932 4282 6960 5102
rect 7300 4826 7328 5238
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7196 4616 7248 4622
rect 7194 4584 7196 4593
rect 7248 4584 7250 4593
rect 7194 4519 7250 4528
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 7392 4146 7420 6598
rect 7484 6458 7512 7346
rect 7668 7342 7696 7686
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7760 6866 7788 7806
rect 7944 7546 7972 10406
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8220 10062 8248 10202
rect 8404 10062 8432 10406
rect 8588 10198 8616 10950
rect 8772 10810 8800 11086
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8576 10192 8628 10198
rect 8576 10134 8628 10140
rect 8772 10130 8800 10746
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8214 9820 8522 9840
rect 8214 9818 8220 9820
rect 8276 9818 8300 9820
rect 8356 9818 8380 9820
rect 8436 9818 8460 9820
rect 8516 9818 8522 9820
rect 8276 9766 8278 9818
rect 8458 9766 8460 9818
rect 8214 9764 8220 9766
rect 8276 9764 8300 9766
rect 8356 9764 8380 9766
rect 8436 9764 8460 9766
rect 8516 9764 8522 9766
rect 8214 9744 8522 9764
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8036 8906 8064 9522
rect 8404 9178 8432 9590
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8496 9178 8524 9454
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 8214 8732 8522 8752
rect 8214 8730 8220 8732
rect 8276 8730 8300 8732
rect 8356 8730 8380 8732
rect 8436 8730 8460 8732
rect 8516 8730 8522 8732
rect 8276 8678 8278 8730
rect 8458 8678 8460 8730
rect 8214 8676 8220 8678
rect 8276 8676 8300 8678
rect 8356 8676 8380 8678
rect 8436 8676 8460 8678
rect 8516 8676 8522 8678
rect 8214 8656 8522 8676
rect 8214 7644 8522 7664
rect 8214 7642 8220 7644
rect 8276 7642 8300 7644
rect 8356 7642 8380 7644
rect 8436 7642 8460 7644
rect 8516 7642 8522 7644
rect 8276 7590 8278 7642
rect 8458 7590 8460 7642
rect 8214 7588 8220 7590
rect 8276 7588 8300 7590
rect 8356 7588 8380 7590
rect 8436 7588 8460 7590
rect 8516 7588 8522 7590
rect 8214 7568 8522 7588
rect 8588 7546 8616 8910
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8680 7886 8708 8434
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8772 8022 8800 8298
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8680 7410 8708 7822
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8404 6934 8432 7346
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 7760 6746 7788 6802
rect 7668 6718 7788 6746
rect 7932 6724 7984 6730
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7484 6225 7512 6258
rect 7470 6216 7526 6225
rect 7668 6186 7696 6718
rect 7932 6666 7984 6672
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7760 6390 7788 6598
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7470 6151 7526 6160
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 7944 5914 7972 6666
rect 8036 6662 8064 6802
rect 8680 6730 8708 7210
rect 8772 6798 8800 7686
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8214 6556 8522 6576
rect 8214 6554 8220 6556
rect 8276 6554 8300 6556
rect 8356 6554 8380 6556
rect 8436 6554 8460 6556
rect 8516 6554 8522 6556
rect 8276 6502 8278 6554
rect 8458 6502 8460 6554
rect 8214 6500 8220 6502
rect 8276 6500 8300 6502
rect 8356 6500 8380 6502
rect 8436 6500 8460 6502
rect 8516 6500 8522 6502
rect 8214 6480 8522 6500
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 8036 5914 8064 6122
rect 8220 5930 8248 6258
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8312 6118 8340 6190
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8220 5914 8340 5930
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 8024 5908 8076 5914
rect 8220 5908 8352 5914
rect 8220 5902 8300 5908
rect 8024 5850 8076 5856
rect 8300 5850 8352 5856
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7562 5672 7618 5681
rect 7562 5607 7618 5616
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7484 4622 7512 5510
rect 7576 5098 7604 5607
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5828 2310 5856 2994
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 5920 2378 5948 2790
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5724 2100 5776 2106
rect 5724 2042 5776 2048
rect 5264 1964 5316 1970
rect 5264 1906 5316 1912
rect 5448 1964 5500 1970
rect 5448 1906 5500 1912
rect 5276 1290 5304 1906
rect 5356 1760 5408 1766
rect 5356 1702 5408 1708
rect 5368 1426 5396 1702
rect 5356 1420 5408 1426
rect 5356 1362 5408 1368
rect 5264 1284 5316 1290
rect 5264 1226 5316 1232
rect 5460 1222 5488 1906
rect 5736 1834 5764 2042
rect 5724 1828 5776 1834
rect 5724 1770 5776 1776
rect 5828 1562 5856 2246
rect 6012 1970 6040 3606
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 6000 1964 6052 1970
rect 6000 1906 6052 1912
rect 5816 1556 5868 1562
rect 5816 1498 5868 1504
rect 5828 1426 5856 1498
rect 5816 1420 5868 1426
rect 5816 1362 5868 1368
rect 6196 1358 6224 2790
rect 6656 2650 6684 3470
rect 6840 3466 6868 3946
rect 7024 3602 7052 4082
rect 7484 3942 7512 4558
rect 7576 4486 7604 5034
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 7484 3534 7512 3878
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 7472 3392 7524 3398
rect 7576 3380 7604 4422
rect 7668 3738 7696 5714
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7852 5302 7880 5646
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 8036 4690 8064 5850
rect 8404 5642 8432 6258
rect 8588 6254 8616 6598
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8680 5710 8708 6666
rect 8772 5896 8800 6734
rect 8864 6458 8892 12786
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 9048 11830 9076 12242
rect 9036 11824 9088 11830
rect 9036 11766 9088 11772
rect 9128 10804 9180 10810
rect 8956 10764 9128 10792
rect 8956 10266 8984 10764
rect 9128 10746 9180 10752
rect 9140 10674 9168 10746
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9048 10266 9076 10610
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9232 10198 9260 10542
rect 9220 10192 9272 10198
rect 9220 10134 9272 10140
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8956 7886 8984 9522
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9048 9042 9076 9318
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9324 8090 9352 13126
rect 9416 12986 9444 13330
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9600 12850 9628 13398
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9692 12442 9720 14200
rect 10888 13530 10916 14447
rect 11242 14200 11298 15000
rect 12714 14200 12770 15000
rect 14186 14200 14242 15000
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 9784 12918 9812 13466
rect 10046 13424 10102 13433
rect 10046 13359 10102 13368
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9600 11762 9628 12174
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9692 11830 9720 12106
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9784 11762 9812 12854
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9784 11234 9812 11698
rect 9876 11694 9904 12378
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9876 11354 9904 11630
rect 9968 11558 9996 12174
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9692 11218 9812 11234
rect 9680 11212 9812 11218
rect 9732 11206 9812 11212
rect 9680 11154 9732 11160
rect 9692 11082 9720 11154
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9692 9926 9720 11018
rect 9784 10674 9812 11086
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9692 9178 9720 9862
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9600 8566 9628 8774
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9140 7342 9168 7754
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 9048 6934 9076 7210
rect 9036 6928 9088 6934
rect 9036 6870 9088 6876
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8956 6458 8984 6598
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 9048 6322 9076 6870
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8772 5868 8892 5896
rect 8760 5772 8812 5778
rect 8760 5714 8812 5720
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8128 5098 8156 5578
rect 8666 5536 8722 5545
rect 8214 5468 8522 5488
rect 8666 5471 8722 5480
rect 8214 5466 8220 5468
rect 8276 5466 8300 5468
rect 8356 5466 8380 5468
rect 8436 5466 8460 5468
rect 8516 5466 8522 5468
rect 8276 5414 8278 5466
rect 8458 5414 8460 5466
rect 8214 5412 8220 5414
rect 8276 5412 8300 5414
rect 8356 5412 8380 5414
rect 8436 5412 8460 5414
rect 8516 5412 8522 5414
rect 8214 5392 8522 5412
rect 8680 5370 8708 5471
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8576 5296 8628 5302
rect 8576 5238 8628 5244
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 7838 4584 7894 4593
rect 7838 4519 7840 4528
rect 7892 4519 7894 4528
rect 7840 4490 7892 4496
rect 8036 4214 8064 4626
rect 8404 4622 8432 4966
rect 8588 4622 8616 5238
rect 8772 4758 8800 5714
rect 8760 4752 8812 4758
rect 8760 4694 8812 4700
rect 8392 4616 8444 4622
rect 8576 4616 8628 4622
rect 8392 4558 8444 4564
rect 8574 4584 8576 4593
rect 8628 4584 8630 4593
rect 8574 4519 8630 4528
rect 8214 4380 8522 4400
rect 8214 4378 8220 4380
rect 8276 4378 8300 4380
rect 8356 4378 8380 4380
rect 8436 4378 8460 4380
rect 8516 4378 8522 4380
rect 8276 4326 8278 4378
rect 8458 4326 8460 4378
rect 8214 4324 8220 4326
rect 8276 4324 8300 4326
rect 8356 4324 8380 4326
rect 8436 4324 8460 4326
rect 8516 4324 8522 4326
rect 8214 4304 8522 4324
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7852 3534 7880 4082
rect 8300 4072 8352 4078
rect 8588 4026 8616 4519
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8300 4014 8352 4020
rect 8312 3670 8340 4014
rect 8496 3998 8616 4026
rect 8300 3664 8352 3670
rect 8300 3606 8352 3612
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 8392 3528 8444 3534
rect 8496 3516 8524 3998
rect 8680 3942 8708 4422
rect 8864 4010 8892 5868
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8956 5234 8984 5646
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8956 5137 8984 5170
rect 8942 5128 8998 5137
rect 8942 5063 8998 5072
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8852 4004 8904 4010
rect 8852 3946 8904 3952
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8588 3534 8616 3878
rect 8444 3488 8524 3516
rect 8576 3528 8628 3534
rect 8392 3470 8444 3476
rect 8576 3470 8628 3476
rect 7524 3352 7604 3380
rect 7656 3392 7708 3398
rect 7472 3334 7524 3340
rect 7656 3334 7708 3340
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 7024 2514 7052 3130
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7484 2582 7512 3062
rect 7668 2582 7696 3334
rect 7852 3058 7880 3470
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 7944 3126 7972 3334
rect 8128 3194 8156 3334
rect 8214 3292 8522 3312
rect 8214 3290 8220 3292
rect 8276 3290 8300 3292
rect 8356 3290 8380 3292
rect 8436 3290 8460 3292
rect 8516 3290 8522 3292
rect 8276 3238 8278 3290
rect 8458 3238 8460 3290
rect 8214 3236 8220 3238
rect 8276 3236 8300 3238
rect 8356 3236 8380 3238
rect 8436 3236 8460 3238
rect 8516 3236 8522 3238
rect 8214 3216 8522 3236
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 8128 2582 8156 2994
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6472 1970 6500 2246
rect 7760 2106 7788 2382
rect 8576 2372 8628 2378
rect 8576 2314 8628 2320
rect 8214 2204 8522 2224
rect 8214 2202 8220 2204
rect 8276 2202 8300 2204
rect 8356 2202 8380 2204
rect 8436 2202 8460 2204
rect 8516 2202 8522 2204
rect 8276 2150 8278 2202
rect 8458 2150 8460 2202
rect 8214 2148 8220 2150
rect 8276 2148 8300 2150
rect 8356 2148 8380 2150
rect 8436 2148 8460 2150
rect 8516 2148 8522 2150
rect 8214 2128 8522 2148
rect 7748 2100 7800 2106
rect 7748 2042 7800 2048
rect 6460 1964 6512 1970
rect 6460 1906 6512 1912
rect 7564 1964 7616 1970
rect 7564 1906 7616 1912
rect 7012 1760 7064 1766
rect 7012 1702 7064 1708
rect 6552 1556 6604 1562
rect 6552 1498 6604 1504
rect 6184 1352 6236 1358
rect 6184 1294 6236 1300
rect 5448 1216 5500 1222
rect 5448 1158 5500 1164
rect 6564 800 6592 1498
rect 7024 1358 7052 1702
rect 7576 1494 7604 1906
rect 7564 1488 7616 1494
rect 7564 1430 7616 1436
rect 7760 1358 7788 2042
rect 8588 1834 8616 2314
rect 8576 1828 8628 1834
rect 8576 1770 8628 1776
rect 8588 1494 8616 1770
rect 8576 1488 8628 1494
rect 8576 1430 8628 1436
rect 7012 1352 7064 1358
rect 7012 1294 7064 1300
rect 7748 1352 7800 1358
rect 7748 1294 7800 1300
rect 8214 1116 8522 1136
rect 8214 1114 8220 1116
rect 8276 1114 8300 1116
rect 8356 1114 8380 1116
rect 8436 1114 8460 1116
rect 8516 1114 8522 1116
rect 8276 1062 8278 1114
rect 8458 1062 8460 1114
rect 8214 1060 8220 1062
rect 8276 1060 8300 1062
rect 8356 1060 8380 1062
rect 8436 1060 8460 1062
rect 8516 1060 8522 1062
rect 8214 1040 8522 1060
rect 8404 870 8524 898
rect 8404 800 8432 870
rect 4724 734 4936 762
rect 6550 0 6606 800
rect 8390 0 8446 800
rect 8496 762 8524 870
rect 8680 762 8708 3878
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8772 3369 8800 3470
rect 8864 3398 8892 3946
rect 8956 3942 8984 4626
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8956 3398 8984 3878
rect 9048 3534 9076 5578
rect 9140 4078 9168 6666
rect 9232 5284 9260 7958
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9416 7546 9444 7822
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9312 7472 9364 7478
rect 9364 7420 9444 7426
rect 9312 7414 9444 7420
rect 9324 7398 9444 7414
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9324 6322 9352 7278
rect 9416 7154 9444 7398
rect 9508 7154 9536 7890
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9416 7126 9536 7154
rect 9416 6866 9444 7126
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9324 5953 9352 6258
rect 9310 5944 9366 5953
rect 9310 5879 9366 5888
rect 9312 5704 9364 5710
rect 9310 5672 9312 5681
rect 9364 5672 9366 5681
rect 9310 5607 9366 5616
rect 9312 5296 9364 5302
rect 9232 5256 9312 5284
rect 9312 5238 9364 5244
rect 9310 5128 9366 5137
rect 9310 5063 9366 5072
rect 9324 4622 9352 5063
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9416 4468 9444 6802
rect 9508 6730 9536 6938
rect 9600 6914 9628 7414
rect 9784 7410 9812 10610
rect 9968 8090 9996 10610
rect 10060 10198 10088 13359
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10520 12170 10548 12786
rect 10704 12238 10732 13126
rect 11164 12918 11192 13262
rect 11152 12912 11204 12918
rect 11152 12854 11204 12860
rect 10782 12744 10838 12753
rect 10782 12679 10838 12688
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10520 11762 10548 12106
rect 10796 11914 10824 12679
rect 10876 12164 10928 12170
rect 10876 12106 10928 12112
rect 10704 11898 10824 11914
rect 10692 11892 10824 11898
rect 10744 11886 10824 11892
rect 10692 11834 10744 11840
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10152 10742 10180 11698
rect 10796 11626 10824 11886
rect 10888 11762 10916 12106
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10980 11898 11008 12038
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 10784 11620 10836 11626
rect 10784 11562 10836 11568
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10600 11008 10652 11014
rect 10322 10976 10378 10985
rect 10600 10950 10652 10956
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10322 10911 10378 10920
rect 10336 10810 10364 10911
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 10612 10674 10640 10950
rect 10704 10674 10732 10950
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10520 10266 10548 10406
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10048 10192 10100 10198
rect 10520 10169 10548 10202
rect 10048 10134 10100 10140
rect 10506 10160 10562 10169
rect 10506 10095 10562 10104
rect 10704 9994 10732 10610
rect 10692 9988 10744 9994
rect 10692 9930 10744 9936
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10060 8634 10088 9522
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10508 9444 10560 9450
rect 10508 9386 10560 9392
rect 10414 9072 10470 9081
rect 10414 9007 10470 9016
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10060 7818 10088 7958
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 10324 7812 10376 7818
rect 10324 7754 10376 7760
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9600 6886 9720 6914
rect 9692 6780 9720 6886
rect 9772 6792 9824 6798
rect 9692 6752 9772 6780
rect 9772 6734 9824 6740
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9496 6248 9548 6254
rect 9494 6216 9496 6225
rect 9548 6216 9550 6225
rect 9692 6186 9720 6598
rect 9494 6151 9550 6160
rect 9680 6180 9732 6186
rect 9680 6122 9732 6128
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9232 4440 9444 4468
rect 9232 4146 9260 4440
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9324 3652 9352 4150
rect 9416 3738 9444 4440
rect 9508 4049 9536 6054
rect 9692 5846 9720 6122
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9600 5273 9628 5714
rect 9784 5352 9812 6734
rect 9876 6730 9904 7210
rect 9968 6866 9996 7414
rect 10060 7410 10088 7754
rect 10336 7478 10364 7754
rect 10324 7472 10376 7478
rect 10324 7414 10376 7420
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10244 6934 10272 7210
rect 10232 6928 10284 6934
rect 10232 6870 10284 6876
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9864 6724 9916 6730
rect 9864 6666 9916 6672
rect 9784 5324 9904 5352
rect 9586 5264 9642 5273
rect 9876 5250 9904 5324
rect 9586 5199 9642 5208
rect 9784 5222 9904 5250
rect 9600 5166 9628 5199
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9494 4040 9550 4049
rect 9494 3975 9550 3984
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9232 3624 9352 3652
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8852 3392 8904 3398
rect 8758 3360 8814 3369
rect 8852 3334 8904 3340
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8758 3295 8814 3304
rect 8956 2990 8984 3334
rect 9232 3058 9260 3624
rect 9416 3398 9444 3674
rect 9784 3528 9812 5222
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9876 4826 9904 4966
rect 9968 4865 9996 6802
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10060 5574 10088 6054
rect 10152 5681 10180 6598
rect 10244 6186 10272 6870
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10336 6458 10364 6802
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 10138 5672 10194 5681
rect 10138 5607 10194 5616
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10060 5137 10088 5510
rect 10152 5370 10180 5510
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10046 5128 10102 5137
rect 10244 5098 10272 5782
rect 10428 5386 10456 9007
rect 10520 8974 10548 9386
rect 10612 8974 10640 9454
rect 10704 9110 10732 9930
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10520 5914 10548 8366
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10336 5358 10456 5386
rect 10046 5063 10102 5072
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 9954 4856 10010 4865
rect 9864 4820 9916 4826
rect 9954 4791 10010 4800
rect 9864 4762 9916 4768
rect 9968 4622 9996 4791
rect 10152 4622 10180 4966
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 10060 4146 10088 4422
rect 10152 4214 10180 4558
rect 10140 4208 10192 4214
rect 10140 4150 10192 4156
rect 10244 4146 10272 4558
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9772 3522 9824 3528
rect 9772 3464 9824 3470
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9402 3224 9458 3233
rect 9402 3159 9458 3168
rect 9588 3188 9640 3194
rect 9416 3058 9444 3159
rect 9588 3130 9640 3136
rect 9600 3097 9628 3130
rect 9586 3088 9642 3097
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9404 3052 9456 3058
rect 9586 3023 9642 3032
rect 9404 2994 9456 3000
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 9600 2650 9628 3023
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 8956 2106 8984 2382
rect 9312 2372 9364 2378
rect 9312 2314 9364 2320
rect 8944 2100 8996 2106
rect 8944 2042 8996 2048
rect 9324 1426 9352 2314
rect 9508 1562 9536 2518
rect 9692 2514 9720 2926
rect 9680 2508 9732 2514
rect 9876 2496 9904 3878
rect 9968 3670 9996 4082
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 9680 2450 9732 2456
rect 9784 2468 9904 2496
rect 9784 2310 9812 2468
rect 9864 2372 9916 2378
rect 9864 2314 9916 2320
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9600 1970 9628 2246
rect 9876 2038 9904 2314
rect 9864 2032 9916 2038
rect 9864 1974 9916 1980
rect 9588 1964 9640 1970
rect 9588 1906 9640 1912
rect 9496 1556 9548 1562
rect 9496 1498 9548 1504
rect 9312 1420 9364 1426
rect 9312 1362 9364 1368
rect 9600 1358 9628 1906
rect 9876 1494 9904 1974
rect 9864 1488 9916 1494
rect 9864 1430 9916 1436
rect 9588 1352 9640 1358
rect 9588 1294 9640 1300
rect 9968 1290 9996 2858
rect 10060 2106 10088 3334
rect 10244 3194 10272 3334
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10048 2100 10100 2106
rect 10048 2042 10100 2048
rect 10336 2038 10364 5358
rect 10506 5264 10562 5273
rect 10506 5199 10508 5208
rect 10560 5199 10562 5208
rect 10508 5170 10560 5176
rect 10416 5092 10468 5098
rect 10416 5034 10468 5040
rect 10428 4690 10456 5034
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10520 4622 10548 4762
rect 10508 4616 10560 4622
rect 10414 4584 10470 4593
rect 10508 4558 10560 4564
rect 10414 4519 10416 4528
rect 10468 4519 10470 4528
rect 10416 4490 10468 4496
rect 10428 4128 10456 4490
rect 10428 4100 10548 4128
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 10428 3369 10456 3946
rect 10520 3670 10548 4100
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10414 3360 10470 3369
rect 10414 3295 10470 3304
rect 10428 3058 10456 3295
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10508 2916 10560 2922
rect 10508 2858 10560 2864
rect 10520 2650 10548 2858
rect 10612 2854 10640 8910
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10704 6798 10732 7822
rect 10888 7546 10916 8978
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10888 6934 10916 7482
rect 10980 7002 11008 11494
rect 11072 11286 11100 11698
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 11072 10742 11100 11222
rect 11060 10736 11112 10742
rect 11060 10678 11112 10684
rect 11256 9042 11284 14200
rect 12214 13628 12522 13648
rect 12214 13626 12220 13628
rect 12276 13626 12300 13628
rect 12356 13626 12380 13628
rect 12436 13626 12460 13628
rect 12516 13626 12522 13628
rect 12276 13574 12278 13626
rect 12458 13574 12460 13626
rect 12214 13572 12220 13574
rect 12276 13572 12300 13574
rect 12356 13572 12380 13574
rect 12436 13572 12460 13574
rect 12516 13572 12522 13574
rect 12214 13552 12522 13572
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11716 12850 11744 13126
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11704 12708 11756 12714
rect 11704 12650 11756 12656
rect 11716 12306 11744 12650
rect 11992 12374 12020 13126
rect 12084 12374 12112 13262
rect 12214 12540 12522 12560
rect 12214 12538 12220 12540
rect 12276 12538 12300 12540
rect 12356 12538 12380 12540
rect 12436 12538 12460 12540
rect 12516 12538 12522 12540
rect 12276 12486 12278 12538
rect 12458 12486 12460 12538
rect 12214 12484 12220 12486
rect 12276 12484 12300 12486
rect 12356 12484 12380 12486
rect 12436 12484 12460 12486
rect 12516 12484 12522 12486
rect 12214 12464 12522 12484
rect 11980 12368 12032 12374
rect 11980 12310 12032 12316
rect 12072 12368 12124 12374
rect 12072 12310 12124 12316
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 12636 12238 12664 13262
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 11440 11558 11468 12174
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11624 11937 11652 12038
rect 11610 11928 11666 11937
rect 11610 11863 11666 11872
rect 12728 11778 12756 14200
rect 13176 13252 13228 13258
rect 13176 13194 13228 13200
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13188 12238 13216 13194
rect 13280 12986 13308 13194
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 13280 12374 13308 12650
rect 13268 12368 13320 12374
rect 13268 12310 13320 12316
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13280 11830 13308 12310
rect 13372 12170 13400 12786
rect 13464 12306 13492 13126
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13360 12164 13412 12170
rect 13360 12106 13412 12112
rect 13268 11824 13320 11830
rect 12728 11750 12940 11778
rect 13268 11766 13320 11772
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11900 11218 11928 11630
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 12214 11452 12522 11472
rect 12214 11450 12220 11452
rect 12276 11450 12300 11452
rect 12356 11450 12380 11452
rect 12436 11450 12460 11452
rect 12516 11450 12522 11452
rect 12276 11398 12278 11450
rect 12458 11398 12460 11450
rect 12214 11396 12220 11398
rect 12276 11396 12300 11398
rect 12356 11396 12380 11398
rect 12436 11396 12460 11398
rect 12516 11396 12522 11398
rect 12214 11376 12522 11396
rect 12820 11286 12848 11562
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 12452 10742 12480 11222
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11624 9994 11652 10610
rect 12728 10606 12756 11086
rect 12808 11076 12860 11082
rect 12808 11018 12860 11024
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11808 10130 11836 10406
rect 12214 10364 12522 10384
rect 12214 10362 12220 10364
rect 12276 10362 12300 10364
rect 12356 10362 12380 10364
rect 12436 10362 12460 10364
rect 12516 10362 12522 10364
rect 12276 10310 12278 10362
rect 12458 10310 12460 10362
rect 12214 10308 12220 10310
rect 12276 10308 12300 10310
rect 12356 10308 12380 10310
rect 12436 10308 12460 10310
rect 12516 10308 12522 10310
rect 12214 10288 12522 10308
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11532 9178 11560 9522
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11164 8022 11192 8774
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 11532 7886 11560 8434
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 10876 6928 10928 6934
rect 10796 6888 10876 6916
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10704 5914 10732 6734
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10796 5778 10824 6888
rect 10876 6870 10928 6876
rect 11348 6866 11376 7142
rect 11532 6934 11560 7822
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11520 6928 11572 6934
rect 11520 6870 11572 6876
rect 11624 6866 11652 7142
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11152 6792 11204 6798
rect 11072 6752 11152 6780
rect 11072 6390 11100 6752
rect 11152 6734 11204 6740
rect 11348 6633 11376 6802
rect 11334 6624 11390 6633
rect 11334 6559 11390 6568
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 10876 6248 10928 6254
rect 10874 6216 10876 6225
rect 10928 6216 10930 6225
rect 10874 6151 10930 6160
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10888 5642 10916 6054
rect 11072 5710 11100 6326
rect 11716 5914 11744 9998
rect 12452 9586 12480 9998
rect 12636 9586 12664 10474
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12214 9276 12522 9296
rect 12214 9274 12220 9276
rect 12276 9274 12300 9276
rect 12356 9274 12380 9276
rect 12436 9274 12460 9276
rect 12516 9274 12522 9276
rect 12276 9222 12278 9274
rect 12458 9222 12460 9274
rect 12214 9220 12220 9222
rect 12276 9220 12300 9222
rect 12356 9220 12380 9222
rect 12436 9220 12460 9222
rect 12516 9220 12522 9222
rect 12214 9200 12522 9220
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12636 8634 12664 9046
rect 12728 8634 12756 10542
rect 12820 10266 12848 11018
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12912 10112 12940 11750
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13464 11150 13492 11698
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 13188 10742 13216 11018
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 12820 10084 12940 10112
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 11808 7886 11836 8366
rect 12214 8188 12522 8208
rect 12214 8186 12220 8188
rect 12276 8186 12300 8188
rect 12356 8186 12380 8188
rect 12436 8186 12460 8188
rect 12516 8186 12522 8188
rect 12276 8134 12278 8186
rect 12458 8134 12460 8186
rect 12214 8132 12220 8134
rect 12276 8132 12300 8134
rect 12356 8132 12380 8134
rect 12436 8132 12460 8134
rect 12516 8132 12522 8134
rect 12214 8112 12522 8132
rect 12636 8022 12664 8366
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 11796 7880 11848 7886
rect 11848 7828 11928 7834
rect 11796 7822 11928 7828
rect 11808 7806 11928 7822
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11808 7410 11836 7686
rect 11900 7546 11928 7806
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 12214 7100 12522 7120
rect 12214 7098 12220 7100
rect 12276 7098 12300 7100
rect 12356 7098 12380 7100
rect 12436 7098 12460 7100
rect 12516 7098 12522 7100
rect 12276 7046 12278 7098
rect 12458 7046 12460 7098
rect 12214 7044 12220 7046
rect 12276 7044 12300 7046
rect 12356 7044 12380 7046
rect 12436 7044 12460 7046
rect 12516 7044 12522 7046
rect 12214 7024 12522 7044
rect 12636 6914 12664 7958
rect 12820 7546 12848 10084
rect 13188 10062 13216 10678
rect 13464 10674 13492 11086
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 12900 9988 12952 9994
rect 12900 9930 12952 9936
rect 12912 9450 12940 9930
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13372 9654 13400 9862
rect 14200 9722 14228 14200
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 12912 8974 12940 9386
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 13096 8906 13124 9522
rect 13372 9110 13400 9590
rect 13360 9104 13412 9110
rect 13360 9046 13412 9052
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12912 7478 12940 8502
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12912 7002 12940 7414
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12544 6886 12664 6914
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10690 5264 10746 5273
rect 10690 5199 10692 5208
rect 10744 5199 10746 5208
rect 10692 5170 10744 5176
rect 10796 5098 10824 5510
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10784 5092 10836 5098
rect 10784 5034 10836 5040
rect 10704 4554 10732 5034
rect 10796 4826 10824 5034
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10704 3058 10732 4150
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 10324 2032 10376 2038
rect 10324 1974 10376 1980
rect 10612 1902 10640 2450
rect 10796 2378 10824 3946
rect 10888 2582 10916 5578
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 10980 5273 11008 5306
rect 10966 5264 11022 5273
rect 11072 5234 11100 5646
rect 10966 5199 11022 5208
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11164 5114 11192 5782
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 11072 5086 11192 5114
rect 11072 5030 11100 5086
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 11072 4214 11100 4966
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10968 3664 11020 3670
rect 10968 3606 11020 3612
rect 10980 2922 11008 3606
rect 11072 3466 11100 3878
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 11058 3360 11114 3369
rect 11058 3295 11114 3304
rect 11072 3058 11100 3295
rect 11060 3052 11112 3058
rect 11112 3012 11192 3040
rect 11060 2994 11112 3000
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 10876 2576 10928 2582
rect 11072 2530 11100 2858
rect 10876 2518 10928 2524
rect 10980 2502 11100 2530
rect 10784 2372 10836 2378
rect 10784 2314 10836 2320
rect 10690 2136 10746 2145
rect 10690 2071 10746 2080
rect 10600 1896 10652 1902
rect 10600 1838 10652 1844
rect 10324 1760 10376 1766
rect 10324 1702 10376 1708
rect 10336 1426 10364 1702
rect 10612 1562 10640 1838
rect 10600 1556 10652 1562
rect 10600 1498 10652 1504
rect 10324 1420 10376 1426
rect 10324 1362 10376 1368
rect 10704 1358 10732 2071
rect 10876 1896 10928 1902
rect 10876 1838 10928 1844
rect 10888 1358 10916 1838
rect 10692 1352 10744 1358
rect 10692 1294 10744 1300
rect 10876 1352 10928 1358
rect 10876 1294 10928 1300
rect 9956 1284 10008 1290
rect 9956 1226 10008 1232
rect 10244 870 10364 898
rect 10244 800 10272 870
rect 8496 734 8708 762
rect 10230 0 10286 800
rect 10336 762 10364 870
rect 10980 762 11008 2502
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11072 1426 11100 2382
rect 11164 2310 11192 3012
rect 11256 2650 11284 5714
rect 11520 5296 11572 5302
rect 11520 5238 11572 5244
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 11440 4865 11468 5102
rect 11426 4856 11482 4865
rect 11426 4791 11482 4800
rect 11532 4622 11560 5238
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11532 4214 11560 4558
rect 11808 4282 11836 6734
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11992 6458 12020 6598
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11980 6248 12032 6254
rect 11978 6216 11980 6225
rect 12032 6216 12034 6225
rect 11978 6151 12034 6160
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11900 5710 11928 6054
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 11992 5370 12020 6151
rect 12084 5778 12112 6734
rect 12544 6390 12572 6886
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12532 6384 12584 6390
rect 12532 6326 12584 6332
rect 12214 6012 12522 6032
rect 12214 6010 12220 6012
rect 12276 6010 12300 6012
rect 12356 6010 12380 6012
rect 12436 6010 12460 6012
rect 12516 6010 12522 6012
rect 12276 5958 12278 6010
rect 12458 5958 12460 6010
rect 12214 5956 12220 5958
rect 12276 5956 12300 5958
rect 12356 5956 12380 5958
rect 12436 5956 12460 5958
rect 12516 5956 12522 5958
rect 12214 5936 12522 5956
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 12084 5681 12112 5714
rect 12532 5704 12584 5710
rect 12070 5672 12126 5681
rect 12636 5692 12664 6598
rect 13096 6322 13124 8434
rect 13188 7886 13216 8842
rect 13268 8424 13320 8430
rect 13266 8392 13268 8401
rect 13320 8392 13322 8401
rect 13266 8327 13322 8336
rect 13280 8090 13308 8327
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13266 7440 13322 7449
rect 13266 7375 13322 7384
rect 13280 6458 13308 7375
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 12584 5664 12664 5692
rect 12532 5646 12584 5652
rect 12070 5607 12126 5616
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 12544 5234 12572 5646
rect 12912 5234 12940 6122
rect 13280 5914 13308 6394
rect 13372 6254 13400 6734
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13372 5846 13400 6190
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 12992 5636 13044 5642
rect 12992 5578 13044 5584
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12214 4924 12522 4944
rect 12214 4922 12220 4924
rect 12276 4922 12300 4924
rect 12356 4922 12380 4924
rect 12436 4922 12460 4924
rect 12516 4922 12522 4924
rect 12276 4870 12278 4922
rect 12458 4870 12460 4922
rect 12214 4868 12220 4870
rect 12276 4868 12300 4870
rect 12356 4868 12380 4870
rect 12436 4868 12460 4870
rect 12516 4868 12522 4870
rect 12214 4848 12522 4868
rect 12912 4622 12940 5170
rect 13004 5098 13032 5578
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 12992 5092 13044 5098
rect 12992 5034 13044 5040
rect 13004 4622 13032 5034
rect 13188 4758 13216 5510
rect 13372 4826 13400 5782
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13176 4752 13228 4758
rect 13176 4694 13228 4700
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 13280 4146 13308 4422
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 11532 3534 11560 4014
rect 11704 4004 11756 4010
rect 11704 3946 11756 3952
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11256 2514 11284 2586
rect 11244 2508 11296 2514
rect 11244 2450 11296 2456
rect 11440 2446 11468 3402
rect 11532 2922 11560 3470
rect 11716 3466 11744 3946
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 11716 3126 11744 3402
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 11900 2990 11928 3878
rect 11992 3534 12020 4014
rect 12900 4004 12952 4010
rect 12900 3946 12952 3952
rect 12214 3836 12522 3856
rect 12214 3834 12220 3836
rect 12276 3834 12300 3836
rect 12356 3834 12380 3836
rect 12436 3834 12460 3836
rect 12516 3834 12522 3836
rect 12276 3782 12278 3834
rect 12458 3782 12460 3834
rect 12214 3780 12220 3782
rect 12276 3780 12300 3782
rect 12356 3780 12380 3782
rect 12436 3780 12460 3782
rect 12516 3780 12522 3782
rect 12214 3760 12522 3780
rect 12912 3670 12940 3946
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11992 3194 12020 3470
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 11888 2984 11940 2990
rect 12072 2984 12124 2990
rect 11888 2926 11940 2932
rect 11992 2944 12072 2972
rect 11520 2916 11572 2922
rect 11520 2858 11572 2864
rect 11992 2514 12020 2944
rect 12072 2926 12124 2932
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 11348 2106 11376 2382
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 11336 2100 11388 2106
rect 11336 2042 11388 2048
rect 11624 1834 11652 2314
rect 12084 2310 12112 2790
rect 12214 2748 12522 2768
rect 12214 2746 12220 2748
rect 12276 2746 12300 2748
rect 12356 2746 12380 2748
rect 12436 2746 12460 2748
rect 12516 2746 12522 2748
rect 12276 2694 12278 2746
rect 12458 2694 12460 2746
rect 12214 2692 12220 2694
rect 12276 2692 12300 2694
rect 12356 2692 12380 2694
rect 12436 2692 12460 2694
rect 12516 2692 12522 2694
rect 12214 2672 12522 2692
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 11612 1828 11664 1834
rect 11612 1770 11664 1776
rect 12084 1442 12112 2246
rect 12214 1660 12522 1680
rect 12214 1658 12220 1660
rect 12276 1658 12300 1660
rect 12356 1658 12380 1660
rect 12436 1658 12460 1660
rect 12516 1658 12522 1660
rect 12276 1606 12278 1658
rect 12458 1606 12460 1658
rect 12214 1604 12220 1606
rect 12276 1604 12300 1606
rect 12356 1604 12380 1606
rect 12436 1604 12460 1606
rect 12516 1604 12522 1606
rect 12214 1584 12522 1604
rect 11060 1420 11112 1426
rect 12084 1414 12204 1442
rect 11060 1362 11112 1368
rect 11704 1352 11756 1358
rect 11702 1320 11704 1329
rect 11756 1320 11758 1329
rect 11702 1255 11758 1264
rect 12176 800 12204 1414
rect 12636 1358 12664 2246
rect 12912 2038 12940 3606
rect 13004 3194 13032 4014
rect 13280 3534 13308 4082
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13084 2372 13136 2378
rect 13084 2314 13136 2320
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12900 2032 12952 2038
rect 12900 1974 12952 1980
rect 13096 1358 13124 2314
rect 13280 1562 13308 2314
rect 13360 1896 13412 1902
rect 13360 1838 13412 1844
rect 13268 1556 13320 1562
rect 13268 1498 13320 1504
rect 13372 1358 13400 1838
rect 14004 1420 14056 1426
rect 14004 1362 14056 1368
rect 12624 1352 12676 1358
rect 12624 1294 12676 1300
rect 13084 1352 13136 1358
rect 13084 1294 13136 1300
rect 13360 1352 13412 1358
rect 13360 1294 13412 1300
rect 14016 800 14044 1362
rect 10336 734 11008 762
rect 12162 0 12218 800
rect 13912 536 13964 542
rect 13910 504 13912 513
rect 13964 504 13966 513
rect 13910 439 13966 448
rect 14002 0 14058 800
<< via2 >>
rect 10874 14456 10930 14512
rect 1490 11192 1546 11248
rect 2594 10920 2650 10976
rect 2686 10648 2742 10704
rect 2410 10376 2466 10432
rect 3054 10784 3110 10840
rect 2870 10668 2926 10704
rect 2870 10648 2872 10668
rect 2872 10648 2924 10668
rect 2924 10648 2926 10668
rect 3238 10920 3294 10976
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4342 11756 4398 11792
rect 4342 11736 4344 11756
rect 4344 11736 4396 11756
rect 4396 11736 4398 11756
rect 4710 11736 4766 11792
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 3790 10376 3846 10432
rect 8220 13082 8276 13084
rect 8300 13082 8356 13084
rect 8380 13082 8436 13084
rect 8460 13082 8516 13084
rect 8220 13030 8266 13082
rect 8266 13030 8276 13082
rect 8300 13030 8330 13082
rect 8330 13030 8342 13082
rect 8342 13030 8356 13082
rect 8380 13030 8394 13082
rect 8394 13030 8406 13082
rect 8406 13030 8436 13082
rect 8460 13030 8470 13082
rect 8470 13030 8516 13082
rect 8220 13028 8276 13030
rect 8300 13028 8356 13030
rect 8380 13028 8436 13030
rect 8460 13028 8516 13030
rect 5630 11736 5686 11792
rect 4526 10668 4582 10704
rect 4526 10648 4528 10668
rect 4528 10648 4580 10668
rect 4580 10648 4582 10668
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4710 10784 4766 10840
rect 8220 11994 8276 11996
rect 8300 11994 8356 11996
rect 8380 11994 8436 11996
rect 8460 11994 8516 11996
rect 8220 11942 8266 11994
rect 8266 11942 8276 11994
rect 8300 11942 8330 11994
rect 8330 11942 8342 11994
rect 8342 11942 8356 11994
rect 8380 11942 8394 11994
rect 8394 11942 8406 11994
rect 8406 11942 8436 11994
rect 8460 11942 8470 11994
rect 8470 11942 8516 11994
rect 8220 11940 8276 11942
rect 8300 11940 8356 11942
rect 8380 11940 8436 11942
rect 8460 11940 8516 11942
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 1582 3732 1638 3768
rect 1582 3712 1584 3732
rect 1584 3712 1636 3732
rect 1636 3712 1638 3732
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3606 6432 3662 6488
rect 3422 6316 3478 6352
rect 3422 6296 3424 6316
rect 3424 6296 3476 6316
rect 3476 6296 3478 6316
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4526 5752 4582 5808
rect 4894 6452 4950 6488
rect 4894 6432 4896 6452
rect 4896 6432 4948 6452
rect 4948 6432 4950 6452
rect 4894 6296 4950 6352
rect 4710 5652 4712 5672
rect 4712 5652 4764 5672
rect 4764 5652 4766 5672
rect 4710 5616 4766 5652
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 5170 6860 5226 6896
rect 8220 10906 8276 10908
rect 8300 10906 8356 10908
rect 8380 10906 8436 10908
rect 8460 10906 8516 10908
rect 8220 10854 8266 10906
rect 8266 10854 8276 10906
rect 8300 10854 8330 10906
rect 8330 10854 8342 10906
rect 8342 10854 8356 10906
rect 8380 10854 8394 10906
rect 8394 10854 8406 10906
rect 8406 10854 8436 10906
rect 8460 10854 8470 10906
rect 8470 10854 8516 10906
rect 8220 10852 8276 10854
rect 8300 10852 8356 10854
rect 8380 10852 8436 10854
rect 8460 10852 8516 10854
rect 5170 6840 5172 6860
rect 5172 6840 5224 6860
rect 5224 6840 5226 6860
rect 5354 6316 5410 6352
rect 5354 6296 5356 6316
rect 5356 6296 5408 6316
rect 5408 6296 5410 6316
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 7286 6840 7342 6896
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4220 1658 4276 1660
rect 4300 1658 4356 1660
rect 4380 1658 4436 1660
rect 4460 1658 4516 1660
rect 4220 1606 4266 1658
rect 4266 1606 4276 1658
rect 4300 1606 4330 1658
rect 4330 1606 4342 1658
rect 4342 1606 4356 1658
rect 4380 1606 4394 1658
rect 4394 1606 4406 1658
rect 4406 1606 4436 1658
rect 4460 1606 4470 1658
rect 4470 1606 4516 1658
rect 4220 1604 4276 1606
rect 4300 1604 4356 1606
rect 4380 1604 4436 1606
rect 4460 1604 4516 1606
rect 7102 5752 7158 5808
rect 7194 4564 7196 4584
rect 7196 4564 7248 4584
rect 7248 4564 7250 4584
rect 7194 4528 7250 4564
rect 8220 9818 8276 9820
rect 8300 9818 8356 9820
rect 8380 9818 8436 9820
rect 8460 9818 8516 9820
rect 8220 9766 8266 9818
rect 8266 9766 8276 9818
rect 8300 9766 8330 9818
rect 8330 9766 8342 9818
rect 8342 9766 8356 9818
rect 8380 9766 8394 9818
rect 8394 9766 8406 9818
rect 8406 9766 8436 9818
rect 8460 9766 8470 9818
rect 8470 9766 8516 9818
rect 8220 9764 8276 9766
rect 8300 9764 8356 9766
rect 8380 9764 8436 9766
rect 8460 9764 8516 9766
rect 8220 8730 8276 8732
rect 8300 8730 8356 8732
rect 8380 8730 8436 8732
rect 8460 8730 8516 8732
rect 8220 8678 8266 8730
rect 8266 8678 8276 8730
rect 8300 8678 8330 8730
rect 8330 8678 8342 8730
rect 8342 8678 8356 8730
rect 8380 8678 8394 8730
rect 8394 8678 8406 8730
rect 8406 8678 8436 8730
rect 8460 8678 8470 8730
rect 8470 8678 8516 8730
rect 8220 8676 8276 8678
rect 8300 8676 8356 8678
rect 8380 8676 8436 8678
rect 8460 8676 8516 8678
rect 8220 7642 8276 7644
rect 8300 7642 8356 7644
rect 8380 7642 8436 7644
rect 8460 7642 8516 7644
rect 8220 7590 8266 7642
rect 8266 7590 8276 7642
rect 8300 7590 8330 7642
rect 8330 7590 8342 7642
rect 8342 7590 8356 7642
rect 8380 7590 8394 7642
rect 8394 7590 8406 7642
rect 8406 7590 8436 7642
rect 8460 7590 8470 7642
rect 8470 7590 8516 7642
rect 8220 7588 8276 7590
rect 8300 7588 8356 7590
rect 8380 7588 8436 7590
rect 8460 7588 8516 7590
rect 7470 6160 7526 6216
rect 8220 6554 8276 6556
rect 8300 6554 8356 6556
rect 8380 6554 8436 6556
rect 8460 6554 8516 6556
rect 8220 6502 8266 6554
rect 8266 6502 8276 6554
rect 8300 6502 8330 6554
rect 8330 6502 8342 6554
rect 8342 6502 8356 6554
rect 8380 6502 8394 6554
rect 8394 6502 8406 6554
rect 8406 6502 8436 6554
rect 8460 6502 8470 6554
rect 8470 6502 8516 6554
rect 8220 6500 8276 6502
rect 8300 6500 8356 6502
rect 8380 6500 8436 6502
rect 8460 6500 8516 6502
rect 7562 5616 7618 5672
rect 10046 13368 10102 13424
rect 8666 5480 8722 5536
rect 8220 5466 8276 5468
rect 8300 5466 8356 5468
rect 8380 5466 8436 5468
rect 8460 5466 8516 5468
rect 8220 5414 8266 5466
rect 8266 5414 8276 5466
rect 8300 5414 8330 5466
rect 8330 5414 8342 5466
rect 8342 5414 8356 5466
rect 8380 5414 8394 5466
rect 8394 5414 8406 5466
rect 8406 5414 8436 5466
rect 8460 5414 8470 5466
rect 8470 5414 8516 5466
rect 8220 5412 8276 5414
rect 8300 5412 8356 5414
rect 8380 5412 8436 5414
rect 8460 5412 8516 5414
rect 7838 4548 7894 4584
rect 7838 4528 7840 4548
rect 7840 4528 7892 4548
rect 7892 4528 7894 4548
rect 8574 4564 8576 4584
rect 8576 4564 8628 4584
rect 8628 4564 8630 4584
rect 8574 4528 8630 4564
rect 8220 4378 8276 4380
rect 8300 4378 8356 4380
rect 8380 4378 8436 4380
rect 8460 4378 8516 4380
rect 8220 4326 8266 4378
rect 8266 4326 8276 4378
rect 8300 4326 8330 4378
rect 8330 4326 8342 4378
rect 8342 4326 8356 4378
rect 8380 4326 8394 4378
rect 8394 4326 8406 4378
rect 8406 4326 8436 4378
rect 8460 4326 8470 4378
rect 8470 4326 8516 4378
rect 8220 4324 8276 4326
rect 8300 4324 8356 4326
rect 8380 4324 8436 4326
rect 8460 4324 8516 4326
rect 8942 5072 8998 5128
rect 8220 3290 8276 3292
rect 8300 3290 8356 3292
rect 8380 3290 8436 3292
rect 8460 3290 8516 3292
rect 8220 3238 8266 3290
rect 8266 3238 8276 3290
rect 8300 3238 8330 3290
rect 8330 3238 8342 3290
rect 8342 3238 8356 3290
rect 8380 3238 8394 3290
rect 8394 3238 8406 3290
rect 8406 3238 8436 3290
rect 8460 3238 8470 3290
rect 8470 3238 8516 3290
rect 8220 3236 8276 3238
rect 8300 3236 8356 3238
rect 8380 3236 8436 3238
rect 8460 3236 8516 3238
rect 8220 2202 8276 2204
rect 8300 2202 8356 2204
rect 8380 2202 8436 2204
rect 8460 2202 8516 2204
rect 8220 2150 8266 2202
rect 8266 2150 8276 2202
rect 8300 2150 8330 2202
rect 8330 2150 8342 2202
rect 8342 2150 8356 2202
rect 8380 2150 8394 2202
rect 8394 2150 8406 2202
rect 8406 2150 8436 2202
rect 8460 2150 8470 2202
rect 8470 2150 8516 2202
rect 8220 2148 8276 2150
rect 8300 2148 8356 2150
rect 8380 2148 8436 2150
rect 8460 2148 8516 2150
rect 8220 1114 8276 1116
rect 8300 1114 8356 1116
rect 8380 1114 8436 1116
rect 8460 1114 8516 1116
rect 8220 1062 8266 1114
rect 8266 1062 8276 1114
rect 8300 1062 8330 1114
rect 8330 1062 8342 1114
rect 8342 1062 8356 1114
rect 8380 1062 8394 1114
rect 8394 1062 8406 1114
rect 8406 1062 8436 1114
rect 8460 1062 8470 1114
rect 8470 1062 8516 1114
rect 8220 1060 8276 1062
rect 8300 1060 8356 1062
rect 8380 1060 8436 1062
rect 8460 1060 8516 1062
rect 9310 5888 9366 5944
rect 9310 5652 9312 5672
rect 9312 5652 9364 5672
rect 9364 5652 9366 5672
rect 9310 5616 9366 5652
rect 9310 5072 9366 5128
rect 10782 12688 10838 12744
rect 10322 10920 10378 10976
rect 10506 10104 10562 10160
rect 10414 9016 10470 9072
rect 9494 6196 9496 6216
rect 9496 6196 9548 6216
rect 9548 6196 9550 6216
rect 9494 6160 9550 6196
rect 9586 5208 9642 5264
rect 9494 3984 9550 4040
rect 8758 3304 8814 3360
rect 10138 5616 10194 5672
rect 10046 5072 10102 5128
rect 9954 4800 10010 4856
rect 9402 3168 9458 3224
rect 9586 3032 9642 3088
rect 10506 5228 10562 5264
rect 10506 5208 10508 5228
rect 10508 5208 10560 5228
rect 10560 5208 10562 5228
rect 10414 4548 10470 4584
rect 10414 4528 10416 4548
rect 10416 4528 10468 4548
rect 10468 4528 10470 4548
rect 10414 3304 10470 3360
rect 12220 13626 12276 13628
rect 12300 13626 12356 13628
rect 12380 13626 12436 13628
rect 12460 13626 12516 13628
rect 12220 13574 12266 13626
rect 12266 13574 12276 13626
rect 12300 13574 12330 13626
rect 12330 13574 12342 13626
rect 12342 13574 12356 13626
rect 12380 13574 12394 13626
rect 12394 13574 12406 13626
rect 12406 13574 12436 13626
rect 12460 13574 12470 13626
rect 12470 13574 12516 13626
rect 12220 13572 12276 13574
rect 12300 13572 12356 13574
rect 12380 13572 12436 13574
rect 12460 13572 12516 13574
rect 12220 12538 12276 12540
rect 12300 12538 12356 12540
rect 12380 12538 12436 12540
rect 12460 12538 12516 12540
rect 12220 12486 12266 12538
rect 12266 12486 12276 12538
rect 12300 12486 12330 12538
rect 12330 12486 12342 12538
rect 12342 12486 12356 12538
rect 12380 12486 12394 12538
rect 12394 12486 12406 12538
rect 12406 12486 12436 12538
rect 12460 12486 12470 12538
rect 12470 12486 12516 12538
rect 12220 12484 12276 12486
rect 12300 12484 12356 12486
rect 12380 12484 12436 12486
rect 12460 12484 12516 12486
rect 11610 11872 11666 11928
rect 12220 11450 12276 11452
rect 12300 11450 12356 11452
rect 12380 11450 12436 11452
rect 12460 11450 12516 11452
rect 12220 11398 12266 11450
rect 12266 11398 12276 11450
rect 12300 11398 12330 11450
rect 12330 11398 12342 11450
rect 12342 11398 12356 11450
rect 12380 11398 12394 11450
rect 12394 11398 12406 11450
rect 12406 11398 12436 11450
rect 12460 11398 12470 11450
rect 12470 11398 12516 11450
rect 12220 11396 12276 11398
rect 12300 11396 12356 11398
rect 12380 11396 12436 11398
rect 12460 11396 12516 11398
rect 12220 10362 12276 10364
rect 12300 10362 12356 10364
rect 12380 10362 12436 10364
rect 12460 10362 12516 10364
rect 12220 10310 12266 10362
rect 12266 10310 12276 10362
rect 12300 10310 12330 10362
rect 12330 10310 12342 10362
rect 12342 10310 12356 10362
rect 12380 10310 12394 10362
rect 12394 10310 12406 10362
rect 12406 10310 12436 10362
rect 12460 10310 12470 10362
rect 12470 10310 12516 10362
rect 12220 10308 12276 10310
rect 12300 10308 12356 10310
rect 12380 10308 12436 10310
rect 12460 10308 12516 10310
rect 11334 6568 11390 6624
rect 10874 6196 10876 6216
rect 10876 6196 10928 6216
rect 10928 6196 10930 6216
rect 10874 6160 10930 6196
rect 12220 9274 12276 9276
rect 12300 9274 12356 9276
rect 12380 9274 12436 9276
rect 12460 9274 12516 9276
rect 12220 9222 12266 9274
rect 12266 9222 12276 9274
rect 12300 9222 12330 9274
rect 12330 9222 12342 9274
rect 12342 9222 12356 9274
rect 12380 9222 12394 9274
rect 12394 9222 12406 9274
rect 12406 9222 12436 9274
rect 12460 9222 12470 9274
rect 12470 9222 12516 9274
rect 12220 9220 12276 9222
rect 12300 9220 12356 9222
rect 12380 9220 12436 9222
rect 12460 9220 12516 9222
rect 12220 8186 12276 8188
rect 12300 8186 12356 8188
rect 12380 8186 12436 8188
rect 12460 8186 12516 8188
rect 12220 8134 12266 8186
rect 12266 8134 12276 8186
rect 12300 8134 12330 8186
rect 12330 8134 12342 8186
rect 12342 8134 12356 8186
rect 12380 8134 12394 8186
rect 12394 8134 12406 8186
rect 12406 8134 12436 8186
rect 12460 8134 12470 8186
rect 12470 8134 12516 8186
rect 12220 8132 12276 8134
rect 12300 8132 12356 8134
rect 12380 8132 12436 8134
rect 12460 8132 12516 8134
rect 12220 7098 12276 7100
rect 12300 7098 12356 7100
rect 12380 7098 12436 7100
rect 12460 7098 12516 7100
rect 12220 7046 12266 7098
rect 12266 7046 12276 7098
rect 12300 7046 12330 7098
rect 12330 7046 12342 7098
rect 12342 7046 12356 7098
rect 12380 7046 12394 7098
rect 12394 7046 12406 7098
rect 12406 7046 12436 7098
rect 12460 7046 12470 7098
rect 12470 7046 12516 7098
rect 12220 7044 12276 7046
rect 12300 7044 12356 7046
rect 12380 7044 12436 7046
rect 12460 7044 12516 7046
rect 10690 5228 10746 5264
rect 10690 5208 10692 5228
rect 10692 5208 10744 5228
rect 10744 5208 10746 5228
rect 10966 5208 11022 5264
rect 11058 3304 11114 3360
rect 10690 2080 10746 2136
rect 11426 4800 11482 4856
rect 11978 6196 11980 6216
rect 11980 6196 12032 6216
rect 12032 6196 12034 6216
rect 11978 6160 12034 6196
rect 12220 6010 12276 6012
rect 12300 6010 12356 6012
rect 12380 6010 12436 6012
rect 12460 6010 12516 6012
rect 12220 5958 12266 6010
rect 12266 5958 12276 6010
rect 12300 5958 12330 6010
rect 12330 5958 12342 6010
rect 12342 5958 12356 6010
rect 12380 5958 12394 6010
rect 12394 5958 12406 6010
rect 12406 5958 12436 6010
rect 12460 5958 12470 6010
rect 12470 5958 12516 6010
rect 12220 5956 12276 5958
rect 12300 5956 12356 5958
rect 12380 5956 12436 5958
rect 12460 5956 12516 5958
rect 12070 5616 12126 5672
rect 13266 8372 13268 8392
rect 13268 8372 13320 8392
rect 13320 8372 13322 8392
rect 13266 8336 13322 8372
rect 13266 7384 13322 7440
rect 12220 4922 12276 4924
rect 12300 4922 12356 4924
rect 12380 4922 12436 4924
rect 12460 4922 12516 4924
rect 12220 4870 12266 4922
rect 12266 4870 12276 4922
rect 12300 4870 12330 4922
rect 12330 4870 12342 4922
rect 12342 4870 12356 4922
rect 12380 4870 12394 4922
rect 12394 4870 12406 4922
rect 12406 4870 12436 4922
rect 12460 4870 12470 4922
rect 12470 4870 12516 4922
rect 12220 4868 12276 4870
rect 12300 4868 12356 4870
rect 12380 4868 12436 4870
rect 12460 4868 12516 4870
rect 12220 3834 12276 3836
rect 12300 3834 12356 3836
rect 12380 3834 12436 3836
rect 12460 3834 12516 3836
rect 12220 3782 12266 3834
rect 12266 3782 12276 3834
rect 12300 3782 12330 3834
rect 12330 3782 12342 3834
rect 12342 3782 12356 3834
rect 12380 3782 12394 3834
rect 12394 3782 12406 3834
rect 12406 3782 12436 3834
rect 12460 3782 12470 3834
rect 12470 3782 12516 3834
rect 12220 3780 12276 3782
rect 12300 3780 12356 3782
rect 12380 3780 12436 3782
rect 12460 3780 12516 3782
rect 12220 2746 12276 2748
rect 12300 2746 12356 2748
rect 12380 2746 12436 2748
rect 12460 2746 12516 2748
rect 12220 2694 12266 2746
rect 12266 2694 12276 2746
rect 12300 2694 12330 2746
rect 12330 2694 12342 2746
rect 12342 2694 12356 2746
rect 12380 2694 12394 2746
rect 12394 2694 12406 2746
rect 12406 2694 12436 2746
rect 12460 2694 12470 2746
rect 12470 2694 12516 2746
rect 12220 2692 12276 2694
rect 12300 2692 12356 2694
rect 12380 2692 12436 2694
rect 12460 2692 12516 2694
rect 12220 1658 12276 1660
rect 12300 1658 12356 1660
rect 12380 1658 12436 1660
rect 12460 1658 12516 1660
rect 12220 1606 12266 1658
rect 12266 1606 12276 1658
rect 12300 1606 12330 1658
rect 12330 1606 12342 1658
rect 12342 1606 12356 1658
rect 12380 1606 12394 1658
rect 12394 1606 12406 1658
rect 12406 1606 12436 1658
rect 12460 1606 12470 1658
rect 12470 1606 12516 1658
rect 12220 1604 12276 1606
rect 12300 1604 12356 1606
rect 12380 1604 12436 1606
rect 12460 1604 12516 1606
rect 11702 1300 11704 1320
rect 11704 1300 11756 1320
rect 11756 1300 11758 1320
rect 11702 1264 11758 1300
rect 13910 484 13912 504
rect 13912 484 13964 504
rect 13964 484 13966 504
rect 13910 448 13966 484
<< metal3 >>
rect 10869 14514 10935 14517
rect 14200 14514 15000 14544
rect 10869 14512 15000 14514
rect 10869 14456 10874 14512
rect 10930 14456 15000 14512
rect 10869 14454 15000 14456
rect 10869 14451 10935 14454
rect 14200 14424 15000 14454
rect 14200 13698 15000 13728
rect 12758 13638 15000 13698
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 12208 13632 12528 13633
rect 12208 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12528 13632
rect 12208 13567 12528 13568
rect 10041 13426 10107 13429
rect 12758 13426 12818 13638
rect 14200 13608 15000 13638
rect 10041 13424 12818 13426
rect 10041 13368 10046 13424
rect 10102 13368 12818 13424
rect 10041 13366 12818 13368
rect 10041 13363 10107 13366
rect 8208 13088 8528 13089
rect 8208 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8528 13088
rect 8208 13023 8528 13024
rect 10777 12746 10843 12749
rect 14200 12746 15000 12776
rect 10777 12744 15000 12746
rect 10777 12688 10782 12744
rect 10838 12688 15000 12744
rect 10777 12686 15000 12688
rect 10777 12683 10843 12686
rect 14200 12656 15000 12686
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 12208 12544 12528 12545
rect 12208 12480 12216 12544
rect 12280 12480 12296 12544
rect 12360 12480 12376 12544
rect 12440 12480 12456 12544
rect 12520 12480 12528 12544
rect 12208 12479 12528 12480
rect 8208 12000 8528 12001
rect 8208 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8528 12000
rect 8208 11935 8528 11936
rect 11605 11930 11671 11933
rect 14200 11930 15000 11960
rect 11605 11928 15000 11930
rect 11605 11872 11610 11928
rect 11666 11872 15000 11928
rect 11605 11870 15000 11872
rect 11605 11867 11671 11870
rect 14200 11840 15000 11870
rect 4337 11794 4403 11797
rect 4705 11794 4771 11797
rect 5625 11794 5691 11797
rect 4337 11792 5691 11794
rect 4337 11736 4342 11792
rect 4398 11736 4710 11792
rect 4766 11736 5630 11792
rect 5686 11736 5691 11792
rect 4337 11734 5691 11736
rect 4337 11731 4403 11734
rect 4705 11731 4771 11734
rect 5625 11731 5691 11734
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 12208 11456 12528 11457
rect 12208 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12528 11456
rect 12208 11391 12528 11392
rect 0 11250 800 11280
rect 1485 11250 1551 11253
rect 0 11248 1551 11250
rect 0 11192 1490 11248
rect 1546 11192 1551 11248
rect 0 11190 1551 11192
rect 0 11160 800 11190
rect 1485 11187 1551 11190
rect 2589 10978 2655 10981
rect 3233 10978 3299 10981
rect 2589 10976 3299 10978
rect 2589 10920 2594 10976
rect 2650 10920 3238 10976
rect 3294 10920 3299 10976
rect 2589 10918 3299 10920
rect 2589 10915 2655 10918
rect 3233 10915 3299 10918
rect 10317 10978 10383 10981
rect 14200 10978 15000 11008
rect 10317 10976 15000 10978
rect 10317 10920 10322 10976
rect 10378 10920 15000 10976
rect 10317 10918 15000 10920
rect 10317 10915 10383 10918
rect 8208 10912 8528 10913
rect 8208 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8528 10912
rect 14200 10888 15000 10918
rect 8208 10847 8528 10848
rect 3049 10842 3115 10845
rect 4705 10842 4771 10845
rect 3049 10840 4771 10842
rect 3049 10784 3054 10840
rect 3110 10784 4710 10840
rect 4766 10784 4771 10840
rect 3049 10782 4771 10784
rect 3049 10779 3115 10782
rect 4705 10779 4771 10782
rect 2681 10706 2747 10709
rect 2865 10706 2931 10709
rect 4521 10706 4587 10709
rect 2681 10704 4587 10706
rect 2681 10648 2686 10704
rect 2742 10648 2870 10704
rect 2926 10648 4526 10704
rect 4582 10648 4587 10704
rect 2681 10646 4587 10648
rect 2681 10643 2747 10646
rect 2865 10643 2931 10646
rect 4521 10643 4587 10646
rect 2405 10434 2471 10437
rect 3785 10434 3851 10437
rect 2405 10432 3851 10434
rect 2405 10376 2410 10432
rect 2466 10376 3790 10432
rect 3846 10376 3851 10432
rect 2405 10374 3851 10376
rect 2405 10371 2471 10374
rect 3785 10371 3851 10374
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 12208 10368 12528 10369
rect 12208 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12528 10368
rect 12208 10303 12528 10304
rect 10501 10162 10567 10165
rect 14200 10162 15000 10192
rect 10501 10160 15000 10162
rect 10501 10104 10506 10160
rect 10562 10104 15000 10160
rect 10501 10102 15000 10104
rect 10501 10099 10567 10102
rect 14200 10072 15000 10102
rect 8208 9824 8528 9825
rect 8208 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8528 9824
rect 8208 9759 8528 9760
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 12208 9280 12528 9281
rect 12208 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12528 9280
rect 12208 9215 12528 9216
rect 14200 9210 15000 9240
rect 12758 9150 15000 9210
rect 10409 9074 10475 9077
rect 12758 9074 12818 9150
rect 14200 9120 15000 9150
rect 10409 9072 12818 9074
rect 10409 9016 10414 9072
rect 10470 9016 12818 9072
rect 10409 9014 12818 9016
rect 10409 9011 10475 9014
rect 8208 8736 8528 8737
rect 8208 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8528 8736
rect 8208 8671 8528 8672
rect 13261 8394 13327 8397
rect 14200 8394 15000 8424
rect 13261 8392 15000 8394
rect 13261 8336 13266 8392
rect 13322 8336 15000 8392
rect 13261 8334 15000 8336
rect 13261 8331 13327 8334
rect 14200 8304 15000 8334
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 12208 8192 12528 8193
rect 12208 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12528 8192
rect 12208 8127 12528 8128
rect 8208 7648 8528 7649
rect 8208 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8528 7648
rect 8208 7583 8528 7584
rect 13261 7442 13327 7445
rect 14200 7442 15000 7472
rect 13261 7440 15000 7442
rect 13261 7384 13266 7440
rect 13322 7384 15000 7440
rect 13261 7382 15000 7384
rect 13261 7379 13327 7382
rect 14200 7352 15000 7382
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 12208 7104 12528 7105
rect 12208 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12528 7104
rect 12208 7039 12528 7040
rect 5165 6898 5231 6901
rect 7281 6898 7347 6901
rect 5165 6896 7347 6898
rect 5165 6840 5170 6896
rect 5226 6840 7286 6896
rect 7342 6840 7347 6896
rect 5165 6838 7347 6840
rect 5165 6835 5231 6838
rect 7281 6835 7347 6838
rect 11329 6626 11395 6629
rect 14200 6626 15000 6656
rect 11329 6624 15000 6626
rect 11329 6568 11334 6624
rect 11390 6568 15000 6624
rect 11329 6566 15000 6568
rect 11329 6563 11395 6566
rect 8208 6560 8528 6561
rect 8208 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8528 6560
rect 14200 6536 15000 6566
rect 8208 6495 8528 6496
rect 3601 6490 3667 6493
rect 4889 6490 4955 6493
rect 3601 6488 4955 6490
rect 3601 6432 3606 6488
rect 3662 6432 4894 6488
rect 4950 6432 4955 6488
rect 3601 6430 4955 6432
rect 3601 6427 3667 6430
rect 4889 6427 4955 6430
rect 3417 6354 3483 6357
rect 4889 6354 4955 6357
rect 5349 6354 5415 6357
rect 3417 6352 5415 6354
rect 3417 6296 3422 6352
rect 3478 6296 4894 6352
rect 4950 6296 5354 6352
rect 5410 6296 5415 6352
rect 3417 6294 5415 6296
rect 3417 6291 3483 6294
rect 4889 6291 4955 6294
rect 5349 6291 5415 6294
rect 7465 6218 7531 6221
rect 9489 6218 9555 6221
rect 7465 6216 9555 6218
rect 7465 6160 7470 6216
rect 7526 6160 9494 6216
rect 9550 6160 9555 6216
rect 7465 6158 9555 6160
rect 7465 6155 7531 6158
rect 9489 6155 9555 6158
rect 10869 6218 10935 6221
rect 11973 6218 12039 6221
rect 10869 6216 12039 6218
rect 10869 6160 10874 6216
rect 10930 6160 11978 6216
rect 12034 6160 12039 6216
rect 10869 6158 12039 6160
rect 10869 6155 10935 6158
rect 11973 6155 12039 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 12208 6016 12528 6017
rect 12208 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12528 6016
rect 12208 5951 12528 5952
rect 9305 5948 9371 5949
rect 9254 5884 9260 5948
rect 9324 5946 9371 5948
rect 9324 5944 9416 5946
rect 9366 5888 9416 5944
rect 9324 5886 9416 5888
rect 9324 5884 9371 5886
rect 9305 5883 9371 5884
rect 4521 5810 4587 5813
rect 7097 5810 7163 5813
rect 4521 5808 7163 5810
rect 4521 5752 4526 5808
rect 4582 5752 7102 5808
rect 7158 5752 7163 5808
rect 4521 5750 7163 5752
rect 4521 5747 4587 5750
rect 7097 5747 7163 5750
rect 4705 5674 4771 5677
rect 7557 5674 7623 5677
rect 9305 5674 9371 5677
rect 4705 5672 9371 5674
rect 4705 5616 4710 5672
rect 4766 5616 7562 5672
rect 7618 5616 9310 5672
rect 9366 5616 9371 5672
rect 4705 5614 9371 5616
rect 4705 5611 4771 5614
rect 7557 5611 7623 5614
rect 9305 5611 9371 5614
rect 10133 5672 10199 5677
rect 10133 5616 10138 5672
rect 10194 5616 10199 5672
rect 10133 5611 10199 5616
rect 12065 5674 12131 5677
rect 14200 5674 15000 5704
rect 12065 5672 15000 5674
rect 12065 5616 12070 5672
rect 12126 5616 15000 5672
rect 12065 5614 15000 5616
rect 12065 5611 12131 5614
rect 8661 5538 8727 5541
rect 10136 5538 10196 5611
rect 14200 5584 15000 5614
rect 8661 5536 10196 5538
rect 8661 5480 8666 5536
rect 8722 5480 10196 5536
rect 8661 5478 10196 5480
rect 8661 5475 8727 5478
rect 8208 5472 8528 5473
rect 8208 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8528 5472
rect 8208 5407 8528 5408
rect 9581 5266 9647 5269
rect 10501 5266 10567 5269
rect 9581 5264 10567 5266
rect 9581 5208 9586 5264
rect 9642 5208 10506 5264
rect 10562 5208 10567 5264
rect 9581 5206 10567 5208
rect 9581 5203 9647 5206
rect 10501 5203 10567 5206
rect 10685 5266 10751 5269
rect 10961 5266 11027 5269
rect 10685 5264 11027 5266
rect 10685 5208 10690 5264
rect 10746 5208 10966 5264
rect 11022 5208 11027 5264
rect 10685 5206 11027 5208
rect 10685 5203 10751 5206
rect 10961 5203 11027 5206
rect 8937 5130 9003 5133
rect 9305 5130 9371 5133
rect 8937 5128 9371 5130
rect 8937 5072 8942 5128
rect 8998 5072 9310 5128
rect 9366 5072 9371 5128
rect 8937 5070 9371 5072
rect 8937 5067 9003 5070
rect 9305 5067 9371 5070
rect 10041 5130 10107 5133
rect 10041 5128 12818 5130
rect 10041 5072 10046 5128
rect 10102 5072 12818 5128
rect 10041 5070 12818 5072
rect 10041 5067 10107 5070
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 12208 4928 12528 4929
rect 12208 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12528 4928
rect 12208 4863 12528 4864
rect 9949 4858 10015 4861
rect 11421 4858 11487 4861
rect 9949 4856 11487 4858
rect 9949 4800 9954 4856
rect 10010 4800 11426 4856
rect 11482 4800 11487 4856
rect 9949 4798 11487 4800
rect 12758 4858 12818 5070
rect 14200 4858 15000 4888
rect 12758 4798 15000 4858
rect 9949 4795 10015 4798
rect 11421 4795 11487 4798
rect 14200 4768 15000 4798
rect 7189 4586 7255 4589
rect 7833 4586 7899 4589
rect 7189 4584 7899 4586
rect 7189 4528 7194 4584
rect 7250 4528 7838 4584
rect 7894 4528 7899 4584
rect 7189 4526 7899 4528
rect 7189 4523 7255 4526
rect 7833 4523 7899 4526
rect 8569 4586 8635 4589
rect 10409 4586 10475 4589
rect 8569 4584 10475 4586
rect 8569 4528 8574 4584
rect 8630 4528 10414 4584
rect 10470 4528 10475 4584
rect 8569 4526 10475 4528
rect 8569 4523 8635 4526
rect 10409 4523 10475 4526
rect 8208 4384 8528 4385
rect 8208 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8528 4384
rect 8208 4319 8528 4320
rect 9489 4042 9555 4045
rect 9489 4040 12818 4042
rect 9489 3984 9494 4040
rect 9550 3984 12818 4040
rect 9489 3982 12818 3984
rect 9489 3979 9555 3982
rect 12758 3906 12818 3982
rect 14200 3906 15000 3936
rect 12758 3846 15000 3906
rect 4208 3840 4528 3841
rect 0 3770 800 3800
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 12208 3840 12528 3841
rect 12208 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12528 3840
rect 14200 3816 15000 3846
rect 12208 3775 12528 3776
rect 1577 3770 1643 3773
rect 0 3768 1643 3770
rect 0 3712 1582 3768
rect 1638 3712 1643 3768
rect 0 3710 1643 3712
rect 0 3680 800 3710
rect 1577 3707 1643 3710
rect 8753 3362 8819 3365
rect 10409 3362 10475 3365
rect 11053 3362 11119 3365
rect 8753 3360 11119 3362
rect 8753 3304 8758 3360
rect 8814 3304 10414 3360
rect 10470 3304 11058 3360
rect 11114 3304 11119 3360
rect 8753 3302 11119 3304
rect 8753 3299 8819 3302
rect 10409 3299 10475 3302
rect 11053 3299 11119 3302
rect 8208 3296 8528 3297
rect 8208 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8528 3296
rect 8208 3231 8528 3232
rect 9254 3164 9260 3228
rect 9324 3226 9330 3228
rect 9397 3226 9463 3229
rect 9324 3224 9463 3226
rect 9324 3168 9402 3224
rect 9458 3168 9463 3224
rect 9324 3166 9463 3168
rect 9324 3164 9330 3166
rect 9397 3163 9463 3166
rect 9581 3090 9647 3093
rect 14200 3090 15000 3120
rect 9581 3088 15000 3090
rect 9581 3032 9586 3088
rect 9642 3032 15000 3088
rect 9581 3030 15000 3032
rect 9581 3027 9647 3030
rect 14200 3000 15000 3030
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 12208 2752 12528 2753
rect 12208 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12528 2752
rect 12208 2687 12528 2688
rect 8208 2208 8528 2209
rect 8208 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8528 2208
rect 8208 2143 8528 2144
rect 10685 2138 10751 2141
rect 14200 2138 15000 2168
rect 10685 2136 15000 2138
rect 10685 2080 10690 2136
rect 10746 2080 15000 2136
rect 10685 2078 15000 2080
rect 10685 2075 10751 2078
rect 14200 2048 15000 2078
rect 4208 1664 4528 1665
rect 4208 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4528 1664
rect 4208 1599 4528 1600
rect 12208 1664 12528 1665
rect 12208 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12528 1664
rect 12208 1599 12528 1600
rect 11697 1322 11763 1325
rect 14200 1322 15000 1352
rect 11697 1320 15000 1322
rect 11697 1264 11702 1320
rect 11758 1264 15000 1320
rect 11697 1262 15000 1264
rect 11697 1259 11763 1262
rect 14200 1232 15000 1262
rect 8208 1120 8528 1121
rect 8208 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8528 1120
rect 8208 1055 8528 1056
rect 13905 506 13971 509
rect 14200 506 15000 536
rect 13905 504 15000 506
rect 13905 448 13910 504
rect 13966 448 15000 504
rect 13905 446 15000 448
rect 13905 443 13971 446
rect 14200 416 15000 446
<< via3 >>
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 12216 13628 12280 13632
rect 12216 13572 12220 13628
rect 12220 13572 12276 13628
rect 12276 13572 12280 13628
rect 12216 13568 12280 13572
rect 12296 13628 12360 13632
rect 12296 13572 12300 13628
rect 12300 13572 12356 13628
rect 12356 13572 12360 13628
rect 12296 13568 12360 13572
rect 12376 13628 12440 13632
rect 12376 13572 12380 13628
rect 12380 13572 12436 13628
rect 12436 13572 12440 13628
rect 12376 13568 12440 13572
rect 12456 13628 12520 13632
rect 12456 13572 12460 13628
rect 12460 13572 12516 13628
rect 12516 13572 12520 13628
rect 12456 13568 12520 13572
rect 8216 13084 8280 13088
rect 8216 13028 8220 13084
rect 8220 13028 8276 13084
rect 8276 13028 8280 13084
rect 8216 13024 8280 13028
rect 8296 13084 8360 13088
rect 8296 13028 8300 13084
rect 8300 13028 8356 13084
rect 8356 13028 8360 13084
rect 8296 13024 8360 13028
rect 8376 13084 8440 13088
rect 8376 13028 8380 13084
rect 8380 13028 8436 13084
rect 8436 13028 8440 13084
rect 8376 13024 8440 13028
rect 8456 13084 8520 13088
rect 8456 13028 8460 13084
rect 8460 13028 8516 13084
rect 8516 13028 8520 13084
rect 8456 13024 8520 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 12216 12540 12280 12544
rect 12216 12484 12220 12540
rect 12220 12484 12276 12540
rect 12276 12484 12280 12540
rect 12216 12480 12280 12484
rect 12296 12540 12360 12544
rect 12296 12484 12300 12540
rect 12300 12484 12356 12540
rect 12356 12484 12360 12540
rect 12296 12480 12360 12484
rect 12376 12540 12440 12544
rect 12376 12484 12380 12540
rect 12380 12484 12436 12540
rect 12436 12484 12440 12540
rect 12376 12480 12440 12484
rect 12456 12540 12520 12544
rect 12456 12484 12460 12540
rect 12460 12484 12516 12540
rect 12516 12484 12520 12540
rect 12456 12480 12520 12484
rect 8216 11996 8280 12000
rect 8216 11940 8220 11996
rect 8220 11940 8276 11996
rect 8276 11940 8280 11996
rect 8216 11936 8280 11940
rect 8296 11996 8360 12000
rect 8296 11940 8300 11996
rect 8300 11940 8356 11996
rect 8356 11940 8360 11996
rect 8296 11936 8360 11940
rect 8376 11996 8440 12000
rect 8376 11940 8380 11996
rect 8380 11940 8436 11996
rect 8436 11940 8440 11996
rect 8376 11936 8440 11940
rect 8456 11996 8520 12000
rect 8456 11940 8460 11996
rect 8460 11940 8516 11996
rect 8516 11940 8520 11996
rect 8456 11936 8520 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 12216 11452 12280 11456
rect 12216 11396 12220 11452
rect 12220 11396 12276 11452
rect 12276 11396 12280 11452
rect 12216 11392 12280 11396
rect 12296 11452 12360 11456
rect 12296 11396 12300 11452
rect 12300 11396 12356 11452
rect 12356 11396 12360 11452
rect 12296 11392 12360 11396
rect 12376 11452 12440 11456
rect 12376 11396 12380 11452
rect 12380 11396 12436 11452
rect 12436 11396 12440 11452
rect 12376 11392 12440 11396
rect 12456 11452 12520 11456
rect 12456 11396 12460 11452
rect 12460 11396 12516 11452
rect 12516 11396 12520 11452
rect 12456 11392 12520 11396
rect 8216 10908 8280 10912
rect 8216 10852 8220 10908
rect 8220 10852 8276 10908
rect 8276 10852 8280 10908
rect 8216 10848 8280 10852
rect 8296 10908 8360 10912
rect 8296 10852 8300 10908
rect 8300 10852 8356 10908
rect 8356 10852 8360 10908
rect 8296 10848 8360 10852
rect 8376 10908 8440 10912
rect 8376 10852 8380 10908
rect 8380 10852 8436 10908
rect 8436 10852 8440 10908
rect 8376 10848 8440 10852
rect 8456 10908 8520 10912
rect 8456 10852 8460 10908
rect 8460 10852 8516 10908
rect 8516 10852 8520 10908
rect 8456 10848 8520 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 12216 10364 12280 10368
rect 12216 10308 12220 10364
rect 12220 10308 12276 10364
rect 12276 10308 12280 10364
rect 12216 10304 12280 10308
rect 12296 10364 12360 10368
rect 12296 10308 12300 10364
rect 12300 10308 12356 10364
rect 12356 10308 12360 10364
rect 12296 10304 12360 10308
rect 12376 10364 12440 10368
rect 12376 10308 12380 10364
rect 12380 10308 12436 10364
rect 12436 10308 12440 10364
rect 12376 10304 12440 10308
rect 12456 10364 12520 10368
rect 12456 10308 12460 10364
rect 12460 10308 12516 10364
rect 12516 10308 12520 10364
rect 12456 10304 12520 10308
rect 8216 9820 8280 9824
rect 8216 9764 8220 9820
rect 8220 9764 8276 9820
rect 8276 9764 8280 9820
rect 8216 9760 8280 9764
rect 8296 9820 8360 9824
rect 8296 9764 8300 9820
rect 8300 9764 8356 9820
rect 8356 9764 8360 9820
rect 8296 9760 8360 9764
rect 8376 9820 8440 9824
rect 8376 9764 8380 9820
rect 8380 9764 8436 9820
rect 8436 9764 8440 9820
rect 8376 9760 8440 9764
rect 8456 9820 8520 9824
rect 8456 9764 8460 9820
rect 8460 9764 8516 9820
rect 8516 9764 8520 9820
rect 8456 9760 8520 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 12216 9276 12280 9280
rect 12216 9220 12220 9276
rect 12220 9220 12276 9276
rect 12276 9220 12280 9276
rect 12216 9216 12280 9220
rect 12296 9276 12360 9280
rect 12296 9220 12300 9276
rect 12300 9220 12356 9276
rect 12356 9220 12360 9276
rect 12296 9216 12360 9220
rect 12376 9276 12440 9280
rect 12376 9220 12380 9276
rect 12380 9220 12436 9276
rect 12436 9220 12440 9276
rect 12376 9216 12440 9220
rect 12456 9276 12520 9280
rect 12456 9220 12460 9276
rect 12460 9220 12516 9276
rect 12516 9220 12520 9276
rect 12456 9216 12520 9220
rect 8216 8732 8280 8736
rect 8216 8676 8220 8732
rect 8220 8676 8276 8732
rect 8276 8676 8280 8732
rect 8216 8672 8280 8676
rect 8296 8732 8360 8736
rect 8296 8676 8300 8732
rect 8300 8676 8356 8732
rect 8356 8676 8360 8732
rect 8296 8672 8360 8676
rect 8376 8732 8440 8736
rect 8376 8676 8380 8732
rect 8380 8676 8436 8732
rect 8436 8676 8440 8732
rect 8376 8672 8440 8676
rect 8456 8732 8520 8736
rect 8456 8676 8460 8732
rect 8460 8676 8516 8732
rect 8516 8676 8520 8732
rect 8456 8672 8520 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 12216 8188 12280 8192
rect 12216 8132 12220 8188
rect 12220 8132 12276 8188
rect 12276 8132 12280 8188
rect 12216 8128 12280 8132
rect 12296 8188 12360 8192
rect 12296 8132 12300 8188
rect 12300 8132 12356 8188
rect 12356 8132 12360 8188
rect 12296 8128 12360 8132
rect 12376 8188 12440 8192
rect 12376 8132 12380 8188
rect 12380 8132 12436 8188
rect 12436 8132 12440 8188
rect 12376 8128 12440 8132
rect 12456 8188 12520 8192
rect 12456 8132 12460 8188
rect 12460 8132 12516 8188
rect 12516 8132 12520 8188
rect 12456 8128 12520 8132
rect 8216 7644 8280 7648
rect 8216 7588 8220 7644
rect 8220 7588 8276 7644
rect 8276 7588 8280 7644
rect 8216 7584 8280 7588
rect 8296 7644 8360 7648
rect 8296 7588 8300 7644
rect 8300 7588 8356 7644
rect 8356 7588 8360 7644
rect 8296 7584 8360 7588
rect 8376 7644 8440 7648
rect 8376 7588 8380 7644
rect 8380 7588 8436 7644
rect 8436 7588 8440 7644
rect 8376 7584 8440 7588
rect 8456 7644 8520 7648
rect 8456 7588 8460 7644
rect 8460 7588 8516 7644
rect 8516 7588 8520 7644
rect 8456 7584 8520 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 12216 7100 12280 7104
rect 12216 7044 12220 7100
rect 12220 7044 12276 7100
rect 12276 7044 12280 7100
rect 12216 7040 12280 7044
rect 12296 7100 12360 7104
rect 12296 7044 12300 7100
rect 12300 7044 12356 7100
rect 12356 7044 12360 7100
rect 12296 7040 12360 7044
rect 12376 7100 12440 7104
rect 12376 7044 12380 7100
rect 12380 7044 12436 7100
rect 12436 7044 12440 7100
rect 12376 7040 12440 7044
rect 12456 7100 12520 7104
rect 12456 7044 12460 7100
rect 12460 7044 12516 7100
rect 12516 7044 12520 7100
rect 12456 7040 12520 7044
rect 8216 6556 8280 6560
rect 8216 6500 8220 6556
rect 8220 6500 8276 6556
rect 8276 6500 8280 6556
rect 8216 6496 8280 6500
rect 8296 6556 8360 6560
rect 8296 6500 8300 6556
rect 8300 6500 8356 6556
rect 8356 6500 8360 6556
rect 8296 6496 8360 6500
rect 8376 6556 8440 6560
rect 8376 6500 8380 6556
rect 8380 6500 8436 6556
rect 8436 6500 8440 6556
rect 8376 6496 8440 6500
rect 8456 6556 8520 6560
rect 8456 6500 8460 6556
rect 8460 6500 8516 6556
rect 8516 6500 8520 6556
rect 8456 6496 8520 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 12216 6012 12280 6016
rect 12216 5956 12220 6012
rect 12220 5956 12276 6012
rect 12276 5956 12280 6012
rect 12216 5952 12280 5956
rect 12296 6012 12360 6016
rect 12296 5956 12300 6012
rect 12300 5956 12356 6012
rect 12356 5956 12360 6012
rect 12296 5952 12360 5956
rect 12376 6012 12440 6016
rect 12376 5956 12380 6012
rect 12380 5956 12436 6012
rect 12436 5956 12440 6012
rect 12376 5952 12440 5956
rect 12456 6012 12520 6016
rect 12456 5956 12460 6012
rect 12460 5956 12516 6012
rect 12516 5956 12520 6012
rect 12456 5952 12520 5956
rect 9260 5944 9324 5948
rect 9260 5888 9310 5944
rect 9310 5888 9324 5944
rect 9260 5884 9324 5888
rect 8216 5468 8280 5472
rect 8216 5412 8220 5468
rect 8220 5412 8276 5468
rect 8276 5412 8280 5468
rect 8216 5408 8280 5412
rect 8296 5468 8360 5472
rect 8296 5412 8300 5468
rect 8300 5412 8356 5468
rect 8356 5412 8360 5468
rect 8296 5408 8360 5412
rect 8376 5468 8440 5472
rect 8376 5412 8380 5468
rect 8380 5412 8436 5468
rect 8436 5412 8440 5468
rect 8376 5408 8440 5412
rect 8456 5468 8520 5472
rect 8456 5412 8460 5468
rect 8460 5412 8516 5468
rect 8516 5412 8520 5468
rect 8456 5408 8520 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 12216 4924 12280 4928
rect 12216 4868 12220 4924
rect 12220 4868 12276 4924
rect 12276 4868 12280 4924
rect 12216 4864 12280 4868
rect 12296 4924 12360 4928
rect 12296 4868 12300 4924
rect 12300 4868 12356 4924
rect 12356 4868 12360 4924
rect 12296 4864 12360 4868
rect 12376 4924 12440 4928
rect 12376 4868 12380 4924
rect 12380 4868 12436 4924
rect 12436 4868 12440 4924
rect 12376 4864 12440 4868
rect 12456 4924 12520 4928
rect 12456 4868 12460 4924
rect 12460 4868 12516 4924
rect 12516 4868 12520 4924
rect 12456 4864 12520 4868
rect 8216 4380 8280 4384
rect 8216 4324 8220 4380
rect 8220 4324 8276 4380
rect 8276 4324 8280 4380
rect 8216 4320 8280 4324
rect 8296 4380 8360 4384
rect 8296 4324 8300 4380
rect 8300 4324 8356 4380
rect 8356 4324 8360 4380
rect 8296 4320 8360 4324
rect 8376 4380 8440 4384
rect 8376 4324 8380 4380
rect 8380 4324 8436 4380
rect 8436 4324 8440 4380
rect 8376 4320 8440 4324
rect 8456 4380 8520 4384
rect 8456 4324 8460 4380
rect 8460 4324 8516 4380
rect 8516 4324 8520 4380
rect 8456 4320 8520 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 12216 3836 12280 3840
rect 12216 3780 12220 3836
rect 12220 3780 12276 3836
rect 12276 3780 12280 3836
rect 12216 3776 12280 3780
rect 12296 3836 12360 3840
rect 12296 3780 12300 3836
rect 12300 3780 12356 3836
rect 12356 3780 12360 3836
rect 12296 3776 12360 3780
rect 12376 3836 12440 3840
rect 12376 3780 12380 3836
rect 12380 3780 12436 3836
rect 12436 3780 12440 3836
rect 12376 3776 12440 3780
rect 12456 3836 12520 3840
rect 12456 3780 12460 3836
rect 12460 3780 12516 3836
rect 12516 3780 12520 3836
rect 12456 3776 12520 3780
rect 8216 3292 8280 3296
rect 8216 3236 8220 3292
rect 8220 3236 8276 3292
rect 8276 3236 8280 3292
rect 8216 3232 8280 3236
rect 8296 3292 8360 3296
rect 8296 3236 8300 3292
rect 8300 3236 8356 3292
rect 8356 3236 8360 3292
rect 8296 3232 8360 3236
rect 8376 3292 8440 3296
rect 8376 3236 8380 3292
rect 8380 3236 8436 3292
rect 8436 3236 8440 3292
rect 8376 3232 8440 3236
rect 8456 3292 8520 3296
rect 8456 3236 8460 3292
rect 8460 3236 8516 3292
rect 8516 3236 8520 3292
rect 8456 3232 8520 3236
rect 9260 3164 9324 3228
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 12216 2748 12280 2752
rect 12216 2692 12220 2748
rect 12220 2692 12276 2748
rect 12276 2692 12280 2748
rect 12216 2688 12280 2692
rect 12296 2748 12360 2752
rect 12296 2692 12300 2748
rect 12300 2692 12356 2748
rect 12356 2692 12360 2748
rect 12296 2688 12360 2692
rect 12376 2748 12440 2752
rect 12376 2692 12380 2748
rect 12380 2692 12436 2748
rect 12436 2692 12440 2748
rect 12376 2688 12440 2692
rect 12456 2748 12520 2752
rect 12456 2692 12460 2748
rect 12460 2692 12516 2748
rect 12516 2692 12520 2748
rect 12456 2688 12520 2692
rect 8216 2204 8280 2208
rect 8216 2148 8220 2204
rect 8220 2148 8276 2204
rect 8276 2148 8280 2204
rect 8216 2144 8280 2148
rect 8296 2204 8360 2208
rect 8296 2148 8300 2204
rect 8300 2148 8356 2204
rect 8356 2148 8360 2204
rect 8296 2144 8360 2148
rect 8376 2204 8440 2208
rect 8376 2148 8380 2204
rect 8380 2148 8436 2204
rect 8436 2148 8440 2204
rect 8376 2144 8440 2148
rect 8456 2204 8520 2208
rect 8456 2148 8460 2204
rect 8460 2148 8516 2204
rect 8516 2148 8520 2204
rect 8456 2144 8520 2148
rect 4216 1660 4280 1664
rect 4216 1604 4220 1660
rect 4220 1604 4276 1660
rect 4276 1604 4280 1660
rect 4216 1600 4280 1604
rect 4296 1660 4360 1664
rect 4296 1604 4300 1660
rect 4300 1604 4356 1660
rect 4356 1604 4360 1660
rect 4296 1600 4360 1604
rect 4376 1660 4440 1664
rect 4376 1604 4380 1660
rect 4380 1604 4436 1660
rect 4436 1604 4440 1660
rect 4376 1600 4440 1604
rect 4456 1660 4520 1664
rect 4456 1604 4460 1660
rect 4460 1604 4516 1660
rect 4516 1604 4520 1660
rect 4456 1600 4520 1604
rect 12216 1660 12280 1664
rect 12216 1604 12220 1660
rect 12220 1604 12276 1660
rect 12276 1604 12280 1660
rect 12216 1600 12280 1604
rect 12296 1660 12360 1664
rect 12296 1604 12300 1660
rect 12300 1604 12356 1660
rect 12356 1604 12360 1660
rect 12296 1600 12360 1604
rect 12376 1660 12440 1664
rect 12376 1604 12380 1660
rect 12380 1604 12436 1660
rect 12436 1604 12440 1660
rect 12376 1600 12440 1604
rect 12456 1660 12520 1664
rect 12456 1604 12460 1660
rect 12460 1604 12516 1660
rect 12516 1604 12520 1660
rect 12456 1600 12520 1604
rect 8216 1116 8280 1120
rect 8216 1060 8220 1116
rect 8220 1060 8276 1116
rect 8276 1060 8280 1116
rect 8216 1056 8280 1060
rect 8296 1116 8360 1120
rect 8296 1060 8300 1116
rect 8300 1060 8356 1116
rect 8356 1060 8360 1116
rect 8296 1056 8360 1060
rect 8376 1116 8440 1120
rect 8376 1060 8380 1116
rect 8380 1060 8436 1116
rect 8436 1060 8440 1116
rect 8376 1056 8440 1060
rect 8456 1116 8520 1120
rect 8456 1060 8460 1116
rect 8460 1060 8516 1116
rect 8516 1060 8520 1116
rect 8456 1056 8520 1060
<< metal4 >>
rect 4208 13632 4528 13648
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12488 4296 12544
rect 4360 12488 4376 12544
rect 4440 12488 4456 12544
rect 4520 12480 4528 12544
rect 4208 12252 4250 12480
rect 4486 12252 4528 12480
rect 4208 11456 4528 12252
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4488 4528 4864
rect 4208 4252 4250 4488
rect 4486 4252 4528 4488
rect 4208 3840 4528 4252
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 1664 4528 2688
rect 4208 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4528 1664
rect 4208 1040 4528 1600
rect 8208 13088 8528 13648
rect 8208 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8528 13088
rect 8208 12000 8528 13024
rect 8208 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8528 12000
rect 8208 10912 8528 11936
rect 8208 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8528 10912
rect 8208 9824 8528 10848
rect 8208 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8528 9824
rect 8208 8736 8528 9760
rect 8208 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8528 8736
rect 8208 8488 8528 8672
rect 8208 8252 8250 8488
rect 8486 8252 8528 8488
rect 8208 7648 8528 8252
rect 8208 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8528 7648
rect 8208 6560 8528 7584
rect 8208 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8528 6560
rect 8208 5472 8528 6496
rect 12208 13632 12528 13648
rect 12208 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12528 13632
rect 12208 12544 12528 13568
rect 12208 12480 12216 12544
rect 12280 12488 12296 12544
rect 12360 12488 12376 12544
rect 12440 12488 12456 12544
rect 12520 12480 12528 12544
rect 12208 12252 12250 12480
rect 12486 12252 12528 12480
rect 12208 11456 12528 12252
rect 12208 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12528 11456
rect 12208 10368 12528 11392
rect 12208 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12528 10368
rect 12208 9280 12528 10304
rect 12208 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12528 9280
rect 12208 8192 12528 9216
rect 12208 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12528 8192
rect 12208 7104 12528 8128
rect 12208 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12528 7104
rect 12208 6016 12528 7040
rect 12208 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12528 6016
rect 9259 5948 9325 5949
rect 9259 5884 9260 5948
rect 9324 5884 9325 5948
rect 9259 5883 9325 5884
rect 8208 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8528 5472
rect 8208 4384 8528 5408
rect 8208 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8528 4384
rect 8208 3296 8528 4320
rect 8208 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8528 3296
rect 8208 2208 8528 3232
rect 9262 3229 9322 5883
rect 12208 4928 12528 5952
rect 12208 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12528 4928
rect 12208 4488 12528 4864
rect 12208 4252 12250 4488
rect 12486 4252 12528 4488
rect 12208 3840 12528 4252
rect 12208 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12528 3840
rect 9259 3228 9325 3229
rect 9259 3164 9260 3228
rect 9324 3164 9325 3228
rect 9259 3163 9325 3164
rect 8208 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8528 2208
rect 8208 1120 8528 2144
rect 8208 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8528 1120
rect 8208 1040 8528 1056
rect 12208 2752 12528 3776
rect 12208 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12528 2752
rect 12208 1664 12528 2688
rect 12208 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12528 1664
rect 12208 1040 12528 1600
<< via4 >>
rect 4250 12480 4280 12488
rect 4280 12480 4296 12488
rect 4296 12480 4360 12488
rect 4360 12480 4376 12488
rect 4376 12480 4440 12488
rect 4440 12480 4456 12488
rect 4456 12480 4486 12488
rect 4250 12252 4486 12480
rect 4250 4252 4486 4488
rect 8250 8252 8486 8488
rect 12250 12480 12280 12488
rect 12280 12480 12296 12488
rect 12296 12480 12360 12488
rect 12360 12480 12376 12488
rect 12376 12480 12440 12488
rect 12440 12480 12456 12488
rect 12456 12480 12486 12488
rect 12250 12252 12486 12480
rect 12250 4252 12486 4488
<< metal5 >>
rect 1104 12488 13892 12530
rect 1104 12252 4250 12488
rect 4486 12252 12250 12488
rect 12486 12252 13892 12488
rect 1104 12210 13892 12252
rect 1104 8488 13892 8530
rect 1104 8252 8250 8488
rect 8486 8252 13892 8488
rect 1104 8210 13892 8252
rect 1104 4488 13892 4530
rect 1104 4252 4250 4488
rect 4486 4252 12250 4488
rect 12486 4252 13892 4488
rect 1104 4210 13892 4252
use sky130_fd_sc_hd__decap_8  FILLER_0_13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2300 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3036 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1380 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1932 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1636915332
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2024 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _356_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1380 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__D $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 3680 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _324_
timestamp 1636915332
transform 1 0 3220 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _357_
timestamp 1636915332
transform -1 0 5244 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _367_
timestamp 1636915332
transform -1 0 5704 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__o2bb2a_2  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5244 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 6256 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50
timestamp 1636915332
transform 1 0 5704 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1636915332
transform -1 0 6256 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 7268 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 6440 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1636915332
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1636915332
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 1636915332
transform 1 0 6348 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 7544 0 1 1088
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75
timestamp 1636915332
transform 1 0 8004 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1636915332
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1636915332
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _354_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8924 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8924 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8004 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8096 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.iss.delayenb0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7268 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen1
timestamp 1636915332
transform 1 0 9752 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_1_88
timestamp 1636915332
transform 1 0 9200 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10304 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _330_
timestamp 1636915332
transform -1 0 11408 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1636915332
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A1
timestamp 1636915332
transform 1 0 10948 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__S
timestamp 1636915332
transform 1 0 10764 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A1
timestamp 1636915332
transform 1 0 10580 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__S
timestamp 1636915332
transform 1 0 10396 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9292 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1636915332
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1636915332
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_118
timestamp 1636915332
transform 1 0 11960 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp 1636915332
transform 1 0 11500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__S
timestamp 1636915332
transform 1 0 12144 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__S
timestamp 1636915332
transform 1 0 11776 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__A1
timestamp 1636915332
transform 1 0 11592 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 13156 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb1
timestamp 1636915332
transform 1 0 12328 0 1 1088
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp 1636915332
transform 1 0 11500 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_1_135
timestamp 1636915332
transform 1 0 13524 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1636915332
transform -1 0 13892 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1636915332
transform -1 0 13892 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1636915332
transform 1 0 13340 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1636915332
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1636915332
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _358_
timestamp 1636915332
transform 1 0 1564 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1636915332
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_39
timestamp 1636915332
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1636915332
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _313_
timestamp 1636915332
transform 1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _314_
timestamp 1636915332
transform 1 0 4140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _370_
timestamp 1636915332
transform 1 0 4876 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__B
timestamp 1636915332
transform -1 0 6992 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen1
timestamp 1636915332
transform 1 0 6992 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A1
timestamp 1636915332
transform -1 0 9200 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__S
timestamp 1636915332
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_80
timestamp 1636915332
transform 1 0 8464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1636915332
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1636915332
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0
timestamp 1636915332
transform -1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.reseten0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7636 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__S
timestamp 1636915332
transform 1 0 10948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_106
timestamp 1636915332
transform 1 0 10856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_88
timestamp 1636915332
transform 1 0 9200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _278_
timestamp 1636915332
transform -1 0 10856 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1636915332
transform 1 0 9568 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen0
timestamp 1636915332
transform 1 0 11132 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 9568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_116
timestamp 1636915332
transform 1 0 11776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _331_
timestamp 1636915332
transform -1 0 12696 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen1
timestamp 1636915332
transform 1 0 12696 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1636915332
transform -1 0 13892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1636915332
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1636915332
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_2  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2760 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _323_
timestamp 1636915332
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _368_
timestamp 1636915332
transform 1 0 3588 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A
timestamp 1636915332
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_48
timestamp 1636915332
transform 1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1636915332
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_59
timestamp 1636915332
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1636915332
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _311_
timestamp 1636915332
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[0\].id.delayenb1
timestamp 1636915332
transform 1 0 6808 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A1
timestamp 1636915332
transform 1 0 8832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_73
timestamp 1636915332
transform 1 0 7820 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _288_
timestamp 1636915332
transform -1 0 9476 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1636915332
transform 1 0 8004 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_2  _282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10304 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _326_
timestamp 1636915332
transform 1 0 11040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _339_
timestamp 1636915332
transform -1 0 10304 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A1
timestamp 1636915332
transform -1 0 12512 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1636915332
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1636915332
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _332_
timestamp 1636915332
transform 1 0 12512 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _333_
timestamp 1636915332
transform 1 0 11500 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1636915332
transform -1 0 13892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1636915332
transform 1 0 13340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1636915332
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_19
timestamp 1636915332
transform 1 0 2852 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1636915332
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_8
timestamp 1636915332
transform 1 0 1840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1636915332
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _315_
timestamp 1636915332
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _328_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 1840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1636915332
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_41
timestamp 1636915332
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1636915332
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4968 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _258_
timestamp 1636915332
transform -1 0 3680 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_4_49
timestamp 1636915332
transform 1 0 5612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_59
timestamp 1636915332
transform 1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_63
timestamp 1636915332
transform 1 0 6900 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5796 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0
timestamp 1636915332
transform 1 0 6992 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__S
timestamp 1636915332
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_87
timestamp 1636915332
transform 1 0 9108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1636915332
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_2  _291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8188 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1636915332
transform 1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 1636915332
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_106
timestamp 1636915332
transform 1 0 10856 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o41a_2  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 10120 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_2  _303_
timestamp 1636915332
transform 1 0 10120 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[10\].id.delayenb1
timestamp 1636915332
transform 1 0 10948 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[10\].id.delayenb0
timestamp 1636915332
transform 1 0 11960 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1636915332
transform -1 0 13892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1636915332
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _366_
timestamp 1636915332
transform 1 0 1380 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_5_41
timestamp 1636915332
transform 1 0 4876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _240_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 4876 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _263_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 4140 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1636915332
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1636915332
transform -1 0 6256 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1636915332
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5152 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[0\].id.delayenb0
timestamp 1636915332
transform 1 0 6624 0 -1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A1
timestamp 1636915332
transform 1 0 8740 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__S
timestamp 1636915332
transform 1 0 9016 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1636915332
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_82
timestamp 1636915332
transform 1 0 8648 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_85
timestamp 1636915332
transform 1 0 8924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _229_
timestamp 1636915332
transform 1 0 9200 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1636915332
transform -1 0 11316 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10488 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_2  _304_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9660 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A1
timestamp 1636915332
transform -1 0 12420 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1636915332
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1636915332
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1636915332
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1636915332
transform 1 0 13064 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp 1636915332
transform 1 0 12420 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen1
timestamp 1636915332
transform 1 0 11592 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__A1
timestamp 1636915332
transform -1 0 13616 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_133
timestamp 1636915332
transform 1 0 13340 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1636915332
transform -1 0 13892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_13
timestamp 1636915332
transform 1 0 2300 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1636915332
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_9
timestamp 1636915332
transform 1 0 1932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1636915332
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1636915332
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _266_
timestamp 1636915332
transform 1 0 2392 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _317_
timestamp 1636915332
transform 1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _364_
timestamp 1636915332
transform 1 0 1380 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_2  _262_
timestamp 1636915332
transform -1 0 3680 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _259_
timestamp 1636915332
transform -1 0 4600 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_2  _238_
timestamp 1636915332
transform 1 0 3496 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1636915332
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_24
timestamp 1636915332
transform 1 0 3312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_22
timestamp 1636915332
transform 1 0 3128 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_2  _260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4232 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _257_
timestamp 1636915332
transform 1 0 4784 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_38
timestamp 1636915332
transform 1 0 4600 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_42
timestamp 1636915332
transform 1 0 4968 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_2  _256_
timestamp 1636915332
transform 1 0 5152 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _251_
timestamp 1636915332
transform -1 0 6072 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_6_53
timestamp 1636915332
transform 1 0 5980 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_49
timestamp 1636915332
transform 1 0 5612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_2  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 6348 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_2  _241_
timestamp 1636915332
transform 1 0 6072 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1636915332
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1636915332
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_63
timestamp 1636915332
transform 1 0 6900 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _239_
timestamp 1636915332
transform -1 0 7452 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _221_
timestamp 1636915332
transform 1 0 7268 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1636915332
transform 1 0 7728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1636915332
transform 1 0 7728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _170_
timestamp 1636915332
transform 1 0 7452 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_75
timestamp 1636915332
transform 1 0 8004 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_66
timestamp 1636915332
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_75
timestamp 1636915332
transform 1 0 8004 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _335_
timestamp 1636915332
transform -1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_2  _300_
timestamp 1636915332
transform -1 0 9108 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o41a_2  _296_
timestamp 1636915332
transform 1 0 9108 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__or2_2  _227_
timestamp 1636915332
transform 1 0 8372 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1636915332
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_107
timestamp 1636915332
transform 1 0 10948 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_97
timestamp 1636915332
transform 1 0 10028 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1636915332
transform -1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_2  _293_
timestamp 1636915332
transform -1 0 10948 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _294_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 11408 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_2  _295_
timestamp 1636915332
transform 1 0 10028 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen1
timestamp 1636915332
transform 1 0 11040 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1636915332
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _231_
timestamp 1636915332
transform 1 0 11500 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1636915332
transform -1 0 13340 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1636915332
transform 1 0 12696 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[9\].id.delayenb0
timestamp 1636915332
transform 1 0 11960 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[9\].id.delayenb1
timestamp 1636915332
transform 1 0 11684 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__S
timestamp 1636915332
transform 1 0 13340 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_135
timestamp 1636915332
transform 1 0 13524 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1636915332
transform -1 0 13892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1636915332
transform -1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_13
timestamp 1636915332
transform 1 0 2300 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_21
timestamp 1636915332
transform 1 0 3036 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1636915332
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1636915332
transform 1 0 1932 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1636915332
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _316_
timestamp 1636915332
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1636915332
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1636915332
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1636915332
transform 1 0 3128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1636915332
transform -1 0 3680 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _233_
timestamp 1636915332
transform 1 0 3864 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_2  _235_
timestamp 1636915332
transform 1 0 4416 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_44
timestamp 1636915332
transform 1 0 5152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_63
timestamp 1636915332
transform 1 0 6900 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1636915332
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _242_
timestamp 1636915332
transform -1 0 5980 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _252_
timestamp 1636915332
transform -1 0 6624 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1636915332
transform 1 0 6624 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1636915332
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1636915332
transform 1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _223_
timestamp 1636915332
transform -1 0 7912 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _297_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8188 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_2  _298_
timestamp 1636915332
transform -1 0 9752 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_103
timestamp 1636915332
transform 1 0 10580 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _337_
timestamp 1636915332
transform 1 0 10672 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _349_
timestamp 1636915332
transform -1 0 10580 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__S
timestamp 1636915332
transform 1 0 12328 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _347_
timestamp 1636915332
transform -1 0 12328 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 1636915332
transform 1 0 12512 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1636915332
transform 1 0 13156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A1
timestamp 1636915332
transform -1 0 13616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1636915332
transform -1 0 13892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1636915332
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _365_
timestamp 1636915332
transform 1 0 1380 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1636915332
transform 1 0 5060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_2  _264_
timestamp 1636915332
transform -1 0 5060 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o22ai_2  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3312 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1636915332
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1636915332
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _232_
timestamp 1636915332
transform -1 0 7544 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_2  _243_
timestamp 1636915332
transform -1 0 7084 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _254_
timestamp 1636915332
transform 1 0 5336 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__A1
timestamp 1636915332
transform -1 0 7728 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_72
timestamp 1636915332
transform 1 0 7728 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_82
timestamp 1636915332
transform 1 0 8648 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o31a_2  _283_
timestamp 1636915332
transform 1 0 8740 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1636915332
transform 1 0 7820 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A1
timestamp 1636915332
transform -1 0 10396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A1
timestamp 1636915332
transform -1 0 10212 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__S
timestamp 1636915332
transform 1 0 9844 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A1
timestamp 1636915332
transform 1 0 9476 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__S
timestamp 1636915332
transform 1 0 9660 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_2  _292_
timestamp 1636915332
transform 1 0 10396 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 11408 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_122
timestamp 1636915332
transform 1 0 12328 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1636915332
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _329_
timestamp 1636915332
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _343_
timestamp 1636915332
transform 1 0 12788 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1636915332
transform 1 0 12420 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1636915332
transform -1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1636915332
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1636915332
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1636915332
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _189_
timestamp 1636915332
transform -1 0 2852 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _310_
timestamp 1636915332
transform 1 0 2116 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1636915332
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_43
timestamp 1636915332
transform 1 0 5060 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1636915332
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _224_
timestamp 1636915332
transform -1 0 5060 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _237_
timestamp 1636915332
transform -1 0 4508 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1636915332
transform -1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _369_
timestamp 1636915332
transform 1 0 5428 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__S
timestamp 1636915332
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1636915332
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _280_
timestamp 1636915332
transform 1 0 8188 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1636915332
transform 1 0 7360 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1636915332
transform -1 0 9292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_2  _285_
timestamp 1636915332
transform -1 0 10212 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _345_
timestamp 1636915332
transform -1 0 11040 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen1
timestamp 1636915332
transform 1 0 11040 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__A1
timestamp 1636915332
transform -1 0 12512 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__S
timestamp 1636915332
transform 1 0 12144 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_2  _301_
timestamp 1636915332
transform 1 0 11684 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _334_
timestamp 1636915332
transform 1 0 12512 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__A1
timestamp 1636915332
transform 1 0 13432 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_133
timestamp 1636915332
transform 1 0 13340 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1636915332
transform -1 0 13892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1636915332
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _371_
timestamp 1636915332
transform 1 0 1380 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_11_32
timestamp 1636915332
transform 1 0 4048 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _188_
timestamp 1636915332
transform -1 0 4048 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4416 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_45
timestamp 1636915332
transform 1 0 5244 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1636915332
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1636915332
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1636915332
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1636915332
transform -1 0 6808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _255_
timestamp 1636915332
transform 1 0 5428 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen1
timestamp 1636915332
transform 1 0 6808 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _289_
timestamp 1636915332
transform 1 0 8464 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[1\].id.delayenb1
timestamp 1636915332
transform 1 0 7452 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__S
timestamp 1636915332
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_106
timestamp 1636915332
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_88
timestamp 1636915332
transform 1 0 9200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_96
timestamp 1636915332
transform 1 0 9936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__o31a_2  _281_
timestamp 1636915332
transform -1 0 10856 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9292 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__A1
timestamp 1636915332
transform -1 0 13156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__S
timestamp 1636915332
transform 1 0 12788 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__S
timestamp 1636915332
transform 1 0 13156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A1
timestamp 1636915332
transform -1 0 11408 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1636915332
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_117
timestamp 1636915332
transform 1 0 11868 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1636915332
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _336_
timestamp 1636915332
transform 1 0 11960 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1636915332
transform 1 0 11592 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__S
timestamp 1636915332
transform 1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_135
timestamp 1636915332
transform 1 0 13524 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1636915332
transform -1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1636915332
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _372_
timestamp 1636915332
transform 1 0 1380 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1636915332
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1636915332
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _373_
timestamp 1636915332
transform 1 0 3772 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_12_53
timestamp 1636915332
transform 1 0 5980 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1636915332
transform -1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _219_
timestamp 1636915332
transform 1 0 6532 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _312_
timestamp 1636915332
transform -1 0 7268 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_67
timestamp 1636915332
transform 1 0 7268 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1636915332
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1636915332
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1636915332
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o41a_2  _286_
timestamp 1636915332
transform 1 0 9016 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1636915332
transform 1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp 1636915332
transform 1 0 7820 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1636915332
transform 1 0 7544 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_103
timestamp 1636915332
transform 1 0 10580 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__a31o_2  _290_
timestamp 1636915332
transform -1 0 10580 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[8\].id.delayenb1
timestamp 1636915332
transform 1 0 10764 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[8\].id.delayenb0
timestamp 1636915332
transform 1 0 11776 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A1
timestamp 1636915332
transform -1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1636915332
transform -1 0 13892 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_16
timestamp 1636915332
transform 1 0 2576 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1636915332
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1636915332
transform 1 0 1932 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1636915332
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1636915332
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _309_
timestamp 1636915332
transform 1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _318_
timestamp 1636915332
transform 1 0 2300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _363_
timestamp 1636915332
transform 1 0 1380 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__a21oi_2  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 4416 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3864 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _187_
timestamp 1636915332
transform 1 0 3128 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1636915332
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1636915332
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _319_
timestamp 1636915332
transform 1 0 4692 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _308_
timestamp 1636915332
transform 1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _180_
timestamp 1636915332
transform 1 0 4876 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1636915332
transform 1 0 4416 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _378_
timestamp 1636915332
transform 1 0 4968 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_13_49
timestamp 1636915332
transform 1 0 5612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1636915332
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1636915332
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1636915332
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1636915332
transform 1 0 6900 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _327_
timestamp 1636915332
transform 1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1636915332
transform 1 0 7544 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A1
timestamp 1636915332
transform 1 0 7176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__B1
timestamp 1636915332
transform -1 0 7544 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1636915332
transform 1 0 9108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1636915332
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1636915332
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1636915332
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__S
timestamp 1636915332
transform 1 0 8556 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__S
timestamp 1636915332
transform 1 0 9108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A1
timestamp 1636915332
transform -1 0 8556 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[1\].id.delayenb0
timestamp 1636915332
transform 1 0 7452 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_14_100
timestamp 1636915332
transform 1 0 10304 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_89
timestamp 1636915332
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _338_
timestamp 1636915332
transform -1 0 11592 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1636915332
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp 1636915332
transform 1 0 9660 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen1
timestamp 1636915332
transform 1 0 10488 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[2\].id.delayenb1
timestamp 1636915332
transform -1 0 10488 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1636915332
transform -1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1636915332
transform 1 0 10396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1636915332
transform 1 0 11684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1636915332
transform 1 0 11960 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1636915332
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_118
timestamp 1636915332
transform 1 0 11960 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1636915332
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__S
timestamp 1636915332
transform 1 0 11592 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__A1
timestamp 1636915332
transform -1 0 11960 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1636915332
transform -1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1636915332
transform 1 0 12788 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__S
timestamp 1636915332
transform 1 0 12604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[7\].id.delayenb1
timestamp 1636915332
transform 1 0 12144 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_14_135
timestamp 1636915332
transform 1 0 13524 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1636915332
transform -1 0 13892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1636915332
transform -1 0 13892 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_14
timestamp 1636915332
transform 1 0 2392 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1636915332
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1636915332
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _271_
timestamp 1636915332
transform 1 0 2944 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _307_
timestamp 1636915332
transform -1 0 2392 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _362_
timestamp 1636915332
transform 1 0 3772 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_15_50
timestamp 1636915332
transform 1 0 5704 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1636915332
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _214_
timestamp 1636915332
transform -1 0 6256 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o221ai_2  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_77
timestamp 1636915332
transform 1 0 8188 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _212_
timestamp 1636915332
transform 1 0 7452 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _348_
timestamp 1636915332
transform -1 0 9108 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[2\].id.delayenb0
timestamp 1636915332
transform 1 0 9108 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen1
timestamp 1636915332
transform 1 0 10764 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1636915332
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1636915332
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[7\].id.delayenb0
timestamp 1636915332
transform 1 0 11592 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_15_135
timestamp 1636915332
transform 1 0 13524 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1636915332
transform -1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1636915332
transform 1 0 13248 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1636915332
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _374_
timestamp 1636915332
transform -1 0 3312 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1636915332
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_41
timestamp 1636915332
transform 1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1636915332
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _208_
timestamp 1636915332
transform 1 0 4232 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _269_
timestamp 1636915332
transform -1 0 4232 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _377_
timestamp 1636915332
transform 1 0 5152 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A
timestamp 1636915332
transform 1 0 7820 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A1
timestamp 1636915332
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1636915332
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _211_
timestamp 1636915332
transform 1 0 8004 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _216_
timestamp 1636915332
transform 1 0 8924 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A
timestamp 1636915332
transform 1 0 9660 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1636915332
transform 1 0 9844 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__S
timestamp 1636915332
transform 1 0 10028 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_99
timestamp 1636915332
transform 1 0 10212 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1636915332
transform -1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[3\].id.delayenb1
timestamp 1636915332
transform -1 0 11776 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen1
timestamp 1636915332
transform -1 0 12420 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1636915332
transform -1 0 13340 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1636915332
transform 1 0 12420 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1636915332
transform -1 0 13892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1636915332
transform 1 0 13340 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_13
timestamp 1636915332
transform 1 0 2300 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1636915332
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1636915332
transform 1 0 1932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1636915332
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _186_
timestamp 1636915332
transform 1 0 2392 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _322_
timestamp 1636915332
transform 1 0 2024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_39
timestamp 1636915332
transform 1 0 4692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__o2bb2ai_2  _206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_2  _272_
timestamp 1636915332
transform -1 0 4692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_2  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3128 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1636915332
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1636915332
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1636915332
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _190_
timestamp 1636915332
transform 1 0 6716 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _209_
timestamp 1636915332
transform 1 0 6440 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_66
timestamp 1636915332
transform 1 0 7176 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_2  _207_
timestamp 1636915332
transform 1 0 7360 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _210_
timestamp 1636915332
transform -1 0 9752 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o2111ai_2  _225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A1
timestamp 1636915332
transform 1 0 10212 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__B1
timestamp 1636915332
transform 1 0 10396 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _279_
timestamp 1636915332
transform 1 0 9752 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp 1636915332
transform 1 0 10580 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1636915332
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_119
timestamp 1636915332
transform 1 0 12052 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1636915332
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1636915332
transform -1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1636915332
transform 1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen1
timestamp 1636915332
transform 1 0 12696 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1636915332
transform 1 0 12328 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1636915332
transform -1 0 13892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1636915332
transform 1 0 13340 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1636915332
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _359_
timestamp 1636915332
transform -1 0 3312 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1636915332
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1636915332
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1636915332
transform 1 0 3312 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1636915332
transform 1 0 4692 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _183_
timestamp 1636915332
transform 1 0 4968 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _193_
timestamp 1636915332
transform 1 0 4232 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _276_
timestamp 1636915332
transform 1 0 3772 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _195_
timestamp 1636915332
transform 1 0 5704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_2  _213_
timestamp 1636915332
transform 1 0 6440 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1636915332
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1636915332
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1636915332
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_2  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 7912 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_2  _217_
timestamp 1636915332
transform -1 0 8740 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _346_
timestamp 1636915332
transform -1 0 9844 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[3\].id.delayenb0
timestamp 1636915332
transform 1 0 9844 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__A1
timestamp 1636915332
transform -1 0 11684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__S
timestamp 1636915332
transform 1 0 11684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp 1636915332
transform 1 0 11868 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[6\].id.delayenb1
timestamp 1636915332
transform 1 0 12512 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_18_135
timestamp 1636915332
transform 1 0 13524 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1636915332
transform -1 0 13892 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_11
timestamp 1636915332
transform 1 0 2116 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1636915332
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_16
timestamp 1636915332
transform 1 0 2576 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1636915332
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1636915332
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1636915332
transform -1 0 2668 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _273_
timestamp 1636915332
transform 1 0 2668 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_2  _275_
timestamp 1636915332
transform 1 0 2760 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp11
timestamp 1636915332
transform -1 0 2576 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_19_31
timestamp 1636915332
transform 1 0 3956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1636915332
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_32
timestamp 1636915332
transform 1 0 4048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1636915332
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1636915332
transform -1 0 4048 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _185_
timestamp 1636915332
transform -1 0 4876 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1636915332
transform 1 0 4876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _274_
timestamp 1636915332
transform 1 0 3312 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_2  _375_
timestamp 1636915332
transform 1 0 4140 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__o2bb2a_2  _194_
timestamp 1636915332
transform 1 0 5152 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1636915332
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _306_
timestamp 1636915332
transform -1 0 6348 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _305_
timestamp 1636915332
transform 1 0 6440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_2  _198_
timestamp 1636915332
transform 1 0 6624 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1636915332
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_61
timestamp 1636915332
transform 1 0 6716 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_57
timestamp 1636915332
transform 1 0 6348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 1636915332
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _197_
timestamp 1636915332
transform 1 0 6992 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _205_
timestamp 1636915332
transform -1 0 8004 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1636915332
transform -1 0 8280 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_2  _200_
timestamp 1636915332
transform -1 0 8648 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_69
timestamp 1636915332
transform 1 0 7452 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__A1
timestamp 1636915332
transform 1 0 7544 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__o211a_2  _204_
timestamp 1636915332
transform -1 0 9016 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _202_
timestamp 1636915332
transform -1 0 9476 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_2  _201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8924 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1636915332
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__A1
timestamp 1636915332
transform -1 0 8832 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__A1
timestamp 1636915332
transform -1 0 10580 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_91
timestamp 1636915332
transform 1 0 9476 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _340_
timestamp 1636915332
transform -1 0 10396 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1636915332
transform -1 0 11224 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1636915332
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen1
timestamp 1636915332
transform -1 0 11500 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[4\].id.delayenb1
timestamp 1636915332
transform 1 0 9844 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__B1
timestamp 1636915332
transform -1 0 11684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A
timestamp 1636915332
transform -1 0 11408 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_122
timestamp 1636915332
transform 1 0 12328 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1636915332
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1636915332
transform 1 0 11684 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb1
timestamp 1636915332
transform 1 0 12512 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1636915332
transform 1 0 13156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[6\].id.delayenb0
timestamp 1636915332
transform 1 0 11500 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_19_135
timestamp 1636915332
transform 1 0 13524 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_135
timestamp 1636915332
transform 1 0 13524 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1636915332
transform -1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1636915332
transform -1 0 13892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1636915332
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1636915332
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _361_
timestamp 1636915332
transform 1 0 1564 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_21_26
timestamp 1636915332
transform 1 0 3496 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _360_
timestamp 1636915332
transform 1 0 3588 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1636915332
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _184_
timestamp 1636915332
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _376_
timestamp 1636915332
transform 1 0 6348 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_21_78
timestamp 1636915332
transform 1 0 8280 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _342_
timestamp 1636915332
transform -1 0 9200 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__S
timestamp 1636915332
transform 1 0 9200 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__A1
timestamp 1636915332
transform -1 0 9568 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[4\].id.delayenb0
timestamp 1636915332
transform 1 0 9568 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1636915332
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1636915332
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1636915332
transform -1 0 13432 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[5\].id.delayenb0
timestamp 1636915332
transform 1 0 11500 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_21_134
timestamp 1636915332
transform 1 0 13432 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1636915332
transform -1 0 13892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_11
timestamp 1636915332
transform 1 0 2116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_17
timestamp 1636915332
transform 1 0 2668 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1636915332
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1636915332
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _267_
timestamp 1636915332
transform 1 0 2944 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _320_
timestamp 1636915332
transform 1 0 2392 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1636915332
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_29
timestamp 1636915332
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_35
timestamp 1636915332
transform 1 0 4324 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_39
timestamp 1636915332
transform 1 0 4692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1636915332
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _321_
timestamp 1636915332
transform 1 0 4416 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_51
timestamp 1636915332
transform 1 0 5796 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_55
timestamp 1636915332
transform 1 0 6164 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_57
timestamp 1636915332
transform 1 0 6348 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_65
timestamp 1636915332
transform 1 0 7084 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1636915332
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A1
timestamp 1636915332
transform 1 0 8556 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1636915332
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1636915332
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _192_
timestamp 1636915332
transform 1 0 7820 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1636915332
transform 1 0 8280 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _199_
timestamp 1636915332
transform 1 0 7176 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _344_
timestamp 1636915332
transform -1 0 9752 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__S
timestamp 1636915332
transform 1 0 10764 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_107
timestamp 1636915332
transform 1 0 10948 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_94
timestamp 1636915332
transform 1 0 9752 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1636915332
transform 1 0 9844 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1636915332
transform -1 0 10764 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_111
timestamp 1636915332
transform 1 0 11316 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_121
timestamp 1636915332
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_125
timestamp 1636915332
transform 1 0 12604 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1636915332
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1636915332
transform 1 0 11500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen1
timestamp 1636915332
transform 1 0 12696 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp10
timestamp 1636915332
transform -1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1636915332
transform -1 0 13892 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1636915332
transform 1 0 13340 0 1 13056
box -38 -48 314 592
<< labels >>
rlabel metal5 s 1104 8210 13892 8530 6 VGND
port 0 nsew ground input
rlabel metal4 s 8208 1040 8528 13648 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 4210 13892 4530 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 12210 13892 12530 6 VPWR
port 1 nsew power input
rlabel metal4 s 4208 1040 4528 13648 6 VPWR
port 1 nsew power input
rlabel metal4 s 12208 1040 12528 13648 6 VPWR
port 1 nsew power input
rlabel metal3 s 0 3680 800 3800 6 clockp[0]
port 2 nsew signal tristate
rlabel metal3 s 0 11160 800 11280 6 clockp[1]
port 3 nsew signal tristate
rlabel metal3 s 14200 14424 15000 14544 6 dco
port 4 nsew signal input
rlabel metal3 s 14200 10072 15000 10192 6 div[0]
port 5 nsew signal input
rlabel metal3 s 14200 10888 15000 11008 6 div[1]
port 6 nsew signal input
rlabel metal3 s 14200 11840 15000 11960 6 div[2]
port 7 nsew signal input
rlabel metal3 s 14200 12656 15000 12776 6 div[3]
port 8 nsew signal input
rlabel metal3 s 14200 13608 15000 13728 6 div[4]
port 9 nsew signal input
rlabel metal3 s 14200 9120 15000 9240 6 enable
port 10 nsew signal input
rlabel metal2 s 754 14200 810 15000 6 ext_trim[0]
port 11 nsew signal input
rlabel metal3 s 14200 416 15000 536 6 ext_trim[10]
port 12 nsew signal input
rlabel metal3 s 14200 1232 15000 1352 6 ext_trim[11]
port 13 nsew signal input
rlabel metal3 s 14200 2048 15000 2168 6 ext_trim[12]
port 14 nsew signal input
rlabel metal3 s 14200 3000 15000 3120 6 ext_trim[13]
port 15 nsew signal input
rlabel metal3 s 14200 3816 15000 3936 6 ext_trim[14]
port 16 nsew signal input
rlabel metal3 s 14200 4768 15000 4888 6 ext_trim[15]
port 17 nsew signal input
rlabel metal3 s 14200 5584 15000 5704 6 ext_trim[16]
port 18 nsew signal input
rlabel metal3 s 14200 6536 15000 6656 6 ext_trim[17]
port 19 nsew signal input
rlabel metal3 s 14200 7352 15000 7472 6 ext_trim[18]
port 20 nsew signal input
rlabel metal3 s 14200 8304 15000 8424 6 ext_trim[19]
port 21 nsew signal input
rlabel metal2 s 2226 14200 2282 15000 6 ext_trim[1]
port 22 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 ext_trim[20]
port 23 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 ext_trim[21]
port 24 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 ext_trim[22]
port 25 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 ext_trim[23]
port 26 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 ext_trim[24]
port 27 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 ext_trim[25]
port 28 nsew signal input
rlabel metal2 s 3698 14200 3754 15000 6 ext_trim[2]
port 29 nsew signal input
rlabel metal2 s 5170 14200 5226 15000 6 ext_trim[3]
port 30 nsew signal input
rlabel metal2 s 6734 14200 6790 15000 6 ext_trim[4]
port 31 nsew signal input
rlabel metal2 s 8206 14200 8262 15000 6 ext_trim[5]
port 32 nsew signal input
rlabel metal2 s 9678 14200 9734 15000 6 ext_trim[6]
port 33 nsew signal input
rlabel metal2 s 11242 14200 11298 15000 6 ext_trim[7]
port 34 nsew signal input
rlabel metal2 s 12714 14200 12770 15000 6 ext_trim[8]
port 35 nsew signal input
rlabel metal2 s 14186 14200 14242 15000 6 ext_trim[9]
port 36 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 osc
port 37 nsew signal input
rlabel metal2 s 938 0 994 800 6 resetb
port 38 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 15000 15000
<< end >>
