* NGSPICE file created from digital_pll.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_2 abstract view
.subckt sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_8 abstract view
.subckt sky130_fd_sc_hd__einvn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_4 abstract view
.subckt sky130_fd_sc_hd__einvn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_1 abstract view
.subckt sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

.subckt digital_pll VGND VPWR clockp[0] clockp[1] dco div[0] div[1] div[2] div[3]
+ div[4] enable ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12] ext_trim[13] ext_trim[14]
+ ext_trim[15] ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19] ext_trim[1] ext_trim[20]
+ ext_trim[21] ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25] ext_trim[2] ext_trim[3]
+ ext_trim[4] ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8] ext_trim[9] osc resetb
X_294_ _315_/B _303_/B _294_/C VGND VGND VPWR VPWR _336_/A sky130_fd_sc_hd__and3_2
X_363_ dco _378_/B VGND VGND VPWR VPWR _363_/Y sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[1\].id.delayint0 ringosc.dstage\[1\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_346_ _298_/X _333_/X _345_/Y ext_trim[20] dco VGND VGND VPWR VPWR _346_/X sky130_fd_sc_hd__a32o_2
X_277_ _385_/Q _280_/A _276_/Y _285_/S VGND VGND VPWR VPWR _385_/D sky130_fd_sc_hd__o211a_2
X_200_ _383_/Q _398_/Q VGND VGND VPWR VPWR _218_/B sky130_fd_sc_hd__xor2_2
X_329_ _315_/B _303_/B _248_/B VGND VGND VPWR VPWR _332_/C sky130_fd_sc_hd__a21o_2
Xringosc.dstage\[11\].id.delayen1 ringosc.dstage\[11\].id.delayen1/A _353_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[11\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[10\].id.delayenb0 ringosc.dstage\[10\].id.delayenb1/A _314_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[9\].id.delayenb0 ringosc.dstage\[9\].id.delayenb1/A _312_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[9\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_293_ dco _298_/C VGND VGND VPWR VPWR _294_/C sky130_fd_sc_hd__and2b_2
X_362_ dco _378_/B VGND VGND VPWR VPWR _362_/Y sky130_fd_sc_hd__nor2_2
X_345_ _393_/Q _345_/B VGND VGND VPWR VPWR _345_/Y sky130_fd_sc_hd__nand2_2
X_276_ _386_/Q _278_/B VGND VGND VPWR VPWR _276_/Y sky130_fd_sc_hd__nand2b_2
X_328_ _328_/A _328_/B VGND VGND VPWR VPWR _336_/B sky130_fd_sc_hd__or2_2
XFILLER_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_259_ _259_/A _259_/B VGND VGND VPWR VPWR _259_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_20_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[9\].id.delayenb1 ringosc.dstage\[9\].id.delayenb1/A _350_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[9\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[10\].id.delayenb1 ringosc.dstage\[10\].id.delayenb1/A _351_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XFILLER_15_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_292_ _324_/A _323_/B VGND VGND VPWR VPWR _303_/B sky130_fd_sc_hd__nand2_2
X_361_ dco _378_/B VGND VGND VPWR VPWR _361_/Y sky130_fd_sc_hd__nor2_2
X_344_ _391_/Q _390_/Q _392_/Q VGND VGND VPWR VPWR _345_/B sky130_fd_sc_hd__o21ai_2
X_275_ _386_/Q _278_/B _285_/S VGND VGND VPWR VPWR _386_/D sky130_fd_sc_hd__o21a_2
XFILLER_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[4\].id.delayen0 ringosc.dstage\[4\].id.delayen0/A _302_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_327_ _392_/Q _327_/B VGND VGND VPWR VPWR _327_/X sky130_fd_sc_hd__or2_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_258_ _261_/A _261_/B _247_/B VGND VGND VPWR VPWR _259_/B sky130_fd_sc_hd__a21oi_2
X_189_ _386_/Q _401_/Q VGND VGND VPWR VPWR _190_/B sky130_fd_sc_hd__or2_2
XANTENNA__310__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[9\].id.delaybuf0 ringosc.dstage\[8\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[10\].id.delaybuf0 ringosc.dstage\[9\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[5\].id.delayenb0 ringosc.dstage\[5\].id.delayenb1/A _305_/X VGND
+ VGND VPWR VPWR ringosc.ibufp10/A sky130_fd_sc_hd__einvn_8
X_291_ _392_/Q _307_/C VGND VGND VPWR VPWR _323_/B sky130_fd_sc_hd__nor2_2
X_360_ dco _378_/B VGND VGND VPWR VPWR _360_/Y sky130_fd_sc_hd__nor2_2
X_343_ dco ext_trim[19] _336_/A _336_/B VGND VGND VPWR VPWR _343_/X sky130_fd_sc_hd__a22o_2
X_274_ _385_/Q _280_/A VGND VGND VPWR VPWR _278_/B sky130_fd_sc_hd__and2_2
Xringosc.dstage\[4\].id.delayen1 ringosc.dstage\[4\].id.delayen1/A _341_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_326_ dco ext_trim[14] _304_/X _322_/X VGND VGND VPWR VPWR _326_/X sky130_fd_sc_hd__a22o_2
X_188_ _386_/Q _401_/Q VGND VGND VPWR VPWR _190_/A sky130_fd_sc_hd__nand2_2
X_257_ _393_/Q _271_/B _255_/X _256_/Y VGND VGND VPWR VPWR _393_/D sky130_fd_sc_hd__o22a_2
X_309_ dco ext_trim[7] _336_/A _308_/X VGND VGND VPWR VPWR _309_/X sky130_fd_sc_hd__a22o_2
XANTENNA__310__A2 ext_trim[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__295__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[9\].id.delaybuf1 ringosc.dstage\[9\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[5\].id.delayenb1 ringosc.dstage\[5\].id.delayenb1/A _342_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[5\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[10\].id.delaybuf1 ringosc.dstage\[10\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_290_ _393_/Q _307_/B _391_/Q VGND VGND VPWR VPWR _315_/B sky130_fd_sc_hd__or3_2
XFILLER_3_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_342_ dco ext_trim[18] _324_/B _296_/Y VGND VGND VPWR VPWR _342_/X sky130_fd_sc_hd__a22o_2
X_273_ _384_/Q _383_/Q _382_/Q VGND VGND VPWR VPWR _280_/A sky130_fd_sc_hd__and3_2
X_325_ _328_/A _349_/B VGND VGND VPWR VPWR _325_/X sky130_fd_sc_hd__or2_2
X_187_ _382_/Q _397_/Q _285_/S VGND VGND VPWR VPWR _397_/D sky130_fd_sc_hd__mux2_1
X_256_ _255_/A _255_/B _271_/B VGND VGND VPWR VPWR _256_/Y sky130_fd_sc_hd__o21ai_2
X_308_ _327_/B _328_/B VGND VGND VPWR VPWR _308_/X sky130_fd_sc_hd__or2_2
X_239_ _388_/Q _387_/Q VGND VGND VPWR VPWR _268_/B sky130_fd_sc_hd__nand2_2
XANTENNA__295__A2 ext_trim[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[5\].id.delaybuf0 ringosc.dstage\[4\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_341_ _325_/X _338_/X _340_/X ext_trim[17] dco VGND VGND VPWR VPWR _341_/X sky130_fd_sc_hd__a32o_2
Xringosc.dstage\[1\].id.delayenb0 ringosc.dstage\[1\].id.delayenb1/A _295_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[1\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XANTENNA__361__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_272_ _387_/Q _238_/X _271_/Y VGND VGND VPWR VPWR _387_/D sky130_fd_sc_hd__o21a_2
Xringosc.dstage\[8\].id.delayint0 ringosc.dstage\[8\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__356__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_324_ _324_/A _324_/B VGND VGND VPWR VPWR _347_/C sky130_fd_sc_hd__or2_2
X_186_ _383_/Q _398_/Q _285_/S VGND VGND VPWR VPWR _398_/D sky130_fd_sc_hd__mux2_1
X_255_ _255_/A _255_/B VGND VGND VPWR VPWR _255_/X sky130_fd_sc_hd__and2_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_307_ _393_/Q _307_/B _307_/C VGND VGND VPWR VPWR _328_/B sky130_fd_sc_hd__or3_2
XFILLER_1_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_238_ _380_/Q _238_/B _238_/C _238_/D VGND VGND VPWR VPWR _238_/X sky130_fd_sc_hd__and4_2
XANTENNA__213__B1 div[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__364__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__359__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[5\].id.delaybuf1 ringosc.dstage\[5\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[1\].id.delayenb1 ringosc.dstage\[1\].id.delayenb1/A _326_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[1\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_340_ _340_/A _340_/B _340_/C VGND VGND VPWR VPWR _340_/X sky130_fd_sc_hd__and3_2
X_271_ _387_/Q _271_/B VGND VGND VPWR VPWR _271_/Y sky130_fd_sc_hd__nand2_2
Xringosc.dstage\[1\].id.delayen0 ringosc.dstage\[1\].id.delayen0/A _295_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
X_323_ _393_/Q _323_/B VGND VGND VPWR VPWR _349_/B sky130_fd_sc_hd__nand2_2
XANTENNA__372__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_185_ _384_/Q _399_/Q _285_/S VGND VGND VPWR VPWR _399_/D sky130_fd_sc_hd__mux2_1
X_254_ _393_/Q _269_/A VGND VGND VPWR VPWR _255_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__367__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_306_ dco ext_trim[6] _332_/A _298_/X VGND VGND VPWR VPWR _306_/X sky130_fd_sc_hd__a22o_2
X_237_ _237_/A _237_/B _237_/C VGND VGND VPWR VPWR _238_/D sky130_fd_sc_hd__or3_2
XANTENNA__313__A_N ext_trim[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__222__B2 div[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__222__A1 div[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__289__A1 ext_trim[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__213__A1 div[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__375__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__334__B1 ext_trim[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_270_ _388_/Q _269_/Y _271_/B VGND VGND VPWR VPWR _388_/D sky130_fd_sc_hd__mux2_1
XANTENNA__316__B1 ext_trim[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[1\].id.delayen1 ringosc.dstage\[1\].id.delayen1/A _326_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_399_ _401_/CLK _399_/D _376_/Y VGND VGND VPWR VPWR _399_/Q sky130_fd_sc_hd__dfrtp_2
X_322_ _393_/Q _307_/B _320_/X _321_/Y VGND VGND VPWR VPWR _322_/X sky130_fd_sc_hd__o211a_2
Xringosc.dstage\[1\].id.delaybuf0 ringosc.dstage\[0\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[4\].id.delayint0 ringosc.dstage\[4\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_184_ _385_/Q _400_/Q _285_/S VGND VGND VPWR VPWR _400_/D sky130_fd_sc_hd__mux2_1
X_253_ _259_/A _261_/A _261_/B _324_/B _269_/A VGND VGND VPWR VPWR _255_/A sky130_fd_sc_hd__a32o_2
X_305_ dco ext_trim[5] _304_/X VGND VGND VPWR VPWR _305_/X sky130_fd_sc_hd__a21o_2
X_236_ _236_/A _236_/B _207_/X VGND VGND VPWR VPWR _237_/C sky130_fd_sc_hd__or3b_2
XANTENNA__289__A2 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__378__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__288__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_219_ div[1] _219_/B VGND VGND VPWR VPWR _223_/A sky130_fd_sc_hd__nand2_2
Xringosc.dstage\[9\].id.delayen0 ringosc.dstage\[9\].id.delayen0/A _312_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_16_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__343__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__334__B2 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__316__B2 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_398_ _401_/CLK _398_/D _375_/Y VGND VGND VPWR VPWR _398_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[1\].id.delaybuf1 ringosc.dstage\[1\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_321_ _393_/Q _328_/A _323_/B VGND VGND VPWR VPWR _321_/Y sky130_fd_sc_hd__o21ai_2
X_183_ _386_/Q _401_/Q _285_/S VGND VGND VPWR VPWR _401_/D sky130_fd_sc_hd__mux2_1
X_252_ _339_/A _266_/A _266_/B _327_/B _269_/A VGND VGND VPWR VPWR _261_/B sky130_fd_sc_hd__a32o_2
XFILLER_13_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__225__B1 div[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_304_ _339_/A _303_/B _294_/C _303_/X VGND VGND VPWR VPWR _304_/X sky130_fd_sc_hd__o211a_2
X_235_ div[0] _235_/B VGND VGND VPWR VPWR _236_/A sky130_fd_sc_hd__and2_2
X_218_ _218_/A _218_/B VGND VGND VPWR VPWR _219_/B sky130_fd_sc_hd__xnor2_2
Xringosc.dstage\[9\].id.delayen1 ringosc.dstage\[9\].id.delayen1/A _350_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__343__A2 ext_trim[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__296__B dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_397_ _401_/CLK _397_/D _374_/Y VGND VGND VPWR VPWR _397_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_320_ _392_/Q _327_/B _391_/Q _324_/A VGND VGND VPWR VPWR _320_/X sky130_fd_sc_hd__a211o_2
X_182_ _396_/D _396_/Q VGND VGND VPWR VPWR _287_/B sky130_fd_sc_hd__xor2_2
X_251_ _269_/A _268_/A _268_/B VGND VGND VPWR VPWR _266_/B sky130_fd_sc_hd__a21bo_2
X_303_ _327_/B _303_/B VGND VGND VPWR VPWR _303_/X sky130_fd_sc_hd__or2_2
X_234_ _381_/Q _379_/Q _287_/B VGND VGND VPWR VPWR _238_/C sky130_fd_sc_hd__and3_2
XANTENNA__207__A1 div[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.iss.reseten0 ringosc.iss.const1/HI _378_/B VGND VGND VPWR VPWR ringosc.ibufp00/A
+ sky130_fd_sc_hd__einvp_1
Xringosc.dstage\[0\].id.delayint0 ringosc.dstage\[0\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_217_ _226_/A _217_/B _217_/C VGND VGND VPWR VPWR _237_/A sky130_fd_sc_hd__or3_2
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__346__B1 ext_trim[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[8\].id.delayenb0 ringosc.dstage\[8\].id.delayenb1/A _310_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[8\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
X_396_ _401_/CLK _396_/D _373_/Y VGND VGND VPWR VPWR _396_/Q sky130_fd_sc_hd__dfrtp_2
X_181_ _396_/D _396_/Q VGND VGND VPWR VPWR _285_/S sky130_fd_sc_hd__xnor2_2
X_250_ _347_/B _269_/A VGND VGND VPWR VPWR _266_/A sky130_fd_sc_hd__xnor2_2
X_379_ _401_/CLK _379_/D _356_/Y VGND VGND VPWR VPWR _379_/Q sky130_fd_sc_hd__dfrtp_2
X_302_ dco ext_trim[4] _340_/A VGND VGND VPWR VPWR _302_/X sky130_fd_sc_hd__a21o_2
X_233_ _388_/Q _387_/Q _269_/A _288_/B VGND VGND VPWR VPWR _238_/B sky130_fd_sc_hd__or4bb_2
X_216_ div[2] _216_/B VGND VGND VPWR VPWR _217_/C sky130_fd_sc_hd__nor2_2
Xringosc.iss.delayint0 ringosc.iss.delayen1/Z VGND VGND VPWR VPWR ringosc.iss.delayen0/A
+ sky130_fd_sc_hd__clkinv_1
XANTENNA__346__B2 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__337__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__319__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[8\].id.delayenb1 ringosc.dstage\[8\].id.delayenb1/A _348_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[8\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_395_ _401_/CLK _395_/D _372_/Y VGND VGND VPWR VPWR _396_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_4_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_180_ _389_/Q VGND VGND VPWR VPWR _347_/B sky130_fd_sc_hd__inv_2
X_378_ dco _378_/B VGND VGND VPWR VPWR _378_/Y sky130_fd_sc_hd__nor2_2
X_301_ _390_/Q _315_/B _303_/B _294_/C VGND VGND VPWR VPWR _340_/A sky130_fd_sc_hd__o211a_2
X_232_ _388_/Q _387_/Q VGND VGND VPWR VPWR _268_/A sky130_fd_sc_hd__or2_2
XANTENNA__394__D osc VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[6\].id.delayen0 ringosc.dstage\[6\].id.delayen0/A _306_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
X_215_ _211_/Y _212_/X div[3] VGND VGND VPWR VPWR _226_/B sky130_fd_sc_hd__a21o_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__337__A2 ext_trim[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__319__A2 ext_trim[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_394_ _401_/CLK osc _371_/Y VGND VGND VPWR VPWR _395_/D sky130_fd_sc_hd__dfrtp_2
X_377_ dco _378_/B VGND VGND VPWR VPWR _377_/Y sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[8\].id.delaybuf0 ringosc.dstage\[7\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[4\].id.delayenb0 ringosc.dstage\[4\].id.delayenb1/A _302_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[4\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
X_300_ dco ext_trim[3] _294_/C VGND VGND VPWR VPWR _300_/X sky130_fd_sc_hd__a21o_2
X_231_ _327_/B _298_/C VGND VGND VPWR VPWR _288_/B sky130_fd_sc_hd__nor2_2
XANTENNA__352__A_N dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[10\].id.delayen0 ringosc.dstage\[10\].id.delayen0/A _314_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
Xringosc.dstage\[6\].id.delayen1 ringosc.dstage\[6\].id.delayen1/A _343_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_214_ _211_/Y _212_/X div[3] VGND VGND VPWR VPWR _217_/B sky130_fd_sc_hd__a21oi_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_393_ _401_/CLK _393_/D _370_/Y VGND VGND VPWR VPWR _393_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[8\].id.delaybuf1 ringosc.dstage\[8\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[4\].id.delayenb1 ringosc.dstage\[4\].id.delayenb1/A _341_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[4\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_376_ dco _378_/B VGND VGND VPWR VPWR _376_/Y sky130_fd_sc_hd__nor2_2
X_230_ _393_/Q _324_/B VGND VGND VPWR VPWR _298_/C sky130_fd_sc_hd__or2_2
X_359_ dco _378_/B VGND VGND VPWR VPWR _359_/Y sky130_fd_sc_hd__nor2_2
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__300__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[10\].id.delayen1 ringosc.dstage\[10\].id.delayen1/A _351_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ div[3] _211_/Y _212_/X div[2] _216_/B VGND VGND VPWR VPWR _226_/A sky130_fd_sc_hd__a32o_2
XANTENNA__313__B dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_392_ _401_/CLK _392_/D _369_/Y VGND VGND VPWR VPWR _392_/Q sky130_fd_sc_hd__dfrtp_2
X_375_ dco _378_/B VGND VGND VPWR VPWR _375_/Y sky130_fd_sc_hd__nor2_2
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_358_ dco _378_/B VGND VGND VPWR VPWR _358_/Y sky130_fd_sc_hd__nor2_2
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[4\].id.delaybuf0 ringosc.dstage\[3\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_289_ ext_trim[0] dco _332_/A VGND VGND VPWR VPWR _289_/X sky130_fd_sc_hd__a21o_2
XANTENNA__300__A2 ext_trim[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[7\].id.delayint0 ringosc.dstage\[7\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_212_ _211_/A _211_/B _211_/C VGND VGND VPWR VPWR _212_/X sky130_fd_sc_hd__a21o_2
Xringosc.dstage\[0\].id.delayenb0 ringosc.dstage\[0\].id.delayenb1/A _289_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[0\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_391_ _401_/CLK _391_/D _368_/Y VGND VGND VPWR VPWR _391_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_13_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_374_ dco _378_/B VGND VGND VPWR VPWR _374_/Y sky130_fd_sc_hd__nor2_2
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[3\].id.delayen0 ringosc.dstage\[3\].id.delayen0/A _300_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_357_ dco _378_/B VGND VGND VPWR VPWR _357_/Y sky130_fd_sc_hd__nor2_2
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_288_ dco _288_/B VGND VGND VPWR VPWR _332_/A sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[4\].id.delaybuf1 ringosc.dstage\[4\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_211_ _211_/A _211_/B _211_/C VGND VGND VPWR VPWR _211_/Y sky130_fd_sc_hd__nand3_2
Xringosc.dstage\[0\].id.delayenb1 ringosc.dstage\[0\].id.delayenb1/A _319_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[0\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.iss.delayenb0 ringosc.iss.delayenb1/A ringosc.iss.ctrlen0/X VGND VGND VPWR
+ VPWR ringosc.ibufp00/A sky130_fd_sc_hd__einvn_8
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_390_ _401_/CLK _390_/D _367_/Y VGND VGND VPWR VPWR _390_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__312__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_373_ dco _378_/B VGND VGND VPWR VPWR _373_/Y sky130_fd_sc_hd__nor2_2
X_356_ dco _378_/B VGND VGND VPWR VPWR _356_/Y sky130_fd_sc_hd__nor2_2
X_287_ _379_/Q _287_/B VGND VGND VPWR VPWR _379_/D sky130_fd_sc_hd__or2_2
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[3\].id.delayen1 ringosc.dstage\[3\].id.delayen1/A _337_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_210_ _210_/A _210_/B VGND VGND VPWR VPWR _211_/C sky130_fd_sc_hd__or2_2
X_339_ _339_/A _347_/C VGND VGND VPWR VPWR _340_/C sky130_fd_sc_hd__or2_2
Xringosc.dstage\[0\].id.delaybuf0 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.dstage\[0\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
Xringosc.iss.delayenb1 ringosc.iss.delayenb1/A _354_/X VGND VGND VPWR VPWR ringosc.iss.delayen1/Z
+ sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[3\].id.delayint0 ringosc.dstage\[3\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_372_ dco _378_/B VGND VGND VPWR VPWR _372_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__362__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__312__A2 ext_trim[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__357__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_286_ _380_/Q _379_/Q _287_/B VGND VGND VPWR VPWR _380_/D sky130_fd_sc_hd__mux2_1
X_355_ enable resetb VGND VGND VPWR VPWR _378_/B sky130_fd_sc_hd__nand2_2
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_338_ _265_/A _315_/B _347_/C _248_/B _336_/B VGND VGND VPWR VPWR _338_/X sky130_fd_sc_hd__o221a_2
X_269_ _269_/A _269_/B VGND VGND VPWR VPWR _269_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__370__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[0\].id.delaybuf1 ringosc.dstage\[0\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__365__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.iss.delaybuf0 ringosc.iss.delayenb1/A VGND VGND VPWR VPWR ringosc.iss.delayen1/A
+ sky130_fd_sc_hd__clkbuf_1
X_371_ dco _378_/B VGND VGND VPWR VPWR _371_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__373__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_285_ _380_/Q _381_/Q _285_/S VGND VGND VPWR VPWR _381_/D sky130_fd_sc_hd__mux2_1
X_354_ dco ext_trim[25] _336_/X _340_/C VGND VGND VPWR VPWR _354_/X sky130_fd_sc_hd__a22o_2
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__368__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_337_ dco ext_trim[16] _336_/X VGND VGND VPWR VPWR _337_/X sky130_fd_sc_hd__a21o_2
X_199_ _382_/Q _397_/Q VGND VGND VPWR VPWR _221_/A sky130_fd_sc_hd__nand2_2
X_268_ _268_/A _268_/B VGND VGND VPWR VPWR _269_/B sky130_fd_sc_hd__nand2_2
XANTENNA__351__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__342__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__376__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__306__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_370_ dco _378_/B VGND VGND VPWR VPWR _370_/Y sky130_fd_sc_hd__nor2_2
X_284_ _382_/Q _285_/S _284_/C VGND VGND VPWR VPWR _382_/D sky130_fd_sc_hd__nand3_2
X_353_ dco ext_trim[24] _352_/X VGND VGND VPWR VPWR _353_/X sky130_fd_sc_hd__a21o_2
XANTENNA__215__B1 div[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[0\].id.delayen0 ringosc.dstage\[0\].id.delayen0/A _289_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_336_ _336_/A _336_/B _340_/B VGND VGND VPWR VPWR _336_/X sky130_fd_sc_hd__and3_2
Xringosc.dstage\[7\].id.delayenb0 ringosc.dstage\[7\].id.delayenb1/A _309_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[7\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
X_198_ _382_/Q _397_/Q VGND VGND VPWR VPWR _218_/A sky130_fd_sc_hd__and2_2
X_267_ _271_/B _266_/Y _389_/Q _238_/X VGND VGND VPWR VPWR _389_/D sky130_fd_sc_hd__o2bb2a_2
X_319_ dco ext_trim[13] _336_/A _318_/X VGND VGND VPWR VPWR _319_/X sky130_fd_sc_hd__a22o_2
XANTENNA__351__A2 ext_trim[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__342__A2 ext_trim[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__306__A2 ext_trim[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[0\].id.delayen1 ringosc.dstage\[0\].id.delayen1/A _319_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ _284_/C _282_/Y _287_/B VGND VGND VPWR VPWR _383_/D sky130_fd_sc_hd__a21oi_2
X_352_ dco _392_/Q _393_/Q VGND VGND VPWR VPWR _352_/X sky130_fd_sc_hd__and3b_2
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[7\].id.delayenb1 ringosc.dstage\[7\].id.delayenb1/A _346_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[7\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_335_ _248_/B _328_/B _347_/C _327_/B VGND VGND VPWR VPWR _340_/B sky130_fd_sc_hd__o22a_2
X_197_ _383_/Q _398_/Q VGND VGND VPWR VPWR _197_/X sky130_fd_sc_hd__and2_2
X_266_ _266_/A _266_/B VGND VGND VPWR VPWR _266_/Y sky130_fd_sc_hd__xnor2_2
X_249_ _389_/Q _269_/A VGND VGND VPWR VPWR _249_/Y sky130_fd_sc_hd__nor2_2
X_318_ _390_/Q _328_/B VGND VGND VPWR VPWR _318_/X sky130_fd_sc_hd__or2_2
Xringosc.dstage\[8\].id.delayen0 ringosc.dstage\[8\].id.delayen0/A _310_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[8\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclockp_buffer_0 _401_/CLK VGND VGND VPWR VPWR clockp[0] sky130_fd_sc_hd__clkbuf_16
X_282_ _383_/Q _382_/Q VGND VGND VPWR VPWR _282_/Y sky130_fd_sc_hd__xnor2_2
X_351_ dco ext_trim[23] _296_/Y VGND VGND VPWR VPWR _351_/X sky130_fd_sc_hd__a21o_2
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_334_ _324_/B _296_/Y _327_/X ext_trim[15] dco VGND VGND VPWR VPWR _334_/X sky130_fd_sc_hd__a32o_2
X_196_ _384_/Q _399_/Q VGND VGND VPWR VPWR _208_/B sky130_fd_sc_hd__and2_2
X_265_ _265_/A _265_/B VGND VGND VPWR VPWR _390_/D sky130_fd_sc_hd__xnor2_2
XANTENNA__354__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_317_ dco ext_trim[12] _294_/C _297_/X VGND VGND VPWR VPWR _317_/X sky130_fd_sc_hd__a22o_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_248_ _327_/B _248_/B VGND VGND VPWR VPWR _339_/A sky130_fd_sc_hd__nand2_2
X_179_ _390_/Q VGND VGND VPWR VPWR _265_/A sky130_fd_sc_hd__inv_2
Xringosc.dstage\[7\].id.delaybuf0 ringosc.dstage\[6\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[3\].id.delayenb0 ringosc.dstage\[3\].id.delayenb1/A _300_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[3\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[11\].id.delayint0 ringosc.dstage\[11\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_11_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xringosc.dstage\[8\].id.delayen1 ringosc.dstage\[8\].id.delayen1/A _348_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[8\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_8_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclockp_buffer_1 ringosc.ibufp11/Y VGND VGND VPWR VPWR clockp[1] sky130_fd_sc_hd__clkbuf_16
XANTENNA__309__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_350_ _338_/X _340_/X _349_/X ext_trim[22] dco VGND VGND VPWR VPWR _350_/X sky130_fd_sc_hd__a32o_2
X_281_ _284_/C _280_/X _287_/B VGND VGND VPWR VPWR _384_/D sky130_fd_sc_hd__a21oi_2
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_333_ _333_/A _333_/B _333_/C VGND VGND VPWR VPWR _333_/X sky130_fd_sc_hd__and3_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_195_ _384_/Q _399_/Q VGND VGND VPWR VPWR _211_/A sky130_fd_sc_hd__or2_2
X_264_ _347_/B _266_/B _263_/Y _271_/B VGND VGND VPWR VPWR _265_/B sky130_fd_sc_hd__o211a_2
X_316_ _303_/B _294_/C _315_/X ext_trim[11] dco VGND VGND VPWR VPWR _316_/X sky130_fd_sc_hd__a32o_2
X_247_ _247_/A _247_/B VGND VGND VPWR VPWR _261_/A sky130_fd_sc_hd__nor2_2
XANTENNA__354__A2 ext_trim[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[7\].id.delaybuf1 ringosc.dstage\[7\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[3\].id.delayenb1 ringosc.dstage\[3\].id.delayenb1/A _337_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[3\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_178_ _391_/Q VGND VGND VPWR VPWR _307_/C sky130_fd_sc_hd__inv_2
XANTENNA__309__A2 ext_trim[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_280_ _280_/A _280_/B VGND VGND VPWR VPWR _280_/X sky130_fd_sc_hd__or2_2
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_332_ _332_/A _336_/B _332_/C VGND VGND VPWR VPWR _333_/C sky130_fd_sc_hd__and3_2
X_194_ _384_/Q _399_/Q VGND VGND VPWR VPWR _208_/A sky130_fd_sc_hd__nor2_2
X_401_ _401_/CLK _401_/D _378_/Y VGND VGND VPWR VPWR _401_/Q sky130_fd_sc_hd__dfrtp_2
X_263_ _269_/A _268_/A _249_/Y VGND VGND VPWR VPWR _263_/Y sky130_fd_sc_hd__a21oi_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_315_ _328_/A _315_/B VGND VGND VPWR VPWR _315_/X sky130_fd_sc_hd__or2_2
X_177_ _392_/Q VGND VGND VPWR VPWR _307_/B sky130_fd_sc_hd__inv_2
X_246_ _391_/Q _269_/A VGND VGND VPWR VPWR _247_/B sky130_fd_sc_hd__and2_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_229_ _392_/Q _391_/Q VGND VGND VPWR VPWR _324_/B sky130_fd_sc_hd__or2_2
Xringosc.dstage\[3\].id.delaybuf0 ringosc.dstage\[2\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[6\].id.delayint0 ringosc.dstage\[6\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__216__A div[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.ibufp10 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.ibufp11/A sky130_fd_sc_hd__clkinv_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ _339_/A _303_/B _328_/B _248_/B VGND VGND VPWR VPWR _333_/B sky130_fd_sc_hd__o22a_2
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_193_ _385_/Q _400_/Q VGND VGND VPWR VPWR _210_/B sky130_fd_sc_hd__and2_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_262_ _391_/Q _261_/X _271_/B VGND VGND VPWR VPWR _391_/D sky130_fd_sc_hd__mux2_1
X_400_ _401_/CLK _400_/D _377_/Y VGND VGND VPWR VPWR _400_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__348__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_176_ _393_/Q VGND VGND VPWR VPWR _324_/A sky130_fd_sc_hd__inv_2
X_314_ dco _298_/C _328_/A _313_/Y VGND VGND VPWR VPWR _314_/X sky130_fd_sc_hd__o31a_2
X_245_ _391_/Q _269_/A VGND VGND VPWR VPWR _247_/A sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[5\].id.delayen0 ringosc.dstage\[5\].id.delayen0/A _305_/X VGND VGND
+ VPWR VPWR ringosc.ibufp10/A sky130_fd_sc_hd__einvp_2
Xringosc.dstage\[3\].id.delaybuf1 ringosc.dstage\[3\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_228_ _390_/Q _389_/Q VGND VGND VPWR VPWR _327_/B sky130_fd_sc_hd__or2_2
XFILLER_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__219__A div[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.ibufp00 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.ibufp01/A sky130_fd_sc_hd__clkinv_2
Xringosc.ibufp11 ringosc.ibufp11/A VGND VGND VPWR VPWR ringosc.ibufp11/Y sky130_fd_sc_hd__clkinv_8
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ _265_/A _298_/C _303_/X _315_/X VGND VGND VPWR VPWR _333_/A sky130_fd_sc_hd__o211a_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_192_ _210_/A VGND VGND VPWR VPWR _192_/Y sky130_fd_sc_hd__inv_2
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ _261_/A _261_/B VGND VGND VPWR VPWR _261_/X sky130_fd_sc_hd__xor2_2
XANTENNA__348__A2 ext_trim[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__293__A_N dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_313_ ext_trim[10] dco VGND VGND VPWR VPWR _313_/Y sky130_fd_sc_hd__nand2b_2
X_244_ _307_/B _269_/A VGND VGND VPWR VPWR _259_/A sky130_fd_sc_hd__xnor2_2
Xringosc.dstage\[5\].id.delayen1 ringosc.dstage\[5\].id.delayen1/A _342_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[5\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_227_ _224_/Y _237_/B _226_/X _207_/X VGND VGND VPWR VPWR _269_/A sky130_fd_sc_hd__o31a_2
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__235__A div[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[2\].id.delayint0 ringosc.dstage\[2\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.ibufp01 ringosc.ibufp01/A VGND VGND VPWR VPWR _401_/CLK sky130_fd_sc_hd__clkinv_8
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ _392_/Q _259_/Y _271_/B VGND VGND VPWR VPWR _392_/D sky130_fd_sc_hd__mux2_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_389_ _401_/CLK _389_/D _366_/Y VGND VGND VPWR VPWR _389_/Q sky130_fd_sc_hd__dfrtp_2
X_191_ _385_/Q _400_/Q VGND VGND VPWR VPWR _210_/A sky130_fd_sc_hd__nor2_2
X_312_ dco ext_trim[9] _304_/X _311_/X VGND VGND VPWR VPWR _312_/X sky130_fd_sc_hd__a22o_2
X_243_ _307_/B _269_/A _242_/X _238_/X VGND VGND VPWR VPWR _271_/B sky130_fd_sc_hd__o31a_2
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_226_ _226_/A _226_/B VGND VGND VPWR VPWR _226_/X sky130_fd_sc_hd__and2_2
XFILLER_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xringosc.dstage\[11\].id.delayenb0 ringosc.dstage\[11\].id.delayenb1/A _316_/X VGND
+ VGND VPWR VPWR ringosc.iss.delayenb1/A sky130_fd_sc_hd__einvn_8
X_209_ _209_/A _209_/B VGND VGND VPWR VPWR _216_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__302__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_190_ _190_/A _190_/B VGND VGND VPWR VPWR _206_/A sky130_fd_sc_hd__and2_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_388_ _401_/CLK _388_/D _365_/Y VGND VGND VPWR VPWR _388_/Q sky130_fd_sc_hd__dfrtp_2
X_311_ _327_/B _315_/B _303_/B _248_/B VGND VGND VPWR VPWR _311_/X sky130_fd_sc_hd__o22a_2
X_242_ _324_/A _307_/C _268_/B _248_/B VGND VGND VPWR VPWR _242_/X sky130_fd_sc_hd__or4_2
XFILLER_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[11\].id.delayenb1 ringosc.dstage\[11\].id.delayenb1/A _353_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[11\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_225_ _204_/Y _205_/X div[4] VGND VGND VPWR VPWR _237_/B sky130_fd_sc_hd__o21a_2
X_208_ _208_/A _208_/B VGND VGND VPWR VPWR _209_/B sky130_fd_sc_hd__nor2_2
XANTENNA__302__A2 ext_trim[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_387_ _401_/CLK _387_/D _364_/Y VGND VGND VPWR VPWR _387_/Q sky130_fd_sc_hd__dfrtp_2
X_310_ dco ext_trim[8] _294_/C _303_/X VGND VGND VPWR VPWR _310_/X sky130_fd_sc_hd__a22o_2
XANTENNA__360__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[2\].id.delayen0 ringosc.dstage\[2\].id.delayen0/A _299_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
Xringosc.iss.const1 VGND VGND VPWR VPWR ringosc.iss.const1/HI ringosc.iss.const1/LO
+ sky130_fd_sc_hd__conb_1
X_241_ _390_/Q _389_/Q VGND VGND VPWR VPWR _248_/B sky130_fd_sc_hd__nand2_2
XANTENNA__355__A enable VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__341__B1 ext_trim[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__350__B1 ext_trim[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_224_ _223_/A _236_/B _226_/A _217_/B _217_/C VGND VGND VPWR VPWR _224_/Y sky130_fd_sc_hd__a2111oi_2
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[6\].id.delayenb0 ringosc.dstage\[6\].id.delayenb1/A _306_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[6\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[11\].id.delaybuf0 ringosc.dstage\[10\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_207_ div[4] _204_/Y _206_/Y _190_/A VGND VGND VPWR VPWR _207_/X sky130_fd_sc_hd__o211a_2
XANTENNA__363__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__358__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_386_ _401_/CLK _386_/D _363_/Y VGND VGND VPWR VPWR _386_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[2\].id.delayen1 ringosc.dstage\[2\].id.delayen1/A _334_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_240_ _265_/A _347_/B VGND VGND VPWR VPWR _328_/A sky130_fd_sc_hd__nor2_2
XANTENNA__355__B resetb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_369_ dco _378_/B VGND VGND VPWR VPWR _369_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__350__B2 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_223_ _223_/A _223_/B VGND VGND VPWR VPWR _236_/B sky130_fd_sc_hd__nand2_2
XANTENNA__371__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__341__B2 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__366__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__314__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[6\].id.delayenb1 ringosc.dstage\[6\].id.delayenb1/A _343_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[6\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_206_ _206_/A _206_/B VGND VGND VPWR VPWR _206_/Y sky130_fd_sc_hd__nand2_2
Xringosc.dstage\[11\].id.delaybuf1 ringosc.dstage\[11\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__305__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__214__B1 div[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__374__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_385_ _401_/CLK _385_/D _362_/Y VGND VGND VPWR VPWR _385_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.iss.delayen0 ringosc.iss.delayen0/A _317_/X VGND VGND VPWR VPWR ringosc.ibufp00/A
+ sky130_fd_sc_hd__einvp_2
XANTENNA__369__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_299_ dco ext_trim[2] _303_/B _294_/C VGND VGND VPWR VPWR _299_/X sky130_fd_sc_hd__a22o_2
X_368_ dco _378_/B VGND VGND VPWR VPWR _368_/Y sky130_fd_sc_hd__nor2_2
X_222_ div[1] _219_/B _235_/B div[0] VGND VGND VPWR VPWR _223_/B sky130_fd_sc_hd__o22a_2
XFILLER_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_205_ _206_/A _206_/B VGND VGND VPWR VPWR _205_/X sky130_fd_sc_hd__and2_2
XANTENNA__305__A2 ext_trim[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__377__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__299__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[6\].id.delaybuf0 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.dstage\[6\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[2\].id.delayenb0 ringosc.dstage\[2\].id.delayenb1/A _299_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[2\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[9\].id.delayint0 ringosc.dstage\[9\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[10\].id.delayint0 ringosc.dstage\[10\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_384_ _401_/CLK _384_/D _361_/Y VGND VGND VPWR VPWR _384_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.iss.delayen1 ringosc.iss.delayen1/A _354_/X VGND VGND VPWR VPWR ringosc.iss.delayen1/Z
+ sky130_fd_sc_hd__einvp_2
X_298_ _390_/Q _347_/B _298_/C VGND VGND VPWR VPWR _298_/X sky130_fd_sc_hd__or3_2
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_367_ dco _378_/B VGND VGND VPWR VPWR _367_/Y sky130_fd_sc_hd__nor2_2
X_221_ _221_/A _221_/B VGND VGND VPWR VPWR _235_/B sky130_fd_sc_hd__nand2_2
X_204_ _206_/A _206_/B VGND VGND VPWR VPWR _204_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__299__A2 ext_trim[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[6\].id.delaybuf1 ringosc.dstage\[6\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[2\].id.delayenb1 ringosc.dstage\[2\].id.delayenb1/A _334_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[2\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_383_ _401_/CLK _383_/D _360_/Y VGND VGND VPWR VPWR _383_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__353__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_297_ _390_/Q _303_/B VGND VGND VPWR VPWR _297_/X sky130_fd_sc_hd__or2_2
X_366_ dco _378_/B VGND VGND VPWR VPWR _366_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__326__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_220_ _382_/Q _397_/Q VGND VGND VPWR VPWR _221_/B sky130_fd_sc_hd__or2_2
X_349_ _390_/Q _349_/B VGND VGND VPWR VPWR _349_/X sky130_fd_sc_hd__or2_2
XANTENNA__317__A1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_203_ _192_/Y _211_/A _211_/B _210_/B VGND VGND VPWR VPWR _206_/B sky130_fd_sc_hd__a31o_2
Xringosc.iss.ctrlen0 _378_/B _317_/X VGND VGND VPWR VPWR ringosc.iss.ctrlen0/X sky130_fd_sc_hd__or2_2
XFILLER_18_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[2\].id.delaybuf0 ringosc.dstage\[1\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[5\].id.delayint0 ringosc.dstage\[5\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_382_ _401_/CLK _382_/D _359_/Y VGND VGND VPWR VPWR _382_/Q sky130_fd_sc_hd__dfrtp_2
X_296_ _324_/A dco VGND VGND VPWR VPWR _296_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__353__A2 ext_trim[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_365_ dco _378_/B VGND VGND VPWR VPWR _365_/Y sky130_fd_sc_hd__nor2_2
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__326__A2 ext_trim[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_348_ dco ext_trim[21] _336_/X _347_/X VGND VGND VPWR VPWR _348_/X sky130_fd_sc_hd__a22o_2
XANTENNA__317__A2 ext_trim[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_279_ _383_/Q _382_/Q _384_/Q VGND VGND VPWR VPWR _280_/B sky130_fd_sc_hd__a21oi_2
X_202_ _218_/A _218_/B _208_/B _197_/X VGND VGND VPWR VPWR _211_/B sky130_fd_sc_hd__a211o_2
Xringosc.dstage\[7\].id.delayen0 ringosc.dstage\[7\].id.delayen0/A _309_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[7\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[2\].id.delaybuf1 ringosc.dstage\[2\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_381_ _401_/CLK _381_/D _358_/Y VGND VGND VPWR VPWR _381_/Q sky130_fd_sc_hd__dfrtp_2
X_295_ dco ext_trim[1] _336_/A VGND VGND VPWR VPWR _295_/X sky130_fd_sc_hd__a21o_2
XFILLER_3_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_364_ dco _378_/B VGND VGND VPWR VPWR _364_/Y sky130_fd_sc_hd__nor2_2
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_347_ _390_/Q _347_/B _347_/C VGND VGND VPWR VPWR _347_/X sky130_fd_sc_hd__or3_2
X_278_ _386_/Q _278_/B VGND VGND VPWR VPWR _284_/C sky130_fd_sc_hd__nand2_2
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_201_ _218_/A _218_/B _197_/X VGND VGND VPWR VPWR _209_/A sky130_fd_sc_hd__a21o_2
Xringosc.dstage\[11\].id.delayen0 ringosc.dstage\[11\].id.delayen0/A _316_/X VGND
+ VGND VPWR VPWR ringosc.iss.delayenb1/A sky130_fd_sc_hd__einvp_2
Xringosc.dstage\[7\].id.delayen1 ringosc.dstage\[7\].id.delayen1/A _346_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[7\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_380_ _401_/CLK _380_/D _357_/Y VGND VGND VPWR VPWR _380_/Q sky130_fd_sc_hd__dfrtp_2
.ends

