magic
tech sky130A
magscale 1 2
timestamp 1638876627
<< locali >>
rect 14473 9367 14507 9605
rect 13921 5627 13955 5729
rect 15485 3451 15519 3621
rect 2329 2839 2363 3077
rect 8493 2295 8527 2601
rect 5641 1275 5675 1445
rect 13645 663 13679 833
<< viali >>
rect 7297 10761 7331 10795
rect 10057 10761 10091 10795
rect 13921 10761 13955 10795
rect 18337 10761 18371 10795
rect 8309 10693 8343 10727
rect 9045 10693 9079 10727
rect 9137 10693 9171 10727
rect 10885 10693 10919 10727
rect 12357 10693 12391 10727
rect 18153 10693 18187 10727
rect 1961 10625 1995 10659
rect 2145 10625 2179 10659
rect 3893 10625 3927 10659
rect 6285 10625 6319 10659
rect 7481 10625 7515 10659
rect 7941 10625 7975 10659
rect 8125 10625 8159 10659
rect 10241 10625 10275 10659
rect 12449 10625 12483 10659
rect 13737 10625 13771 10659
rect 14105 10625 14139 10659
rect 15025 10625 15059 10659
rect 15669 10625 15703 10659
rect 16957 10625 16991 10659
rect 18061 10625 18095 10659
rect 18245 10625 18279 10659
rect 18521 10625 18555 10659
rect 3801 10557 3835 10591
rect 8953 10557 8987 10591
rect 12265 10557 12299 10591
rect 17877 10557 17911 10591
rect 8585 10489 8619 10523
rect 2053 10421 2087 10455
rect 4261 10421 4295 10455
rect 6285 10421 6319 10455
rect 7757 10421 7791 10455
rect 12817 10421 12851 10455
rect 13461 10421 13495 10455
rect 14473 10421 14507 10455
rect 14933 10421 14967 10455
rect 16313 10421 16347 10455
rect 16957 10421 16991 10455
rect 3433 10217 3467 10251
rect 3893 10217 3927 10251
rect 7895 10217 7929 10251
rect 12633 10217 12667 10251
rect 15071 10217 15105 10251
rect 17831 10217 17865 10251
rect 8585 10149 8619 10183
rect 8861 10149 8895 10183
rect 1685 10081 1719 10115
rect 1961 10081 1995 10115
rect 6101 10081 6135 10115
rect 8953 10081 8987 10115
rect 10885 10081 10919 10115
rect 11161 10081 11195 10115
rect 13277 10081 13311 10115
rect 13645 10081 13679 10115
rect 16037 10081 16071 10115
rect 489 10013 523 10047
rect 949 10013 983 10047
rect 1133 10013 1167 10047
rect 1317 10013 1351 10047
rect 3709 10013 3743 10047
rect 3893 10013 3927 10047
rect 6469 10013 6503 10047
rect 16405 10013 16439 10047
rect 18245 10013 18279 10047
rect 18521 10013 18555 10047
rect 397 9945 431 9979
rect 1409 9945 1443 9979
rect 1593 9945 1627 9979
rect 9229 9945 9263 9979
rect 949 9877 983 9911
rect 1317 9877 1351 9911
rect 4077 9877 4111 9911
rect 5917 9877 5951 9911
rect 10701 9877 10735 9911
rect 13093 9877 13127 9911
rect 15945 9877 15979 9911
rect 18337 9877 18371 9911
rect 2513 9673 2547 9707
rect 3157 9673 3191 9707
rect 5273 9673 5307 9707
rect 6009 9673 6043 9707
rect 6469 9673 6503 9707
rect 11253 9673 11287 9707
rect 11897 9673 11931 9707
rect 3893 9605 3927 9639
rect 5365 9605 5399 9639
rect 6377 9605 6411 9639
rect 6561 9605 6595 9639
rect 12265 9605 12299 9639
rect 14473 9605 14507 9639
rect 17509 9605 17543 9639
rect 305 9537 339 9571
rect 673 9537 707 9571
rect 2099 9537 2133 9571
rect 2513 9537 2547 9571
rect 2605 9537 2639 9571
rect 2789 9537 2823 9571
rect 2881 9537 2915 9571
rect 3249 9537 3283 9571
rect 3617 9537 3651 9571
rect 3801 9537 3835 9571
rect 3985 9537 4019 9571
rect 4077 9537 4111 9571
rect 4261 9537 4295 9571
rect 5733 9537 5767 9571
rect 5917 9537 5951 9571
rect 6285 9537 6319 9571
rect 6837 9537 6871 9571
rect 7481 9537 7515 9571
rect 9965 9537 9999 9571
rect 4169 9469 4203 9503
rect 5457 9469 5491 9503
rect 7573 9469 7607 9503
rect 7849 9469 7883 9503
rect 12541 9469 12575 9503
rect 12817 9469 12851 9503
rect 9321 9401 9355 9435
rect 14289 9401 14323 9435
rect 14749 9537 14783 9571
rect 15117 9537 15151 9571
rect 16543 9537 16577 9571
rect 16865 9537 16899 9571
rect 2237 9333 2271 9367
rect 4905 9333 4939 9367
rect 6193 9333 6227 9367
rect 6745 9333 6779 9367
rect 9781 9333 9815 9367
rect 12173 9333 12207 9367
rect 14473 9333 14507 9367
rect 14657 9333 14691 9367
rect 1041 9129 1075 9163
rect 1409 9129 1443 9163
rect 5641 9129 5675 9163
rect 8493 9129 8527 9163
rect 11897 9129 11931 9163
rect 15485 9129 15519 9163
rect 9689 9061 9723 9095
rect 10517 9061 10551 9095
rect 10885 9061 10919 9095
rect 4353 8993 4387 9027
rect 10333 8993 10367 9027
rect 11437 8993 11471 9027
rect 12541 8993 12575 9027
rect 13277 8993 13311 9027
rect 17601 8993 17635 9027
rect 949 8925 983 8959
rect 1133 8925 1167 8959
rect 1501 8925 1535 8959
rect 2697 8925 2731 8959
rect 2973 8925 3007 8959
rect 4169 8925 4203 8959
rect 5549 8925 5583 8959
rect 5641 8925 5675 8959
rect 6653 8925 6687 8959
rect 6837 8925 6871 8959
rect 7757 8925 7791 8959
rect 7849 8925 7883 8959
rect 8677 8925 8711 8959
rect 8769 8925 8803 8959
rect 9229 8925 9263 8959
rect 10517 8925 10551 8959
rect 10701 8925 10735 8959
rect 11253 8925 11287 8959
rect 12265 8925 12299 8959
rect 12725 8925 12759 8959
rect 13645 8925 13679 8959
rect 15301 8925 15335 8959
rect 15485 8925 15519 8959
rect 17877 8925 17911 8959
rect 5365 8857 5399 8891
rect 6469 8857 6503 8891
rect 6929 8857 6963 8891
rect 7113 8857 7147 8891
rect 9321 8857 9355 8891
rect 9505 8857 9539 8891
rect 10057 8857 10091 8891
rect 12817 8857 12851 8891
rect 13001 8857 13035 8891
rect 15853 8857 15887 8891
rect 3801 8789 3835 8823
rect 4261 8789 4295 8823
rect 7021 8789 7055 8823
rect 7389 8789 7423 8823
rect 8033 8789 8067 8823
rect 9137 8789 9171 8823
rect 9229 8789 9263 8823
rect 10149 8789 10183 8823
rect 11345 8789 11379 8823
rect 12357 8789 12391 8823
rect 12909 8789 12943 8823
rect 15071 8789 15105 8823
rect 15761 8789 15795 8823
rect 2145 8585 2179 8619
rect 3157 8585 3191 8619
rect 3525 8585 3559 8619
rect 3985 8585 4019 8619
rect 6193 8585 6227 8619
rect 8861 8585 8895 8619
rect 10333 8585 10367 8619
rect 10793 8585 10827 8619
rect 10885 8585 10919 8619
rect 12817 8585 12851 8619
rect 13185 8585 13219 8619
rect 13645 8585 13679 8619
rect 17325 8585 17359 8619
rect 5273 8517 5307 8551
rect 6285 8517 6319 8551
rect 7726 8517 7760 8551
rect 14565 8517 14599 8551
rect 17233 8517 17267 8551
rect 2145 8449 2179 8483
rect 2329 8449 2363 8483
rect 2697 8449 2731 8483
rect 4353 8449 4387 8483
rect 5181 8449 5215 8483
rect 5365 8449 5399 8483
rect 5733 8449 5767 8483
rect 6745 8449 6779 8483
rect 9215 8449 9249 8483
rect 9689 8449 9723 8483
rect 11713 8449 11747 8483
rect 12081 8449 12115 8483
rect 12265 8449 12299 8483
rect 12449 8449 12483 8483
rect 12541 8449 12575 8483
rect 12633 8449 12667 8483
rect 12909 8449 12943 8483
rect 13093 8449 13127 8483
rect 13369 8449 13403 8483
rect 13921 8449 13955 8483
rect 14657 8449 14691 8483
rect 18245 8449 18279 8483
rect 18521 8449 18555 8483
rect 305 8381 339 8415
rect 581 8381 615 8415
rect 2605 8381 2639 8415
rect 3617 8381 3651 8415
rect 3709 8381 3743 8415
rect 4445 8381 4479 8415
rect 4537 8381 4571 8415
rect 6009 8381 6043 8415
rect 6837 8381 6871 8415
rect 7113 8381 7147 8415
rect 7481 8381 7515 8415
rect 9137 8381 9171 8415
rect 10701 8381 10735 8415
rect 13829 8381 13863 8415
rect 14841 8381 14875 8415
rect 15209 8381 15243 8415
rect 17417 8381 17451 8415
rect 3065 8313 3099 8347
rect 9505 8313 9539 8347
rect 11253 8313 11287 8347
rect 14289 8313 14323 8347
rect 16865 8313 16899 8347
rect 18337 8313 18371 8347
rect 2053 8245 2087 8279
rect 5825 8245 5859 8279
rect 5917 8245 5951 8279
rect 11621 8245 11655 8279
rect 12081 8245 12115 8279
rect 16635 8245 16669 8279
rect 1409 8041 1443 8075
rect 1501 8041 1535 8075
rect 2421 8041 2455 8075
rect 2513 8041 2547 8075
rect 11805 8041 11839 8075
rect 5641 7973 5675 8007
rect 13369 7973 13403 8007
rect 15761 7973 15795 8007
rect 1317 7905 1351 7939
rect 1869 7905 1903 7939
rect 3065 7905 3099 7939
rect 6653 7905 6687 7939
rect 8861 7905 8895 7939
rect 11437 7905 11471 7939
rect 13001 7905 13035 7939
rect 14381 7905 14415 7939
rect 15209 7905 15243 7939
rect 17509 7905 17543 7939
rect 1593 7837 1627 7871
rect 2881 7837 2915 7871
rect 5457 7837 5491 7871
rect 6285 7837 6319 7871
rect 11253 7837 11287 7871
rect 11713 7837 11747 7871
rect 11897 7837 11931 7871
rect 12725 7837 12759 7871
rect 12909 7837 12943 7871
rect 13921 7837 13955 7871
rect 14473 7837 14507 7871
rect 14657 7837 14691 7871
rect 14933 7837 14967 7871
rect 15301 7837 15335 7871
rect 17877 7837 17911 7871
rect 2053 7769 2087 7803
rect 10609 7769 10643 7803
rect 11989 7769 12023 7803
rect 1961 7701 1995 7735
rect 2973 7701 3007 7735
rect 6193 7701 6227 7735
rect 8079 7701 8113 7735
rect 10885 7701 10919 7735
rect 11345 7701 11379 7735
rect 12541 7701 12575 7735
rect 2145 7497 2179 7531
rect 5549 7497 5583 7531
rect 7481 7497 7515 7531
rect 8493 7497 8527 7531
rect 17049 7497 17083 7531
rect 1961 7429 1995 7463
rect 3893 7429 3927 7463
rect 7389 7429 7423 7463
rect 11345 7429 11379 7463
rect 12541 7429 12575 7463
rect 14197 7429 14231 7463
rect 2053 7361 2087 7395
rect 2145 7361 2179 7395
rect 2329 7361 2363 7395
rect 2697 7361 2731 7395
rect 4077 7361 4111 7395
rect 4169 7361 4203 7395
rect 4261 7361 4295 7395
rect 4445 7361 4479 7395
rect 4905 7361 4939 7395
rect 5068 7367 5102 7401
rect 5181 7364 5215 7398
rect 5319 7361 5353 7395
rect 5917 7361 5951 7395
rect 6101 7361 6135 7395
rect 6929 7361 6963 7395
rect 8033 7361 8067 7395
rect 8861 7361 8895 7395
rect 10425 7361 10459 7395
rect 10885 7361 10919 7395
rect 11069 7361 11103 7395
rect 12357 7361 12391 7395
rect 12449 7361 12483 7395
rect 12633 7361 12667 7395
rect 13553 7361 13587 7395
rect 13737 7361 13771 7395
rect 13829 7361 13863 7395
rect 14032 7361 14066 7395
rect 14289 7361 14323 7395
rect 14473 7361 14507 7395
rect 16267 7361 16301 7395
rect 16957 7361 16991 7395
rect 2605 7293 2639 7327
rect 6469 7293 6503 7327
rect 6837 7293 6871 7327
rect 8125 7293 8159 7327
rect 8309 7293 8343 7327
rect 8953 7293 8987 7327
rect 9045 7293 9079 7327
rect 10517 7293 10551 7327
rect 10701 7293 10735 7327
rect 12081 7293 12115 7327
rect 13645 7293 13679 7327
rect 14841 7293 14875 7327
rect 4169 7225 4203 7259
rect 6101 7225 6135 7259
rect 7665 7225 7699 7259
rect 10057 7225 10091 7259
rect 3065 7157 3099 7191
rect 4261 7157 4295 7191
rect 7113 7157 7147 7191
rect 11437 7157 11471 7191
rect 12173 7157 12207 7191
rect 12265 7157 12299 7191
rect 16405 7157 16439 7191
rect 6377 6953 6411 6987
rect 8045 6953 8079 6987
rect 12357 6953 12391 6987
rect 14105 6953 14139 6987
rect 5917 6885 5951 6919
rect 2237 6817 2271 6851
rect 3341 6817 3375 6851
rect 3893 6817 3927 6851
rect 10885 6817 10919 6851
rect 15393 6817 15427 6851
rect 17877 6817 17911 6851
rect 949 6749 983 6783
rect 1961 6749 1995 6783
rect 2421 6749 2455 6783
rect 2605 6749 2639 6783
rect 4169 6749 4203 6783
rect 4629 6749 4663 6783
rect 4997 6749 5031 6783
rect 5273 6749 5307 6783
rect 6285 6749 6319 6783
rect 6377 6749 6411 6783
rect 8309 6749 8343 6783
rect 8585 6749 8619 6783
rect 10609 6749 10643 6783
rect 12541 6749 12575 6783
rect 12725 6749 12759 6783
rect 14105 6749 14139 6783
rect 14197 6749 14231 6783
rect 15761 6749 15795 6783
rect 18245 6749 18279 6783
rect 18521 6749 18555 6783
rect 2513 6681 2547 6715
rect 3157 6681 3191 6715
rect 6101 6681 6135 6715
rect 8861 6681 8895 6715
rect 11152 6681 11186 6715
rect 14381 6681 14415 6715
rect 14473 6681 14507 6715
rect 15853 6681 15887 6715
rect 17601 6681 17635 6715
rect 765 6613 799 6647
rect 1593 6613 1627 6647
rect 2053 6613 2087 6647
rect 2697 6613 2731 6647
rect 3065 6613 3099 6647
rect 6561 6613 6595 6647
rect 12265 6613 12299 6647
rect 14749 6613 14783 6647
rect 15117 6613 15151 6647
rect 15209 6613 15243 6647
rect 18337 6613 18371 6647
rect 2053 6409 2087 6443
rect 2605 6409 2639 6443
rect 3525 6409 3559 6443
rect 7481 6409 7515 6443
rect 12725 6409 12759 6443
rect 13461 6409 13495 6443
rect 13921 6409 13955 6443
rect 14749 6409 14783 6443
rect 16957 6409 16991 6443
rect 581 6341 615 6375
rect 3985 6341 4019 6375
rect 5641 6341 5675 6375
rect 2513 6273 2547 6307
rect 2697 6273 2731 6307
rect 3433 6273 3467 6307
rect 4169 6273 4203 6307
rect 5733 6273 5767 6307
rect 6469 6273 6503 6307
rect 7665 6273 7699 6307
rect 7849 6273 7883 6307
rect 8033 6273 8067 6307
rect 8585 6273 8619 6307
rect 11897 6273 11931 6307
rect 13829 6273 13863 6307
rect 14749 6273 14783 6307
rect 16865 6273 16899 6307
rect 17325 6273 17359 6307
rect 17693 6273 17727 6307
rect 305 6205 339 6239
rect 3709 6205 3743 6239
rect 4445 6205 4479 6239
rect 5825 6205 5859 6239
rect 6561 6205 6595 6239
rect 6653 6205 6687 6239
rect 7941 6205 7975 6239
rect 12817 6205 12851 6239
rect 13001 6205 13035 6239
rect 14105 6205 14139 6239
rect 14933 6205 14967 6239
rect 15209 6205 15243 6239
rect 16681 6205 16715 6239
rect 5273 6137 5307 6171
rect 12357 6137 12391 6171
rect 2237 6069 2271 6103
rect 3065 6069 3099 6103
rect 4353 6069 4387 6103
rect 6101 6069 6135 6103
rect 8309 6069 8343 6103
rect 8493 6069 8527 6103
rect 8677 6069 8711 6103
rect 9045 6069 9079 6103
rect 9229 6069 9263 6103
rect 11713 6069 11747 6103
rect 3111 5865 3145 5899
rect 6561 5865 6595 5899
rect 8309 5865 8343 5899
rect 10609 5865 10643 5899
rect 16037 5865 16071 5899
rect 4169 5729 4203 5763
rect 6193 5729 6227 5763
rect 6929 5729 6963 5763
rect 11161 5729 11195 5763
rect 13553 5729 13587 5763
rect 13921 5729 13955 5763
rect 14289 5729 14323 5763
rect 15761 5729 15795 5763
rect 15945 5729 15979 5763
rect 16129 5729 16163 5763
rect 17601 5729 17635 5763
rect 1041 5661 1075 5695
rect 1133 5661 1167 5695
rect 1317 5661 1351 5695
rect 1685 5661 1719 5695
rect 6285 5661 6319 5695
rect 7185 5661 7219 5695
rect 10425 5661 10459 5695
rect 13461 5661 13495 5695
rect 14565 5661 14599 5695
rect 15209 5661 15243 5695
rect 16037 5661 16071 5695
rect 17877 5661 17911 5695
rect 18245 5661 18279 5695
rect 18521 5661 18555 5695
rect 4445 5593 4479 5627
rect 11437 5593 11471 5627
rect 13921 5593 13955 5627
rect 14473 5593 14507 5627
rect 3341 5525 3375 5559
rect 3985 5525 4019 5559
rect 5917 5525 5951 5559
rect 9137 5525 9171 5559
rect 11069 5525 11103 5559
rect 12909 5525 12943 5559
rect 13829 5525 13863 5559
rect 14105 5525 14139 5559
rect 14933 5525 14967 5559
rect 15025 5525 15059 5559
rect 15485 5525 15519 5559
rect 18337 5525 18371 5559
rect 1225 5321 1259 5355
rect 2329 5321 2363 5355
rect 2973 5321 3007 5355
rect 4537 5321 4571 5355
rect 4905 5321 4939 5355
rect 5365 5321 5399 5355
rect 6837 5321 6871 5355
rect 11345 5321 11379 5355
rect 12081 5321 12115 5355
rect 6193 5253 6227 5287
rect 6929 5253 6963 5287
rect 11253 5253 11287 5287
rect 16267 5253 16301 5287
rect 1041 5185 1075 5219
rect 1961 5185 1995 5219
rect 2881 5185 2915 5219
rect 3525 5185 3559 5219
rect 4721 5185 4755 5219
rect 5273 5185 5307 5219
rect 5917 5185 5951 5219
rect 8493 5185 8527 5219
rect 9137 5185 9171 5219
rect 9229 5185 9263 5219
rect 9413 5185 9447 5219
rect 10802 5185 10836 5219
rect 11069 5185 11103 5219
rect 11529 5185 11563 5219
rect 11713 5185 11747 5219
rect 13829 5185 13863 5219
rect 14473 5185 14507 5219
rect 16589 5185 16623 5219
rect 17233 5185 17267 5219
rect 2053 5117 2087 5151
rect 3065 5117 3099 5151
rect 3433 5117 3467 5151
rect 5457 5117 5491 5151
rect 8401 5117 8435 5151
rect 13553 5117 13587 5151
rect 14841 5117 14875 5151
rect 17141 5117 17175 5151
rect 2513 5049 2547 5083
rect 8861 5049 8895 5083
rect 9689 5049 9723 5083
rect 16405 5049 16439 5083
rect 16865 5049 16899 5083
rect 3801 4981 3835 5015
rect 9137 4981 9171 5015
rect 11529 4981 11563 5015
rect 11805 4981 11839 5015
rect 14289 4981 14323 5015
rect 8217 4777 8251 4811
rect 10655 4777 10689 4811
rect 5917 4709 5951 4743
rect 4353 4641 4387 4675
rect 4537 4641 4571 4675
rect 4813 4641 4847 4675
rect 5641 4641 5675 4675
rect 6101 4641 6135 4675
rect 6377 4641 6411 4675
rect 8861 4641 8895 4675
rect 9229 4641 9263 4675
rect 11345 4641 11379 4675
rect 11529 4641 11563 4675
rect 13461 4641 13495 4675
rect 16129 4641 16163 4675
rect 17509 4641 17543 4675
rect 857 4573 891 4607
rect 1317 4573 1351 4607
rect 4077 4573 4111 4607
rect 4169 4573 4203 4607
rect 4721 4573 4755 4607
rect 4905 4573 4939 4607
rect 5549 4573 5583 4607
rect 7941 4573 7975 4607
rect 8217 4573 8251 4607
rect 11253 4573 11287 4607
rect 15761 4573 15795 4607
rect 18153 4573 18187 4607
rect 1593 4505 1627 4539
rect 3249 4505 3283 4539
rect 8125 4505 8159 4539
rect 11897 4505 11931 4539
rect 13737 4505 13771 4539
rect 15485 4505 15519 4539
rect 1041 4437 1075 4471
rect 3065 4437 3099 4471
rect 3709 4437 3743 4471
rect 7849 4437 7883 4471
rect 8769 4437 8803 4471
rect 10885 4437 10919 4471
rect 13369 4437 13403 4471
rect 18245 4437 18279 4471
rect 2973 4233 3007 4267
rect 5641 4233 5675 4267
rect 6101 4233 6135 4267
rect 7389 4233 7423 4267
rect 12449 4233 12483 4267
rect 17969 4233 18003 4267
rect 3065 4165 3099 4199
rect 489 4097 523 4131
rect 2329 4097 2363 4131
rect 3801 4097 3835 4131
rect 3893 4097 3927 4131
rect 4537 4097 4571 4131
rect 5641 4097 5675 4131
rect 5733 4097 5767 4131
rect 7297 4097 7331 4131
rect 7481 4097 7515 4131
rect 8861 4097 8895 4131
rect 10609 4097 10643 4131
rect 11253 4097 11287 4131
rect 12357 4097 12391 4131
rect 14197 4097 14231 4131
rect 14473 4097 14507 4131
rect 16635 4097 16669 4131
rect 18245 4097 18279 4131
rect 857 4029 891 4063
rect 3249 4029 3283 4063
rect 3985 4029 4019 4063
rect 5917 4029 5951 4063
rect 8953 4029 8987 4063
rect 10425 4029 10459 4063
rect 11345 4029 11379 4063
rect 13921 4029 13955 4063
rect 14841 4029 14875 4063
rect 15209 4029 15243 4063
rect 16865 4029 16899 4063
rect 17049 4029 17083 4063
rect 2605 3961 2639 3995
rect 11161 3961 11195 3995
rect 3433 3893 3467 3927
rect 4353 3893 4387 3927
rect 14657 3893 14691 3927
rect 1317 3689 1351 3723
rect 3709 3689 3743 3723
rect 5733 3689 5767 3723
rect 11345 3689 11379 3723
rect 14841 3689 14875 3723
rect 18337 3689 18371 3723
rect 4721 3621 4755 3655
rect 8309 3621 8343 3655
rect 15301 3621 15335 3655
rect 15485 3621 15519 3655
rect 4261 3553 4295 3587
rect 6929 3553 6963 3587
rect 7849 3553 7883 3587
rect 8861 3553 8895 3587
rect 11161 3553 11195 3587
rect 13277 3553 13311 3587
rect 14749 3553 14783 3587
rect 1501 3485 1535 3519
rect 3157 3485 3191 3519
rect 3341 3485 3375 3519
rect 4077 3485 4111 3519
rect 4169 3485 4203 3519
rect 4537 3485 4571 3519
rect 4905 3485 4939 3519
rect 5273 3485 5307 3519
rect 6837 3485 6871 3519
rect 8309 3485 8343 3519
rect 8493 3485 8527 3519
rect 10287 3485 10321 3519
rect 11069 3485 11103 3519
rect 12541 3485 12575 3519
rect 12909 3485 12943 3519
rect 13093 3485 13127 3519
rect 15025 3485 15059 3519
rect 15853 3485 15887 3519
rect 18245 3485 18279 3519
rect 18521 3485 18555 3519
rect 3249 3417 3283 3451
rect 5089 3417 5123 3451
rect 8033 3417 8067 3451
rect 8217 3417 8251 3451
rect 13522 3417 13556 3451
rect 15485 3417 15519 3451
rect 16129 3417 16163 3451
rect 17877 3417 17911 3451
rect 2513 3349 2547 3383
rect 6377 3349 6411 3383
rect 6745 3349 6779 3383
rect 12265 3349 12299 3383
rect 13001 3349 13035 3383
rect 14657 3349 14691 3383
rect 15209 3349 15243 3383
rect 15761 3349 15795 3383
rect 8309 3145 8343 3179
rect 8585 3145 8619 3179
rect 16681 3145 16715 3179
rect 2329 3077 2363 3111
rect 2881 3077 2915 3111
rect 11897 3077 11931 3111
rect 305 3009 339 3043
rect 581 2941 615 2975
rect 2053 2941 2087 2975
rect 3709 3009 3743 3043
rect 3801 3009 3835 3043
rect 4169 3009 4203 3043
rect 4353 3009 4387 3043
rect 4629 3009 4663 3043
rect 4905 3009 4939 3043
rect 5181 3009 5215 3043
rect 7297 3009 7331 3043
rect 7389 3009 7423 3043
rect 7573 3009 7607 3043
rect 8033 3009 8067 3043
rect 8217 3009 8251 3043
rect 8769 3009 8803 3043
rect 8861 3009 8895 3043
rect 8953 3009 8987 3043
rect 9873 3009 9907 3043
rect 12081 3009 12115 3043
rect 14013 3009 14047 3043
rect 14657 3009 14691 3043
rect 14841 3009 14875 3043
rect 14933 3009 14967 3043
rect 17049 3009 17083 3043
rect 17601 3009 17635 3043
rect 17785 3009 17819 3043
rect 2973 2941 3007 2975
rect 3157 2941 3191 2975
rect 3985 2941 4019 2975
rect 5457 2941 5491 2975
rect 6929 2941 6963 2975
rect 8493 2941 8527 2975
rect 9781 2941 9815 2975
rect 12449 2941 12483 2975
rect 14289 2941 14323 2975
rect 15209 2941 15243 2975
rect 2513 2873 2547 2907
rect 3341 2873 3375 2907
rect 7297 2873 7331 2907
rect 14105 2873 14139 2907
rect 14473 2873 14507 2907
rect 16865 2873 16899 2907
rect 17509 2873 17543 2907
rect 2237 2805 2271 2839
rect 2329 2805 2363 2839
rect 4537 2805 4571 2839
rect 5089 2805 5123 2839
rect 13875 2805 13909 2839
rect 14197 2805 14231 2839
rect 17141 2805 17175 2839
rect 17969 2805 18003 2839
rect 765 2601 799 2635
rect 2421 2601 2455 2635
rect 3801 2601 3835 2635
rect 6101 2601 6135 2635
rect 6837 2601 6871 2635
rect 8493 2601 8527 2635
rect 9597 2601 9631 2635
rect 11621 2601 11655 2635
rect 13369 2601 13403 2635
rect 17049 2601 17083 2635
rect 17233 2601 17267 2635
rect 17693 2601 17727 2635
rect 2145 2465 2179 2499
rect 2789 2465 2823 2499
rect 3433 2465 3467 2499
rect 6377 2465 6411 2499
rect 6745 2465 6779 2499
rect 7481 2465 7515 2499
rect 949 2397 983 2431
rect 2053 2397 2087 2431
rect 2697 2397 2731 2431
rect 3525 2397 3559 2431
rect 4261 2397 4295 2431
rect 4537 2397 4571 2431
rect 4721 2397 4755 2431
rect 4813 2397 4847 2431
rect 4905 2397 4939 2431
rect 5917 2397 5951 2431
rect 6285 2397 6319 2431
rect 7297 2397 7331 2431
rect 3249 2329 3283 2363
rect 18429 2533 18463 2567
rect 8585 2465 8619 2499
rect 13461 2465 13495 2499
rect 15669 2465 15703 2499
rect 17601 2465 17635 2499
rect 8677 2397 8711 2431
rect 9781 2397 9815 2431
rect 11069 2397 11103 2431
rect 11437 2397 11471 2431
rect 11989 2397 12023 2431
rect 15936 2397 15970 2431
rect 17141 2397 17175 2431
rect 17877 2397 17911 2431
rect 18061 2397 18095 2431
rect 18153 2397 18187 2431
rect 11161 2329 11195 2363
rect 11345 2329 11379 2363
rect 11529 2329 11563 2363
rect 11713 2329 11747 2363
rect 13737 2329 13771 2363
rect 15485 2329 15519 2363
rect 18337 2329 18371 2363
rect 3065 2261 3099 2295
rect 3525 2261 3559 2295
rect 5181 2261 5215 2295
rect 5457 2261 5491 2295
rect 7205 2261 7239 2295
rect 8493 2261 8527 2295
rect 11069 2261 11103 2295
rect 11897 2261 11931 2295
rect 18061 2261 18095 2295
rect 2237 2057 2271 2091
rect 2513 2057 2547 2091
rect 2881 2057 2915 2091
rect 2973 2057 3007 2091
rect 3341 2057 3375 2091
rect 3709 2057 3743 2091
rect 7757 2057 7791 2091
rect 8585 2057 8619 2091
rect 11621 2057 11655 2091
rect 13185 2057 13219 2091
rect 13829 2057 13863 2091
rect 14933 2057 14967 2091
rect 18245 2057 18279 2091
rect 3801 1989 3835 2023
rect 4261 1989 4295 2023
rect 8309 1989 8343 2023
rect 9689 1989 9723 2023
rect 17110 1989 17144 2023
rect 1041 1921 1075 1955
rect 2151 1921 2185 1955
rect 2329 1921 2363 1955
rect 4169 1921 4203 1955
rect 4353 1921 4387 1955
rect 4629 1921 4663 1955
rect 5089 1921 5123 1955
rect 5457 1921 5491 1955
rect 6009 1921 6043 1955
rect 6653 1921 6687 1955
rect 7297 1921 7331 1955
rect 7389 1921 7423 1955
rect 7573 1921 7607 1955
rect 7849 1921 7883 1955
rect 7941 1921 7975 1955
rect 8125 1921 8159 1955
rect 8217 1921 8251 1955
rect 8401 1921 8435 1955
rect 8493 1921 8527 1955
rect 8677 1921 8711 1955
rect 9229 1921 9263 1955
rect 9321 1921 9355 1955
rect 10149 1921 10183 1955
rect 10885 1921 10919 1955
rect 11069 1921 11103 1955
rect 11161 1921 11195 1955
rect 11437 1921 11471 1955
rect 11713 1921 11747 1955
rect 11897 1921 11931 1955
rect 13093 1921 13127 1955
rect 14013 1921 14047 1955
rect 14197 1921 14231 1955
rect 14841 1921 14875 1955
rect 16221 1921 16255 1955
rect 16313 1921 16347 1955
rect 3157 1853 3191 1887
rect 3985 1853 4019 1887
rect 5825 1853 5859 1887
rect 6561 1853 6595 1887
rect 7021 1853 7055 1887
rect 9505 1853 9539 1887
rect 11345 1853 11379 1887
rect 13369 1853 13403 1887
rect 14289 1853 14323 1887
rect 15025 1853 15059 1887
rect 16037 1853 16071 1887
rect 16865 1853 16899 1887
rect 4445 1785 4479 1819
rect 6377 1785 6411 1819
rect 9413 1785 9447 1819
rect 857 1717 891 1751
rect 7297 1717 7331 1751
rect 7849 1717 7883 1751
rect 10425 1717 10459 1751
rect 12725 1717 12759 1751
rect 14473 1717 14507 1751
rect 16681 1717 16715 1751
rect 3065 1513 3099 1547
rect 5917 1513 5951 1547
rect 10057 1513 10091 1547
rect 14749 1513 14783 1547
rect 5641 1445 5675 1479
rect 5365 1377 5399 1411
rect 857 1309 891 1343
rect 1317 1309 1351 1343
rect 3157 1309 3191 1343
rect 4795 1309 4829 1343
rect 5089 1309 5123 1343
rect 6745 1377 6779 1411
rect 7389 1377 7423 1411
rect 7665 1377 7699 1411
rect 9137 1377 9171 1411
rect 11161 1377 11195 1411
rect 12725 1377 12759 1411
rect 15209 1377 15243 1411
rect 15393 1377 15427 1411
rect 5733 1309 5767 1343
rect 5917 1309 5951 1343
rect 6469 1309 6503 1343
rect 7297 1309 7331 1343
rect 8033 1309 8067 1343
rect 8125 1309 8159 1343
rect 8309 1309 8343 1343
rect 9873 1309 9907 1343
rect 10149 1309 10183 1343
rect 10333 1309 10367 1343
rect 10517 1309 10551 1343
rect 11253 1309 11287 1343
rect 11437 1309 11471 1343
rect 13277 1309 13311 1343
rect 13461 1309 13495 1343
rect 14013 1309 14047 1343
rect 14197 1309 14231 1343
rect 14289 1309 14323 1343
rect 16129 1309 16163 1343
rect 1593 1241 1627 1275
rect 3433 1241 3467 1275
rect 5273 1241 5307 1275
rect 5641 1241 5675 1275
rect 10425 1241 10459 1275
rect 10977 1241 11011 1275
rect 12541 1241 12575 1275
rect 16405 1241 16439 1275
rect 581 1173 615 1207
rect 3801 1173 3835 1207
rect 6101 1173 6135 1207
rect 6561 1173 6595 1207
rect 6929 1173 6963 1207
rect 8493 1173 8527 1207
rect 8861 1173 8895 1207
rect 8953 1173 8987 1207
rect 9413 1173 9447 1207
rect 11253 1173 11287 1207
rect 12173 1173 12207 1207
rect 12633 1173 12667 1207
rect 13277 1173 13311 1207
rect 14013 1173 14047 1207
rect 14565 1173 14599 1207
rect 15117 1173 15151 1207
rect 16037 1173 16071 1207
rect 17877 1173 17911 1207
rect 2881 969 2915 1003
rect 2973 969 3007 1003
rect 3341 969 3375 1003
rect 3709 969 3743 1003
rect 6837 969 6871 1003
rect 13921 969 13955 1003
rect 16405 969 16439 1003
rect 16865 969 16899 1003
rect 17325 969 17359 1003
rect 2191 901 2225 935
rect 8861 901 8895 935
rect 12173 901 12207 935
rect 12909 901 12943 935
rect 397 833 431 867
rect 765 833 799 867
rect 4905 833 4939 867
rect 7021 833 7055 867
rect 9137 833 9171 867
rect 9229 833 9263 867
rect 9873 833 9907 867
rect 12081 833 12115 867
rect 12265 833 12299 867
rect 12449 833 12483 867
rect 12817 833 12851 867
rect 13185 833 13219 867
rect 13277 833 13311 867
rect 13369 833 13403 867
rect 13553 833 13587 867
rect 13645 833 13679 867
rect 14013 833 14047 867
rect 14197 833 14231 867
rect 14473 833 14507 867
rect 16589 833 16623 867
rect 16681 833 16715 867
rect 17233 833 17267 867
rect 18245 833 18279 867
rect 3157 765 3191 799
rect 3801 765 3835 799
rect 3985 765 4019 799
rect 5273 765 5307 799
rect 7389 765 7423 799
rect 9781 765 9815 799
rect 10149 765 10183 799
rect 6699 697 6733 731
rect 13461 697 13495 731
rect 14105 765 14139 799
rect 14841 765 14875 799
rect 16405 765 16439 799
rect 17417 765 17451 799
rect 18521 765 18555 799
rect 2513 629 2547 663
rect 4721 629 4755 663
rect 9229 629 9263 663
rect 11621 629 11655 663
rect 13645 629 13679 663
rect 16267 629 16301 663
rect 1501 425 1535 459
rect 2605 425 2639 459
rect 3433 425 3467 459
rect 4905 425 4939 459
rect 6377 425 6411 459
rect 7297 425 7331 459
rect 7573 425 7607 459
rect 8493 425 8527 459
rect 10609 425 10643 459
rect 12725 425 12759 459
rect 15025 425 15059 459
rect 16957 425 16991 459
rect 17233 425 17267 459
rect 18521 425 18555 459
rect 13001 357 13035 391
rect 3249 289 3283 323
rect 5089 289 5123 323
rect 5181 289 5215 323
rect 6837 289 6871 323
rect 7021 289 7055 323
rect 9045 289 9079 323
rect 12449 289 12483 323
rect 14841 289 14875 323
rect 1317 221 1351 255
rect 3157 221 3191 255
rect 5549 221 5583 255
rect 8861 221 8895 255
rect 8953 221 8987 255
rect 10517 221 10551 255
rect 10701 221 10735 255
rect 10885 221 10919 255
rect 11161 221 11195 255
rect 12357 221 12391 255
rect 12817 221 12851 255
rect 13001 221 13035 255
rect 14749 221 14783 255
rect 16865 221 16899 255
rect 17049 221 17083 255
rect 17325 221 17359 255
rect 6745 153 6779 187
rect 10977 153 11011 187
rect 10885 85 10919 119
<< metal1 >>
rect 0 10906 18860 10928
rect 0 10854 4660 10906
rect 4712 10854 4724 10906
rect 4776 10854 4788 10906
rect 4840 10854 4852 10906
rect 4904 10854 4916 10906
rect 4968 10854 7760 10906
rect 7812 10854 7824 10906
rect 7876 10854 7888 10906
rect 7940 10854 7952 10906
rect 8004 10854 8016 10906
rect 8068 10854 10860 10906
rect 10912 10854 10924 10906
rect 10976 10854 10988 10906
rect 11040 10854 11052 10906
rect 11104 10854 11116 10906
rect 11168 10854 13960 10906
rect 14012 10854 14024 10906
rect 14076 10854 14088 10906
rect 14140 10854 14152 10906
rect 14204 10854 14216 10906
rect 14268 10854 17060 10906
rect 17112 10854 17124 10906
rect 17176 10854 17188 10906
rect 17240 10854 17252 10906
rect 17304 10854 17316 10906
rect 17368 10854 18860 10906
rect 0 10832 18860 10854
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 7285 10795 7343 10801
rect 7285 10792 7297 10795
rect 7156 10764 7297 10792
rect 7156 10752 7162 10764
rect 7285 10761 7297 10764
rect 7331 10761 7343 10795
rect 7285 10755 7343 10761
rect 8846 10752 8852 10804
rect 8904 10792 8910 10804
rect 8904 10764 9168 10792
rect 8904 10752 8910 10764
rect 9140 10733 9168 10764
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10045 10795 10103 10801
rect 10045 10792 10057 10795
rect 10008 10764 10057 10792
rect 10008 10752 10014 10764
rect 10045 10761 10057 10764
rect 10091 10761 10103 10795
rect 10045 10755 10103 10761
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 13909 10795 13967 10801
rect 13909 10792 13921 10795
rect 12860 10764 13921 10792
rect 12860 10752 12866 10764
rect 13909 10761 13921 10764
rect 13955 10761 13967 10795
rect 13909 10755 13967 10761
rect 18325 10795 18383 10801
rect 18325 10761 18337 10795
rect 18371 10761 18383 10795
rect 18325 10755 18383 10761
rect 8297 10727 8355 10733
rect 8297 10693 8309 10727
rect 8343 10724 8355 10727
rect 9033 10727 9091 10733
rect 9033 10724 9045 10727
rect 8343 10696 9045 10724
rect 8343 10693 8355 10696
rect 8297 10687 8355 10693
rect 9033 10693 9045 10696
rect 9079 10693 9091 10727
rect 9033 10687 9091 10693
rect 9125 10727 9183 10733
rect 9125 10693 9137 10727
rect 9171 10724 9183 10727
rect 10870 10724 10876 10736
rect 9171 10696 10876 10724
rect 9171 10693 9183 10696
rect 9125 10687 9183 10693
rect 10870 10684 10876 10696
rect 10928 10684 10934 10736
rect 12345 10727 12403 10733
rect 12345 10693 12357 10727
rect 12391 10724 12403 10727
rect 13078 10724 13084 10736
rect 12391 10696 13084 10724
rect 12391 10693 12403 10696
rect 12345 10687 12403 10693
rect 13078 10684 13084 10696
rect 13136 10684 13142 10736
rect 18141 10727 18199 10733
rect 18141 10724 18153 10727
rect 14108 10696 18153 10724
rect 1949 10659 2007 10665
rect 1949 10625 1961 10659
rect 1995 10625 2007 10659
rect 2130 10656 2136 10668
rect 2091 10628 2136 10656
rect 1949 10619 2007 10625
rect 1964 10588 1992 10619
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 3510 10616 3516 10668
rect 3568 10656 3574 10668
rect 3881 10659 3939 10665
rect 3881 10656 3893 10659
rect 3568 10628 3893 10656
rect 3568 10616 3574 10628
rect 3881 10625 3893 10628
rect 3927 10625 3939 10659
rect 3881 10619 3939 10625
rect 6086 10616 6092 10668
rect 6144 10656 6150 10668
rect 6273 10659 6331 10665
rect 6273 10656 6285 10659
rect 6144 10628 6285 10656
rect 6144 10616 6150 10628
rect 6273 10625 6285 10628
rect 6319 10625 6331 10659
rect 6273 10619 6331 10625
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10625 7527 10659
rect 7469 10619 7527 10625
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10625 7987 10659
rect 7929 10619 7987 10625
rect 8113 10659 8171 10665
rect 8113 10625 8125 10659
rect 8159 10656 8171 10659
rect 10229 10659 10287 10665
rect 8159 10628 10180 10656
rect 8159 10625 8171 10628
rect 8113 10619 8171 10625
rect 2038 10588 2044 10600
rect 1964 10560 2044 10588
rect 2038 10548 2044 10560
rect 2096 10548 2102 10600
rect 3786 10588 3792 10600
rect 3747 10560 3792 10588
rect 3786 10548 3792 10560
rect 3844 10548 3850 10600
rect 7484 10520 7512 10619
rect 7944 10588 7972 10619
rect 8938 10588 8944 10600
rect 7944 10560 8616 10588
rect 8899 10560 8944 10588
rect 8588 10529 8616 10560
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 10152 10588 10180 10628
rect 10229 10625 10241 10659
rect 10275 10656 10287 10659
rect 11882 10656 11888 10668
rect 10275 10628 11888 10656
rect 10275 10625 10287 10628
rect 10229 10619 10287 10625
rect 11882 10616 11888 10628
rect 11940 10616 11946 10668
rect 12437 10659 12495 10665
rect 12437 10625 12449 10659
rect 12483 10656 12495 10659
rect 12894 10656 12900 10668
rect 12483 10628 12900 10656
rect 12483 10625 12495 10628
rect 12437 10619 12495 10625
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 14108 10665 14136 10696
rect 18141 10693 18153 10696
rect 18187 10693 18199 10727
rect 18141 10687 18199 10693
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10625 13783 10659
rect 13725 10619 13783 10625
rect 14093 10659 14151 10665
rect 14093 10625 14105 10659
rect 14139 10625 14151 10659
rect 14093 10619 14151 10625
rect 15013 10659 15071 10665
rect 15013 10625 15025 10659
rect 15059 10625 15071 10659
rect 15013 10619 15071 10625
rect 11238 10588 11244 10600
rect 10152 10560 11244 10588
rect 11238 10548 11244 10560
rect 11296 10548 11302 10600
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10557 12311 10591
rect 12802 10588 12808 10600
rect 12253 10551 12311 10557
rect 12406 10560 12808 10588
rect 8573 10523 8631 10529
rect 7484 10492 8524 10520
rect 1946 10412 1952 10464
rect 2004 10452 2010 10464
rect 2041 10455 2099 10461
rect 2041 10452 2053 10455
rect 2004 10424 2053 10452
rect 2004 10412 2010 10424
rect 2041 10421 2053 10424
rect 2087 10421 2099 10455
rect 2041 10415 2099 10421
rect 4249 10455 4307 10461
rect 4249 10421 4261 10455
rect 4295 10452 4307 10455
rect 5258 10452 5264 10464
rect 4295 10424 5264 10452
rect 4295 10421 4307 10424
rect 4249 10415 4307 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 6273 10455 6331 10461
rect 6273 10452 6285 10455
rect 6052 10424 6285 10452
rect 6052 10412 6058 10424
rect 6273 10421 6285 10424
rect 6319 10421 6331 10455
rect 6273 10415 6331 10421
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 7745 10455 7803 10461
rect 7745 10452 7757 10455
rect 7708 10424 7757 10452
rect 7708 10412 7714 10424
rect 7745 10421 7757 10424
rect 7791 10421 7803 10455
rect 8496 10452 8524 10492
rect 8573 10489 8585 10523
rect 8619 10489 8631 10523
rect 12268 10520 12296 10551
rect 12406 10520 12434 10560
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 13740 10588 13768 10619
rect 15028 10588 15056 10619
rect 15102 10616 15108 10668
rect 15160 10656 15166 10668
rect 15657 10659 15715 10665
rect 15657 10656 15669 10659
rect 15160 10628 15669 10656
rect 15160 10616 15166 10628
rect 15657 10625 15669 10628
rect 15703 10625 15715 10659
rect 15657 10619 15715 10625
rect 16945 10659 17003 10665
rect 16945 10625 16957 10659
rect 16991 10625 17003 10659
rect 18046 10656 18052 10668
rect 18007 10628 18052 10656
rect 16945 10619 17003 10625
rect 16960 10588 16988 10619
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 18233 10659 18291 10665
rect 18233 10625 18245 10659
rect 18279 10656 18291 10659
rect 18340 10656 18368 10755
rect 18279 10628 18368 10656
rect 18509 10659 18567 10665
rect 18279 10625 18291 10628
rect 18233 10619 18291 10625
rect 18509 10625 18521 10659
rect 18555 10656 18567 10659
rect 18782 10656 18788 10668
rect 18555 10628 18788 10656
rect 18555 10625 18567 10628
rect 18509 10619 18567 10625
rect 13740 10560 16988 10588
rect 17865 10591 17923 10597
rect 13740 10520 13768 10560
rect 17865 10557 17877 10591
rect 17911 10588 17923 10591
rect 18524 10588 18552 10619
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 17911 10560 18552 10588
rect 17911 10557 17923 10560
rect 17865 10551 17923 10557
rect 12268 10492 12434 10520
rect 12820 10492 13768 10520
rect 8573 10483 8631 10489
rect 12820 10461 12848 10492
rect 12805 10455 12863 10461
rect 12805 10452 12817 10455
rect 8496 10424 12817 10452
rect 7745 10415 7803 10421
rect 12805 10421 12817 10424
rect 12851 10421 12863 10455
rect 12805 10415 12863 10421
rect 13262 10412 13268 10464
rect 13320 10452 13326 10464
rect 13449 10455 13507 10461
rect 13449 10452 13461 10455
rect 13320 10424 13461 10452
rect 13320 10412 13326 10424
rect 13449 10421 13461 10424
rect 13495 10421 13507 10455
rect 14458 10452 14464 10464
rect 14419 10424 14464 10452
rect 13449 10415 13507 10421
rect 14458 10412 14464 10424
rect 14516 10412 14522 10464
rect 14734 10412 14740 10464
rect 14792 10452 14798 10464
rect 14921 10455 14979 10461
rect 14921 10452 14933 10455
rect 14792 10424 14933 10452
rect 14792 10412 14798 10424
rect 14921 10421 14933 10424
rect 14967 10421 14979 10455
rect 14921 10415 14979 10421
rect 15194 10412 15200 10464
rect 15252 10452 15258 10464
rect 16301 10455 16359 10461
rect 16301 10452 16313 10455
rect 15252 10424 16313 10452
rect 15252 10412 15258 10424
rect 16301 10421 16313 10424
rect 16347 10421 16359 10455
rect 16942 10452 16948 10464
rect 16903 10424 16948 10452
rect 16301 10415 16359 10421
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 0 10362 18860 10384
rect 0 10310 3110 10362
rect 3162 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 3302 10362
rect 3354 10310 3366 10362
rect 3418 10310 6210 10362
rect 6262 10310 6274 10362
rect 6326 10310 6338 10362
rect 6390 10310 6402 10362
rect 6454 10310 6466 10362
rect 6518 10310 9310 10362
rect 9362 10310 9374 10362
rect 9426 10310 9438 10362
rect 9490 10310 9502 10362
rect 9554 10310 9566 10362
rect 9618 10310 12410 10362
rect 12462 10310 12474 10362
rect 12526 10310 12538 10362
rect 12590 10310 12602 10362
rect 12654 10310 12666 10362
rect 12718 10310 15510 10362
rect 15562 10310 15574 10362
rect 15626 10310 15638 10362
rect 15690 10310 15702 10362
rect 15754 10310 15766 10362
rect 15818 10310 18860 10362
rect 0 10288 18860 10310
rect 3421 10251 3479 10257
rect 3421 10217 3433 10251
rect 3467 10248 3479 10251
rect 3510 10248 3516 10260
rect 3467 10220 3516 10248
rect 3467 10217 3479 10220
rect 3421 10211 3479 10217
rect 3510 10208 3516 10220
rect 3568 10208 3574 10260
rect 3786 10208 3792 10260
rect 3844 10248 3850 10260
rect 3881 10251 3939 10257
rect 3881 10248 3893 10251
rect 3844 10220 3893 10248
rect 3844 10208 3850 10220
rect 3881 10217 3893 10220
rect 3927 10217 3939 10251
rect 3881 10211 3939 10217
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 7883 10251 7941 10257
rect 7883 10248 7895 10251
rect 6972 10220 7895 10248
rect 6972 10208 6978 10220
rect 7883 10217 7895 10220
rect 7929 10248 7941 10251
rect 12621 10251 12679 10257
rect 7929 10220 12434 10248
rect 7929 10217 7941 10220
rect 7883 10211 7941 10217
rect 8573 10183 8631 10189
rect 8573 10149 8585 10183
rect 8619 10180 8631 10183
rect 8846 10180 8852 10192
rect 8619 10152 8852 10180
rect 8619 10149 8631 10152
rect 8573 10143 8631 10149
rect 1673 10115 1731 10121
rect 1673 10112 1685 10115
rect 492 10084 1685 10112
rect 290 10004 296 10056
rect 348 10044 354 10056
rect 492 10053 520 10084
rect 1673 10081 1685 10084
rect 1719 10081 1731 10115
rect 1946 10112 1952 10124
rect 1907 10084 1952 10112
rect 1673 10075 1731 10081
rect 1946 10072 1952 10084
rect 2004 10072 2010 10124
rect 5994 10072 6000 10124
rect 6052 10112 6058 10124
rect 6089 10115 6147 10121
rect 6089 10112 6101 10115
rect 6052 10084 6101 10112
rect 6052 10072 6058 10084
rect 6089 10081 6101 10084
rect 6135 10081 6147 10115
rect 6089 10075 6147 10081
rect 477 10047 535 10053
rect 477 10044 489 10047
rect 348 10016 489 10044
rect 348 10004 354 10016
rect 477 10013 489 10016
rect 523 10013 535 10047
rect 934 10044 940 10056
rect 895 10016 940 10044
rect 477 10007 535 10013
rect 934 10004 940 10016
rect 992 10004 998 10056
rect 1121 10047 1179 10053
rect 1121 10013 1133 10047
rect 1167 10013 1179 10047
rect 1121 10007 1179 10013
rect 382 9976 388 9988
rect 343 9948 388 9976
rect 382 9936 388 9948
rect 440 9936 446 9988
rect 1136 9976 1164 10007
rect 1210 10004 1216 10056
rect 1268 10044 1274 10056
rect 1305 10047 1363 10053
rect 1305 10044 1317 10047
rect 1268 10016 1317 10044
rect 1268 10004 1274 10016
rect 1305 10013 1317 10016
rect 1351 10013 1363 10047
rect 3694 10044 3700 10056
rect 3655 10016 3700 10044
rect 1305 10007 1363 10013
rect 3694 10004 3700 10016
rect 3752 10004 3758 10056
rect 3878 10044 3884 10056
rect 3839 10016 3884 10044
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 6454 10044 6460 10056
rect 6415 10016 6460 10044
rect 6454 10004 6460 10016
rect 6512 10004 6518 10056
rect 8588 10044 8616 10143
rect 8846 10140 8852 10152
rect 8904 10140 8910 10192
rect 12406 10180 12434 10220
rect 12621 10217 12633 10251
rect 12667 10248 12679 10251
rect 12802 10248 12808 10260
rect 12667 10220 12808 10248
rect 12667 10217 12679 10220
rect 12621 10211 12679 10217
rect 12802 10208 12808 10220
rect 12860 10208 12866 10260
rect 13814 10248 13820 10260
rect 13096 10220 13820 10248
rect 13096 10180 13124 10220
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 15102 10257 15108 10260
rect 15059 10251 15108 10257
rect 15059 10217 15071 10251
rect 15105 10217 15108 10251
rect 15059 10211 15108 10217
rect 15102 10208 15108 10211
rect 15160 10208 15166 10260
rect 17819 10251 17877 10257
rect 17819 10217 17831 10251
rect 17865 10248 17877 10251
rect 18046 10248 18052 10260
rect 17865 10220 18052 10248
rect 17865 10217 17877 10220
rect 17819 10211 17877 10217
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 12406 10152 13124 10180
rect 8941 10115 8999 10121
rect 8941 10081 8953 10115
rect 8987 10112 8999 10115
rect 9214 10112 9220 10124
rect 8987 10084 9220 10112
rect 8987 10081 8999 10084
rect 8941 10075 8999 10081
rect 9214 10072 9220 10084
rect 9272 10112 9278 10124
rect 10873 10115 10931 10121
rect 10873 10112 10885 10115
rect 9272 10084 10885 10112
rect 9272 10072 9278 10084
rect 10873 10081 10885 10084
rect 10919 10081 10931 10115
rect 10873 10075 10931 10081
rect 11149 10115 11207 10121
rect 11149 10081 11161 10115
rect 11195 10112 11207 10115
rect 11514 10112 11520 10124
rect 11195 10084 11520 10112
rect 11195 10081 11207 10084
rect 11149 10075 11207 10081
rect 11514 10072 11520 10084
rect 11572 10072 11578 10124
rect 13262 10112 13268 10124
rect 13223 10084 13268 10112
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 13633 10115 13691 10121
rect 13633 10081 13645 10115
rect 13679 10112 13691 10115
rect 14458 10112 14464 10124
rect 13679 10084 14464 10112
rect 13679 10081 13691 10084
rect 13633 10075 13691 10081
rect 14458 10072 14464 10084
rect 14516 10072 14522 10124
rect 16025 10115 16083 10121
rect 16025 10081 16037 10115
rect 16071 10112 16083 10115
rect 16942 10112 16948 10124
rect 16071 10084 16948 10112
rect 16071 10081 16083 10084
rect 16025 10075 16083 10081
rect 16942 10072 16948 10084
rect 17000 10072 17006 10124
rect 7484 10016 8616 10044
rect 16393 10047 16451 10053
rect 7484 9988 7512 10016
rect 16393 10013 16405 10047
rect 16439 10044 16451 10047
rect 16482 10044 16488 10056
rect 16439 10016 16488 10044
rect 16439 10013 16451 10016
rect 16393 10007 16451 10013
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 18233 10047 18291 10053
rect 18233 10013 18245 10047
rect 18279 10044 18291 10047
rect 18509 10047 18567 10053
rect 18509 10044 18521 10047
rect 18279 10016 18521 10044
rect 18279 10013 18291 10016
rect 18233 10007 18291 10013
rect 18509 10013 18521 10016
rect 18555 10044 18567 10047
rect 18598 10044 18604 10056
rect 18555 10016 18604 10044
rect 18555 10013 18567 10016
rect 18509 10007 18567 10013
rect 18598 10004 18604 10016
rect 18656 10004 18662 10056
rect 1397 9979 1455 9985
rect 1136 9948 1348 9976
rect 658 9868 664 9920
rect 716 9908 722 9920
rect 1320 9917 1348 9948
rect 1397 9945 1409 9979
rect 1443 9945 1455 9979
rect 1578 9976 1584 9988
rect 1539 9948 1584 9976
rect 1397 9939 1455 9945
rect 937 9911 995 9917
rect 937 9908 949 9911
rect 716 9880 949 9908
rect 716 9868 722 9880
rect 937 9877 949 9880
rect 983 9877 995 9911
rect 937 9871 995 9877
rect 1305 9911 1363 9917
rect 1305 9877 1317 9911
rect 1351 9877 1363 9911
rect 1412 9908 1440 9939
rect 1578 9936 1584 9948
rect 1636 9936 1642 9988
rect 2590 9908 2596 9920
rect 1412 9880 2596 9908
rect 1305 9871 1363 9877
rect 2590 9868 2596 9880
rect 2648 9868 2654 9920
rect 3160 9908 3188 9962
rect 7466 9936 7472 9988
rect 7524 9936 7530 9988
rect 9217 9979 9275 9985
rect 9217 9945 9229 9979
rect 9263 9945 9275 9979
rect 10870 9976 10876 9988
rect 10442 9948 10876 9976
rect 9217 9939 9275 9945
rect 3602 9908 3608 9920
rect 3160 9880 3608 9908
rect 3602 9868 3608 9880
rect 3660 9908 3666 9920
rect 4065 9911 4123 9917
rect 4065 9908 4077 9911
rect 3660 9880 4077 9908
rect 3660 9868 3666 9880
rect 4065 9877 4077 9880
rect 4111 9908 4123 9911
rect 5905 9911 5963 9917
rect 5905 9908 5917 9911
rect 4111 9880 5917 9908
rect 4111 9877 4123 9880
rect 4065 9871 4123 9877
rect 5905 9877 5917 9880
rect 5951 9908 5963 9911
rect 7484 9908 7512 9936
rect 5951 9880 7512 9908
rect 9232 9908 9260 9939
rect 10226 9908 10232 9920
rect 9232 9880 10232 9908
rect 5951 9877 5963 9880
rect 5905 9871 5963 9877
rect 10226 9868 10232 9880
rect 10284 9868 10290 9920
rect 10686 9908 10692 9920
rect 10647 9880 10692 9908
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 10796 9908 10824 9948
rect 10870 9936 10876 9948
rect 10928 9936 10934 9988
rect 12360 9908 12388 9962
rect 12434 9908 12440 9920
rect 10796 9880 12440 9908
rect 12434 9868 12440 9880
rect 12492 9908 12498 9920
rect 13081 9911 13139 9917
rect 13081 9908 13093 9911
rect 12492 9880 13093 9908
rect 12492 9868 12498 9880
rect 13081 9877 13093 9880
rect 13127 9908 13139 9911
rect 14660 9908 14688 9962
rect 15933 9911 15991 9917
rect 15933 9908 15945 9911
rect 13127 9880 15945 9908
rect 13127 9877 13139 9880
rect 13081 9871 13139 9877
rect 15933 9877 15945 9880
rect 15979 9908 15991 9911
rect 16114 9908 16120 9920
rect 15979 9880 16120 9908
rect 15979 9877 15991 9880
rect 15933 9871 15991 9877
rect 16114 9868 16120 9880
rect 16172 9908 16178 9920
rect 16776 9908 16804 9962
rect 18322 9908 18328 9920
rect 16172 9880 16804 9908
rect 18283 9880 18328 9908
rect 16172 9868 16178 9880
rect 18322 9868 18328 9880
rect 18380 9868 18386 9920
rect 0 9818 18860 9840
rect 0 9766 4660 9818
rect 4712 9766 4724 9818
rect 4776 9766 4788 9818
rect 4840 9766 4852 9818
rect 4904 9766 4916 9818
rect 4968 9766 7760 9818
rect 7812 9766 7824 9818
rect 7876 9766 7888 9818
rect 7940 9766 7952 9818
rect 8004 9766 8016 9818
rect 8068 9766 10860 9818
rect 10912 9766 10924 9818
rect 10976 9766 10988 9818
rect 11040 9766 11052 9818
rect 11104 9766 11116 9818
rect 11168 9766 13960 9818
rect 14012 9766 14024 9818
rect 14076 9766 14088 9818
rect 14140 9766 14152 9818
rect 14204 9766 14216 9818
rect 14268 9766 17060 9818
rect 17112 9766 17124 9818
rect 17176 9766 17188 9818
rect 17240 9766 17252 9818
rect 17304 9766 17316 9818
rect 17368 9766 18860 9818
rect 0 9744 18860 9766
rect 2130 9664 2136 9716
rect 2188 9704 2194 9716
rect 2501 9707 2559 9713
rect 2501 9704 2513 9707
rect 2188 9676 2513 9704
rect 2188 9664 2194 9676
rect 2501 9673 2513 9676
rect 2547 9673 2559 9707
rect 2501 9667 2559 9673
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 3145 9707 3203 9713
rect 3145 9704 3157 9707
rect 3016 9676 3157 9704
rect 3016 9664 3022 9676
rect 3145 9673 3157 9676
rect 3191 9673 3203 9707
rect 5258 9704 5264 9716
rect 5219 9676 5264 9704
rect 3145 9667 3203 9673
rect 5258 9664 5264 9676
rect 5316 9664 5322 9716
rect 5997 9707 6055 9713
rect 5997 9673 6009 9707
rect 6043 9673 6055 9707
rect 6454 9704 6460 9716
rect 6415 9676 6460 9704
rect 5997 9667 6055 9673
rect 2222 9636 2228 9648
rect 1702 9608 2228 9636
rect 2222 9596 2228 9608
rect 2280 9596 2286 9648
rect 2682 9636 2688 9648
rect 2424 9608 2688 9636
rect 293 9571 351 9577
rect 293 9537 305 9571
rect 339 9568 351 9571
rect 382 9568 388 9580
rect 339 9540 388 9568
rect 339 9537 351 9540
rect 293 9531 351 9537
rect 382 9528 388 9540
rect 440 9528 446 9580
rect 658 9568 664 9580
rect 619 9540 664 9568
rect 658 9528 664 9540
rect 716 9528 722 9580
rect 1578 9528 1584 9580
rect 1636 9568 1642 9580
rect 2087 9571 2145 9577
rect 2087 9568 2099 9571
rect 1636 9540 2099 9568
rect 1636 9528 1642 9540
rect 2087 9537 2099 9540
rect 2133 9568 2145 9571
rect 2424 9568 2452 9608
rect 2682 9596 2688 9608
rect 2740 9636 2746 9648
rect 3694 9636 3700 9648
rect 2740 9608 3096 9636
rect 2740 9596 2746 9608
rect 2133 9540 2452 9568
rect 2501 9571 2559 9577
rect 2133 9537 2145 9540
rect 2087 9531 2145 9537
rect 2501 9537 2513 9571
rect 2547 9537 2559 9571
rect 2501 9531 2559 9537
rect 1210 9460 1216 9512
rect 1268 9500 1274 9512
rect 2516 9500 2544 9531
rect 2590 9528 2596 9580
rect 2648 9568 2654 9580
rect 2777 9571 2835 9577
rect 2648 9540 2693 9568
rect 2648 9528 2654 9540
rect 2777 9537 2789 9571
rect 2823 9537 2835 9571
rect 2777 9531 2835 9537
rect 1268 9472 2544 9500
rect 2792 9500 2820 9531
rect 2866 9528 2872 9580
rect 2924 9568 2930 9580
rect 3068 9568 3096 9608
rect 3252 9608 3700 9636
rect 3252 9577 3280 9608
rect 3694 9596 3700 9608
rect 3752 9636 3758 9648
rect 3881 9639 3939 9645
rect 3752 9608 3832 9636
rect 3752 9596 3758 9608
rect 3237 9571 3295 9577
rect 3237 9568 3249 9571
rect 2924 9540 2969 9568
rect 3068 9540 3249 9568
rect 2924 9528 2930 9540
rect 3237 9537 3249 9540
rect 3283 9537 3295 9571
rect 3237 9531 3295 9537
rect 3510 9528 3516 9580
rect 3568 9568 3574 9580
rect 3804 9577 3832 9608
rect 3881 9605 3893 9639
rect 3927 9636 3939 9639
rect 5353 9639 5411 9645
rect 3927 9608 4292 9636
rect 3927 9605 3939 9608
rect 3881 9599 3939 9605
rect 4264 9577 4292 9608
rect 5353 9605 5365 9639
rect 5399 9636 5411 9639
rect 5626 9636 5632 9648
rect 5399 9608 5632 9636
rect 5399 9605 5411 9608
rect 5353 9599 5411 9605
rect 5626 9596 5632 9608
rect 5684 9596 5690 9648
rect 6012 9636 6040 9667
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 11238 9704 11244 9716
rect 8220 9676 9168 9704
rect 11199 9676 11244 9704
rect 6365 9639 6423 9645
rect 6365 9636 6377 9639
rect 6012 9608 6377 9636
rect 6365 9605 6377 9608
rect 6411 9605 6423 9639
rect 6365 9599 6423 9605
rect 6549 9639 6607 9645
rect 6549 9605 6561 9639
rect 6595 9636 6607 9639
rect 6638 9636 6644 9648
rect 6595 9608 6644 9636
rect 6595 9605 6607 9608
rect 6549 9599 6607 9605
rect 6638 9596 6644 9608
rect 6696 9636 6702 9648
rect 8220 9636 8248 9676
rect 6696 9608 8248 9636
rect 6696 9596 6702 9608
rect 8846 9596 8852 9648
rect 8904 9596 8910 9648
rect 9140 9636 9168 9676
rect 11238 9664 11244 9676
rect 11296 9664 11302 9716
rect 11885 9707 11943 9713
rect 11885 9673 11897 9707
rect 11931 9704 11943 9707
rect 12434 9704 12440 9716
rect 11931 9676 12440 9704
rect 11931 9673 11943 9676
rect 11885 9667 11943 9673
rect 12434 9664 12440 9676
rect 12492 9664 12498 9716
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 16632 9676 17540 9704
rect 16632 9664 16638 9676
rect 9858 9636 9864 9648
rect 9140 9608 9864 9636
rect 9858 9596 9864 9608
rect 9916 9596 9922 9648
rect 11256 9636 11284 9664
rect 12253 9639 12311 9645
rect 12253 9636 12265 9639
rect 11256 9608 12265 9636
rect 12253 9605 12265 9608
rect 12299 9605 12311 9639
rect 14461 9639 14519 9645
rect 14461 9636 14473 9639
rect 14030 9608 14473 9636
rect 12253 9599 12311 9605
rect 14461 9605 14473 9608
rect 14507 9605 14519 9639
rect 14461 9599 14519 9605
rect 16114 9596 16120 9648
rect 16172 9596 16178 9648
rect 17512 9645 17540 9676
rect 17497 9639 17555 9645
rect 17497 9605 17509 9639
rect 17543 9605 17555 9639
rect 17497 9599 17555 9605
rect 3605 9571 3663 9577
rect 3605 9568 3617 9571
rect 3568 9540 3617 9568
rect 3568 9528 3574 9540
rect 3605 9537 3617 9540
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 3973 9571 4031 9577
rect 3973 9537 3985 9571
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 4249 9571 4307 9577
rect 4249 9537 4261 9571
rect 4295 9537 4307 9571
rect 5721 9571 5779 9577
rect 5721 9568 5733 9571
rect 4249 9531 4307 9537
rect 5000 9540 5733 9568
rect 3620 9500 3648 9531
rect 3988 9500 4016 9531
rect 2792 9472 4016 9500
rect 1268 9460 1274 9472
rect 2516 9432 2544 9472
rect 2516 9404 2774 9432
rect 2222 9364 2228 9376
rect 2183 9336 2228 9364
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 2746 9364 2774 9404
rect 2866 9392 2872 9444
rect 2924 9432 2930 9444
rect 3878 9432 3884 9444
rect 2924 9404 3884 9432
rect 2924 9392 2930 9404
rect 3878 9392 3884 9404
rect 3936 9432 3942 9444
rect 4080 9432 4108 9531
rect 4157 9503 4215 9509
rect 4157 9469 4169 9503
rect 4203 9500 4215 9503
rect 5000 9500 5028 9540
rect 5721 9537 5733 9540
rect 5767 9537 5779 9571
rect 5721 9531 5779 9537
rect 5905 9571 5963 9577
rect 5905 9537 5917 9571
rect 5951 9537 5963 9571
rect 5905 9531 5963 9537
rect 4203 9472 5028 9500
rect 4203 9469 4215 9472
rect 4157 9463 4215 9469
rect 5442 9460 5448 9512
rect 5500 9500 5506 9512
rect 5500 9472 5545 9500
rect 5500 9460 5506 9472
rect 5166 9432 5172 9444
rect 3936 9404 4108 9432
rect 4724 9404 5172 9432
rect 3936 9392 3942 9404
rect 3970 9364 3976 9376
rect 2746 9336 3976 9364
rect 3970 9324 3976 9336
rect 4028 9364 4034 9376
rect 4724 9364 4752 9404
rect 5166 9392 5172 9404
rect 5224 9432 5230 9444
rect 5920 9432 5948 9531
rect 5994 9528 6000 9580
rect 6052 9568 6058 9580
rect 6273 9571 6331 9577
rect 6273 9568 6285 9571
rect 6052 9540 6285 9568
rect 6052 9528 6058 9540
rect 6273 9537 6285 9540
rect 6319 9537 6331 9571
rect 6273 9531 6331 9537
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9568 6883 9571
rect 6914 9568 6920 9580
rect 6871 9540 6920 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7466 9568 7472 9580
rect 7427 9540 7472 9568
rect 7466 9528 7472 9540
rect 7524 9528 7530 9580
rect 9766 9528 9772 9580
rect 9824 9568 9830 9580
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 9824 9540 9965 9568
rect 9824 9528 9830 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 14734 9568 14740 9580
rect 14695 9540 14740 9568
rect 9953 9531 10011 9537
rect 14734 9528 14740 9540
rect 14792 9528 14798 9580
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9568 15163 9571
rect 15194 9568 15200 9580
rect 15151 9540 15200 9568
rect 15151 9537 15163 9540
rect 15105 9531 15163 9537
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 16531 9571 16589 9577
rect 16531 9537 16543 9571
rect 16577 9568 16589 9571
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16577 9540 16865 9568
rect 16577 9537 16589 9540
rect 16531 9531 16589 9537
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 6086 9460 6092 9512
rect 6144 9500 6150 9512
rect 7561 9503 7619 9509
rect 7561 9500 7573 9503
rect 6144 9472 7573 9500
rect 6144 9460 6150 9472
rect 7561 9469 7573 9472
rect 7607 9469 7619 9503
rect 7561 9463 7619 9469
rect 7837 9503 7895 9509
rect 7837 9469 7849 9503
rect 7883 9500 7895 9503
rect 8478 9500 8484 9512
rect 7883 9472 8484 9500
rect 7883 9469 7895 9472
rect 7837 9463 7895 9469
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 9030 9460 9036 9512
rect 9088 9500 9094 9512
rect 9088 9472 9996 9500
rect 9088 9460 9094 9472
rect 5224 9404 5948 9432
rect 5224 9392 5230 9404
rect 8846 9392 8852 9444
rect 8904 9432 8910 9444
rect 9309 9435 9367 9441
rect 9309 9432 9321 9435
rect 8904 9404 9321 9432
rect 8904 9392 8910 9404
rect 9309 9401 9321 9404
rect 9355 9432 9367 9435
rect 9858 9432 9864 9444
rect 9355 9404 9864 9432
rect 9355 9401 9367 9404
rect 9309 9395 9367 9401
rect 9858 9392 9864 9404
rect 9916 9392 9922 9444
rect 9968 9432 9996 9472
rect 12250 9460 12256 9512
rect 12308 9500 12314 9512
rect 12529 9503 12587 9509
rect 12529 9500 12541 9503
rect 12308 9472 12541 9500
rect 12308 9460 12314 9472
rect 12529 9469 12541 9472
rect 12575 9469 12587 9503
rect 12529 9463 12587 9469
rect 12805 9503 12863 9509
rect 12805 9469 12817 9503
rect 12851 9500 12863 9503
rect 18322 9500 18328 9512
rect 12851 9472 18328 9500
rect 12851 9469 12863 9472
rect 12805 9463 12863 9469
rect 18322 9460 18328 9472
rect 18380 9460 18386 9512
rect 14277 9435 14335 9441
rect 9968 9404 12434 9432
rect 4890 9364 4896 9376
rect 4028 9336 4752 9364
rect 4851 9336 4896 9364
rect 4028 9324 4034 9336
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 5592 9336 6193 9364
rect 5592 9324 5598 9336
rect 6181 9333 6193 9336
rect 6227 9364 6239 9367
rect 6733 9367 6791 9373
rect 6733 9364 6745 9367
rect 6227 9336 6745 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 6733 9333 6745 9336
rect 6779 9333 6791 9367
rect 6733 9327 6791 9333
rect 7466 9324 7472 9376
rect 7524 9364 7530 9376
rect 9030 9364 9036 9376
rect 7524 9336 9036 9364
rect 7524 9324 7530 9336
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 9766 9364 9772 9376
rect 9727 9336 9772 9364
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 11330 9364 11336 9376
rect 10008 9336 11336 9364
rect 10008 9324 10014 9336
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 12158 9364 12164 9376
rect 12119 9336 12164 9364
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 12406 9364 12434 9404
rect 14277 9401 14289 9435
rect 14323 9432 14335 9435
rect 14734 9432 14740 9444
rect 14323 9404 14740 9432
rect 14323 9401 14335 9404
rect 14277 9395 14335 9401
rect 14734 9392 14740 9404
rect 14792 9392 14798 9444
rect 12986 9364 12992 9376
rect 12406 9336 12992 9364
rect 12986 9324 12992 9336
rect 13044 9324 13050 9376
rect 14461 9367 14519 9373
rect 14461 9333 14473 9367
rect 14507 9364 14519 9367
rect 14645 9367 14703 9373
rect 14645 9364 14657 9367
rect 14507 9336 14657 9364
rect 14507 9333 14519 9336
rect 14461 9327 14519 9333
rect 14645 9333 14657 9336
rect 14691 9364 14703 9367
rect 15286 9364 15292 9376
rect 14691 9336 15292 9364
rect 14691 9333 14703 9336
rect 14645 9327 14703 9333
rect 15286 9324 15292 9336
rect 15344 9364 15350 9376
rect 16114 9364 16120 9376
rect 15344 9336 16120 9364
rect 15344 9324 15350 9336
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 0 9274 18860 9296
rect 0 9222 3110 9274
rect 3162 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 3302 9274
rect 3354 9222 3366 9274
rect 3418 9222 6210 9274
rect 6262 9222 6274 9274
rect 6326 9222 6338 9274
rect 6390 9222 6402 9274
rect 6454 9222 6466 9274
rect 6518 9222 9310 9274
rect 9362 9222 9374 9274
rect 9426 9222 9438 9274
rect 9490 9222 9502 9274
rect 9554 9222 9566 9274
rect 9618 9222 12410 9274
rect 12462 9222 12474 9274
rect 12526 9222 12538 9274
rect 12590 9222 12602 9274
rect 12654 9222 12666 9274
rect 12718 9222 15510 9274
rect 15562 9222 15574 9274
rect 15626 9222 15638 9274
rect 15690 9222 15702 9274
rect 15754 9222 15766 9274
rect 15818 9222 18860 9274
rect 0 9200 18860 9222
rect 934 9120 940 9172
rect 992 9160 998 9172
rect 1029 9163 1087 9169
rect 1029 9160 1041 9163
rect 992 9132 1041 9160
rect 992 9120 998 9132
rect 1029 9129 1041 9132
rect 1075 9129 1087 9163
rect 1394 9160 1400 9172
rect 1355 9132 1400 9160
rect 1029 9123 1087 9129
rect 1394 9120 1400 9132
rect 1452 9120 1458 9172
rect 5629 9163 5687 9169
rect 5629 9129 5641 9163
rect 5675 9160 5687 9163
rect 5994 9160 6000 9172
rect 5675 9132 6000 9160
rect 5675 9129 5687 9132
rect 5629 9123 5687 9129
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 8478 9160 8484 9172
rect 8439 9132 8484 9160
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 11882 9160 11888 9172
rect 8588 9132 11284 9160
rect 11843 9132 11888 9160
rect 2590 9052 2596 9104
rect 2648 9092 2654 9104
rect 6638 9092 6644 9104
rect 2648 9064 6644 9092
rect 2648 9052 2654 9064
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 7190 9052 7196 9104
rect 7248 9092 7254 9104
rect 8588 9092 8616 9132
rect 7248 9064 8616 9092
rect 9677 9095 9735 9101
rect 7248 9052 7254 9064
rect 9677 9061 9689 9095
rect 9723 9061 9735 9095
rect 10502 9092 10508 9104
rect 10463 9064 10508 9092
rect 9677 9055 9735 9061
rect 2130 9024 2136 9036
rect 1136 8996 2136 9024
rect 1136 8965 1164 8996
rect 2130 8984 2136 8996
rect 2188 8984 2194 9036
rect 3694 8984 3700 9036
rect 3752 9024 3758 9036
rect 4341 9027 4399 9033
rect 4341 9024 4353 9027
rect 3752 8996 4353 9024
rect 3752 8984 3758 8996
rect 4341 8993 4353 8996
rect 4387 8993 4399 9027
rect 8846 9024 8852 9036
rect 4341 8987 4399 8993
rect 6656 8996 8852 9024
rect 937 8959 995 8965
rect 937 8925 949 8959
rect 983 8925 995 8959
rect 937 8919 995 8925
rect 1121 8959 1179 8965
rect 1121 8925 1133 8959
rect 1167 8925 1179 8959
rect 1121 8919 1179 8925
rect 952 8888 980 8919
rect 1394 8916 1400 8968
rect 1452 8956 1458 8968
rect 1489 8959 1547 8965
rect 1489 8956 1501 8959
rect 1452 8928 1501 8956
rect 1452 8916 1458 8928
rect 1489 8925 1501 8928
rect 1535 8925 1547 8959
rect 1489 8919 1547 8925
rect 2222 8916 2228 8968
rect 2280 8956 2286 8968
rect 2685 8959 2743 8965
rect 2685 8956 2697 8959
rect 2280 8928 2697 8956
rect 2280 8916 2286 8928
rect 2685 8925 2697 8928
rect 2731 8956 2743 8959
rect 2961 8959 3019 8965
rect 2961 8956 2973 8959
rect 2731 8928 2973 8956
rect 2731 8925 2743 8928
rect 2685 8919 2743 8925
rect 2961 8925 2973 8928
rect 3007 8956 3019 8959
rect 3602 8956 3608 8968
rect 3007 8928 3608 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 3602 8916 3608 8928
rect 3660 8916 3666 8968
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4890 8956 4896 8968
rect 4203 8928 4896 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 4890 8916 4896 8928
rect 4948 8916 4954 8968
rect 5534 8956 5540 8968
rect 5495 8928 5540 8956
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 5626 8916 5632 8968
rect 5684 8956 5690 8968
rect 6656 8965 6684 8996
rect 8846 8984 8852 8996
rect 8904 8984 8910 9036
rect 9692 9024 9720 9055
rect 10502 9052 10508 9064
rect 10560 9052 10566 9104
rect 10873 9095 10931 9101
rect 10873 9061 10885 9095
rect 10919 9061 10931 9095
rect 10873 9055 10931 9061
rect 10318 9024 10324 9036
rect 9140 8996 9720 9024
rect 10279 8996 10324 9024
rect 6641 8959 6699 8965
rect 5684 8928 5729 8956
rect 5684 8916 5690 8928
rect 6641 8925 6653 8959
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 6825 8959 6883 8965
rect 6825 8925 6837 8959
rect 6871 8956 6883 8959
rect 7282 8956 7288 8968
rect 6871 8928 7288 8956
rect 6871 8925 6883 8928
rect 6825 8919 6883 8925
rect 7282 8916 7288 8928
rect 7340 8956 7346 8968
rect 7466 8956 7472 8968
rect 7340 8928 7472 8956
rect 7340 8916 7346 8928
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 7837 8959 7895 8965
rect 7837 8925 7849 8959
rect 7883 8956 7895 8959
rect 8110 8956 8116 8968
rect 7883 8928 8116 8956
rect 7883 8925 7895 8928
rect 7837 8919 7895 8925
rect 2314 8888 2320 8900
rect 952 8860 2320 8888
rect 2314 8848 2320 8860
rect 2372 8848 2378 8900
rect 2774 8888 2780 8900
rect 2516 8860 2780 8888
rect 2130 8780 2136 8832
rect 2188 8820 2194 8832
rect 2516 8820 2544 8860
rect 2774 8848 2780 8860
rect 2832 8848 2838 8900
rect 2884 8860 3832 8888
rect 2188 8792 2544 8820
rect 2188 8780 2194 8792
rect 2590 8780 2596 8832
rect 2648 8820 2654 8832
rect 2884 8820 2912 8860
rect 3804 8829 3832 8860
rect 4062 8848 4068 8900
rect 4120 8888 4126 8900
rect 5353 8891 5411 8897
rect 5353 8888 5365 8891
rect 4120 8860 5365 8888
rect 4120 8848 4126 8860
rect 5353 8857 5365 8860
rect 5399 8888 5411 8891
rect 5442 8888 5448 8900
rect 5399 8860 5448 8888
rect 5399 8857 5411 8860
rect 5353 8851 5411 8857
rect 5442 8848 5448 8860
rect 5500 8848 5506 8900
rect 6086 8848 6092 8900
rect 6144 8888 6150 8900
rect 6457 8891 6515 8897
rect 6457 8888 6469 8891
rect 6144 8860 6469 8888
rect 6144 8848 6150 8860
rect 6457 8857 6469 8860
rect 6503 8857 6515 8891
rect 6457 8851 6515 8857
rect 6546 8848 6552 8900
rect 6604 8888 6610 8900
rect 6917 8891 6975 8897
rect 6917 8888 6929 8891
rect 6604 8860 6929 8888
rect 6604 8848 6610 8860
rect 6917 8857 6929 8860
rect 6963 8857 6975 8891
rect 7098 8888 7104 8900
rect 7059 8860 7104 8888
rect 6917 8851 6975 8857
rect 7098 8848 7104 8860
rect 7156 8848 7162 8900
rect 7760 8888 7788 8919
rect 8110 8916 8116 8928
rect 8168 8956 8174 8968
rect 8665 8959 8723 8965
rect 8665 8956 8677 8959
rect 8168 8928 8677 8956
rect 8168 8916 8174 8928
rect 8665 8925 8677 8928
rect 8711 8925 8723 8959
rect 8665 8919 8723 8925
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 9140 8956 9168 8996
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 10888 9024 10916 9055
rect 10612 8996 10916 9024
rect 8803 8928 9168 8956
rect 9217 8959 9275 8965
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 9217 8925 9229 8959
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 8478 8888 8484 8900
rect 7760 8860 8484 8888
rect 8478 8848 8484 8860
rect 8536 8848 8542 8900
rect 9030 8848 9036 8900
rect 9088 8888 9094 8900
rect 9232 8888 9260 8919
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 10505 8959 10563 8965
rect 10505 8956 10517 8959
rect 9456 8928 10517 8956
rect 9456 8916 9462 8928
rect 10505 8925 10517 8928
rect 10551 8925 10563 8959
rect 10505 8919 10563 8925
rect 9088 8860 9260 8888
rect 9309 8891 9367 8897
rect 9088 8848 9094 8860
rect 9309 8857 9321 8891
rect 9355 8857 9367 8891
rect 9309 8851 9367 8857
rect 9493 8891 9551 8897
rect 9493 8857 9505 8891
rect 9539 8888 9551 8891
rect 9858 8888 9864 8900
rect 9539 8860 9864 8888
rect 9539 8857 9551 8860
rect 9493 8851 9551 8857
rect 2648 8792 2912 8820
rect 3789 8823 3847 8829
rect 2648 8780 2654 8792
rect 3789 8789 3801 8823
rect 3835 8789 3847 8823
rect 3789 8783 3847 8789
rect 4249 8823 4307 8829
rect 4249 8789 4261 8823
rect 4295 8820 4307 8823
rect 5718 8820 5724 8832
rect 4295 8792 5724 8820
rect 4295 8789 4307 8792
rect 4249 8783 4307 8789
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 7009 8823 7067 8829
rect 7009 8789 7021 8823
rect 7055 8820 7067 8823
rect 7377 8823 7435 8829
rect 7377 8820 7389 8823
rect 7055 8792 7389 8820
rect 7055 8789 7067 8792
rect 7009 8783 7067 8789
rect 7377 8789 7389 8792
rect 7423 8789 7435 8823
rect 7377 8783 7435 8789
rect 7558 8780 7564 8832
rect 7616 8820 7622 8832
rect 8021 8823 8079 8829
rect 8021 8820 8033 8823
rect 7616 8792 8033 8820
rect 7616 8780 7622 8792
rect 8021 8789 8033 8792
rect 8067 8789 8079 8823
rect 8021 8783 8079 8789
rect 9125 8823 9183 8829
rect 9125 8789 9137 8823
rect 9171 8820 9183 8823
rect 9217 8823 9275 8829
rect 9217 8820 9229 8823
rect 9171 8792 9229 8820
rect 9171 8789 9183 8792
rect 9125 8783 9183 8789
rect 9217 8789 9229 8792
rect 9263 8789 9275 8823
rect 9324 8820 9352 8851
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 10045 8891 10103 8897
rect 10045 8857 10057 8891
rect 10091 8888 10103 8891
rect 10612 8888 10640 8996
rect 10689 8959 10747 8965
rect 10689 8925 10701 8959
rect 10735 8956 10747 8959
rect 10778 8956 10784 8968
rect 10735 8928 10784 8956
rect 10735 8925 10747 8928
rect 10689 8919 10747 8925
rect 10778 8916 10784 8928
rect 10836 8916 10842 8968
rect 11256 8965 11284 9132
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 12066 9120 12072 9172
rect 12124 9160 12130 9172
rect 15473 9163 15531 9169
rect 12124 9132 14596 9160
rect 12124 9120 12130 9132
rect 12434 9092 12440 9104
rect 12268 9064 12440 9092
rect 11422 9024 11428 9036
rect 11383 8996 11428 9024
rect 11422 8984 11428 8996
rect 11480 8984 11486 9036
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 11330 8916 11336 8968
rect 11388 8956 11394 8968
rect 12268 8965 12296 9064
rect 12434 9052 12440 9064
rect 12492 9092 12498 9104
rect 12894 9092 12900 9104
rect 12492 9064 12900 9092
rect 12492 9052 12498 9064
rect 12894 9052 12900 9064
rect 12952 9052 12958 9104
rect 12529 9027 12587 9033
rect 12529 8993 12541 9027
rect 12575 9024 12587 9027
rect 12802 9024 12808 9036
rect 12575 8996 12808 9024
rect 12575 8993 12587 8996
rect 12529 8987 12587 8993
rect 12802 8984 12808 8996
rect 12860 8984 12866 9036
rect 13265 9027 13323 9033
rect 13265 8993 13277 9027
rect 13311 9024 13323 9027
rect 14458 9024 14464 9036
rect 13311 8996 14464 9024
rect 13311 8993 13323 8996
rect 13265 8987 13323 8993
rect 14458 8984 14464 8996
rect 14516 8984 14522 9036
rect 12253 8959 12311 8965
rect 11388 8928 12204 8956
rect 11388 8916 11394 8928
rect 10091 8860 10640 8888
rect 10796 8888 10824 8916
rect 11974 8888 11980 8900
rect 10796 8860 11980 8888
rect 10091 8857 10103 8860
rect 10045 8851 10103 8857
rect 11974 8848 11980 8860
rect 12032 8848 12038 8900
rect 12176 8888 12204 8928
rect 12253 8925 12265 8959
rect 12299 8925 12311 8959
rect 12710 8956 12716 8968
rect 12671 8928 12716 8956
rect 12253 8919 12311 8925
rect 12710 8916 12716 8928
rect 12768 8916 12774 8968
rect 13633 8959 13691 8965
rect 13633 8956 13645 8959
rect 12912 8928 13645 8956
rect 12805 8891 12863 8897
rect 12805 8888 12817 8891
rect 12176 8860 12817 8888
rect 12805 8857 12817 8860
rect 12851 8857 12863 8891
rect 12805 8851 12863 8857
rect 9950 8820 9956 8832
rect 9324 8792 9956 8820
rect 9217 8783 9275 8789
rect 9950 8780 9956 8792
rect 10008 8780 10014 8832
rect 10134 8780 10140 8832
rect 10192 8820 10198 8832
rect 11333 8823 11391 8829
rect 11333 8820 11345 8823
rect 10192 8792 11345 8820
rect 10192 8780 10198 8792
rect 11333 8789 11345 8792
rect 11379 8820 11391 8823
rect 12066 8820 12072 8832
rect 11379 8792 12072 8820
rect 11379 8789 11391 8792
rect 11333 8783 11391 8789
rect 12066 8780 12072 8792
rect 12124 8780 12130 8832
rect 12250 8780 12256 8832
rect 12308 8820 12314 8832
rect 12345 8823 12403 8829
rect 12345 8820 12357 8823
rect 12308 8792 12357 8820
rect 12308 8780 12314 8792
rect 12345 8789 12357 8792
rect 12391 8820 12403 8823
rect 12618 8820 12624 8832
rect 12391 8792 12624 8820
rect 12391 8789 12403 8792
rect 12345 8783 12403 8789
rect 12618 8780 12624 8792
rect 12676 8780 12682 8832
rect 12912 8829 12940 8928
rect 13633 8925 13645 8928
rect 13679 8925 13691 8959
rect 14568 8956 14596 9132
rect 15473 9129 15485 9163
rect 15519 9160 15531 9163
rect 17402 9160 17408 9172
rect 15519 9132 17408 9160
rect 15519 9129 15531 9132
rect 15473 9123 15531 9129
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 14734 8984 14740 9036
rect 14792 9024 14798 9036
rect 17589 9027 17647 9033
rect 17589 9024 17601 9027
rect 14792 8996 17601 9024
rect 14792 8984 14798 8996
rect 17589 8993 17601 8996
rect 17635 8993 17647 9027
rect 17589 8987 17647 8993
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 14568 8928 15301 8956
rect 13633 8919 13691 8925
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 15473 8959 15531 8965
rect 15473 8925 15485 8959
rect 15519 8956 15531 8959
rect 15930 8956 15936 8968
rect 15519 8928 15936 8956
rect 15519 8925 15531 8928
rect 15473 8919 15531 8925
rect 12989 8891 13047 8897
rect 12989 8857 13001 8891
rect 13035 8888 13047 8891
rect 13170 8888 13176 8900
rect 13035 8860 13176 8888
rect 13035 8857 13047 8860
rect 12989 8851 13047 8857
rect 13170 8848 13176 8860
rect 13228 8848 13234 8900
rect 15194 8888 15200 8900
rect 14674 8874 15200 8888
rect 14660 8860 15200 8874
rect 12897 8823 12955 8829
rect 12897 8789 12909 8823
rect 12943 8789 12955 8823
rect 12897 8783 12955 8789
rect 13630 8780 13636 8832
rect 13688 8820 13694 8832
rect 14660 8820 14688 8860
rect 15194 8848 15200 8860
rect 15252 8848 15258 8900
rect 13688 8792 14688 8820
rect 13688 8780 13694 8792
rect 14918 8780 14924 8832
rect 14976 8820 14982 8832
rect 15059 8823 15117 8829
rect 15059 8820 15071 8823
rect 14976 8792 15071 8820
rect 14976 8780 14982 8792
rect 15059 8789 15071 8792
rect 15105 8789 15117 8823
rect 15304 8820 15332 8919
rect 15930 8916 15936 8928
rect 15988 8916 15994 8968
rect 17862 8916 17868 8968
rect 17920 8956 17926 8968
rect 17920 8928 17965 8956
rect 17920 8916 17926 8928
rect 15841 8891 15899 8897
rect 15841 8888 15853 8891
rect 15580 8860 15853 8888
rect 15580 8820 15608 8860
rect 15841 8857 15853 8860
rect 15887 8857 15899 8891
rect 15841 8851 15899 8857
rect 15304 8792 15608 8820
rect 15749 8823 15807 8829
rect 15059 8783 15117 8789
rect 15749 8789 15761 8823
rect 15795 8820 15807 8823
rect 16206 8820 16212 8832
rect 15795 8792 16212 8820
rect 15795 8789 15807 8792
rect 15749 8783 15807 8789
rect 16206 8780 16212 8792
rect 16264 8820 16270 8832
rect 16408 8820 16436 8874
rect 16264 8792 16436 8820
rect 16264 8780 16270 8792
rect 0 8730 18860 8752
rect 0 8678 4660 8730
rect 4712 8678 4724 8730
rect 4776 8678 4788 8730
rect 4840 8678 4852 8730
rect 4904 8678 4916 8730
rect 4968 8678 7760 8730
rect 7812 8678 7824 8730
rect 7876 8678 7888 8730
rect 7940 8678 7952 8730
rect 8004 8678 8016 8730
rect 8068 8678 10860 8730
rect 10912 8678 10924 8730
rect 10976 8678 10988 8730
rect 11040 8678 11052 8730
rect 11104 8678 11116 8730
rect 11168 8678 13960 8730
rect 14012 8678 14024 8730
rect 14076 8678 14088 8730
rect 14140 8678 14152 8730
rect 14204 8678 14216 8730
rect 14268 8678 17060 8730
rect 17112 8678 17124 8730
rect 17176 8678 17188 8730
rect 17240 8678 17252 8730
rect 17304 8678 17316 8730
rect 17368 8678 18860 8730
rect 0 8656 18860 8678
rect 2038 8576 2044 8628
rect 2096 8616 2102 8628
rect 2133 8619 2191 8625
rect 2133 8616 2145 8619
rect 2096 8588 2145 8616
rect 2096 8576 2102 8588
rect 2133 8585 2145 8588
rect 2179 8585 2191 8619
rect 2133 8579 2191 8585
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 3145 8619 3203 8625
rect 3145 8616 3157 8619
rect 2372 8588 3157 8616
rect 2372 8576 2378 8588
rect 3145 8585 3157 8588
rect 3191 8585 3203 8619
rect 3145 8579 3203 8585
rect 3513 8619 3571 8625
rect 3513 8585 3525 8619
rect 3559 8616 3571 8619
rect 3973 8619 4031 8625
rect 3973 8616 3985 8619
rect 3559 8588 3985 8616
rect 3559 8585 3571 8588
rect 3513 8579 3571 8585
rect 3973 8585 3985 8588
rect 4019 8585 4031 8619
rect 3973 8579 4031 8585
rect 6181 8619 6239 8625
rect 6181 8585 6193 8619
rect 6227 8616 6239 8619
rect 6638 8616 6644 8628
rect 6227 8588 6644 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 8754 8616 8760 8628
rect 6840 8588 8760 8616
rect 2222 8548 2228 8560
rect 1794 8520 2228 8548
rect 2222 8508 2228 8520
rect 2280 8508 2286 8560
rect 2590 8548 2596 8560
rect 2332 8520 2596 8548
rect 2130 8480 2136 8492
rect 2091 8452 2136 8480
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 2332 8489 2360 8520
rect 2590 8508 2596 8520
rect 2648 8508 2654 8560
rect 2774 8508 2780 8560
rect 2832 8548 2838 8560
rect 5261 8551 5319 8557
rect 5261 8548 5273 8551
rect 2832 8520 5273 8548
rect 2832 8508 2838 8520
rect 5261 8517 5273 8520
rect 5307 8517 5319 8551
rect 5534 8548 5540 8560
rect 5261 8511 5319 8517
rect 5368 8520 5540 8548
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8449 2375 8483
rect 2682 8480 2688 8492
rect 2643 8452 2688 8480
rect 2317 8443 2375 8449
rect 2682 8440 2688 8452
rect 2740 8440 2746 8492
rect 4341 8483 4399 8489
rect 4341 8480 4353 8483
rect 3068 8452 4353 8480
rect 290 8412 296 8424
rect 251 8384 296 8412
rect 290 8372 296 8384
rect 348 8372 354 8424
rect 566 8412 572 8424
rect 527 8384 572 8412
rect 566 8372 572 8384
rect 624 8372 630 8424
rect 2593 8415 2651 8421
rect 2593 8412 2605 8415
rect 2056 8384 2605 8412
rect 2056 8288 2084 8384
rect 2593 8381 2605 8384
rect 2639 8412 2651 8415
rect 2866 8412 2872 8424
rect 2639 8384 2872 8412
rect 2639 8381 2651 8384
rect 2593 8375 2651 8381
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 3068 8353 3096 8452
rect 4341 8449 4353 8452
rect 4387 8449 4399 8483
rect 5166 8480 5172 8492
rect 5127 8452 5172 8480
rect 4341 8443 4399 8449
rect 5166 8440 5172 8452
rect 5224 8440 5230 8492
rect 5368 8489 5396 8520
rect 5534 8508 5540 8520
rect 5592 8548 5598 8560
rect 6273 8551 6331 8557
rect 6273 8548 6285 8551
rect 5592 8520 6285 8548
rect 5592 8508 5598 8520
rect 6273 8517 6285 8520
rect 6319 8548 6331 8551
rect 6546 8548 6552 8560
rect 6319 8520 6552 8548
rect 6319 8517 6331 8520
rect 6273 8511 6331 8517
rect 6546 8508 6552 8520
rect 6604 8508 6610 8560
rect 6840 8548 6868 8588
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 8849 8619 8907 8625
rect 8849 8585 8861 8619
rect 8895 8616 8907 8619
rect 8938 8616 8944 8628
rect 8895 8588 8944 8616
rect 8895 8585 8907 8588
rect 8849 8579 8907 8585
rect 8938 8576 8944 8588
rect 8996 8616 9002 8628
rect 9582 8616 9588 8628
rect 8996 8588 9588 8616
rect 8996 8576 9002 8588
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 10226 8576 10232 8628
rect 10284 8616 10290 8628
rect 10321 8619 10379 8625
rect 10321 8616 10333 8619
rect 10284 8588 10333 8616
rect 10284 8576 10290 8588
rect 10321 8585 10333 8588
rect 10367 8585 10379 8619
rect 10321 8579 10379 8585
rect 10686 8576 10692 8628
rect 10744 8616 10750 8628
rect 10781 8619 10839 8625
rect 10781 8616 10793 8619
rect 10744 8588 10793 8616
rect 10744 8576 10750 8588
rect 10781 8585 10793 8588
rect 10827 8585 10839 8619
rect 10781 8579 10839 8585
rect 10873 8619 10931 8625
rect 10873 8585 10885 8619
rect 10919 8616 10931 8619
rect 12158 8616 12164 8628
rect 10919 8588 12164 8616
rect 10919 8585 10931 8588
rect 10873 8579 10931 8585
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 12710 8576 12716 8628
rect 12768 8616 12774 8628
rect 12805 8619 12863 8625
rect 12805 8616 12817 8619
rect 12768 8588 12817 8616
rect 12768 8576 12774 8588
rect 12805 8585 12817 8588
rect 12851 8585 12863 8619
rect 13170 8616 13176 8628
rect 13131 8588 13176 8616
rect 12805 8579 12863 8585
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 13630 8616 13636 8628
rect 13591 8588 13636 8616
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 14458 8576 14464 8628
rect 14516 8616 14522 8628
rect 17313 8619 17371 8625
rect 17313 8616 17325 8619
rect 14516 8588 17325 8616
rect 14516 8576 14522 8588
rect 17313 8585 17325 8588
rect 17359 8585 17371 8619
rect 17313 8579 17371 8585
rect 6748 8520 6868 8548
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8449 5411 8483
rect 5718 8480 5724 8492
rect 5631 8452 5724 8480
rect 5353 8443 5411 8449
rect 5718 8440 5724 8452
rect 5776 8480 5782 8492
rect 6748 8489 6776 8520
rect 7650 8508 7656 8560
rect 7708 8557 7714 8560
rect 7708 8551 7772 8557
rect 7708 8517 7726 8551
rect 7760 8517 7772 8551
rect 10502 8548 10508 8560
rect 7708 8511 7772 8517
rect 8036 8520 10508 8548
rect 7708 8508 7714 8511
rect 6733 8483 6791 8489
rect 5776 8452 6132 8480
rect 5776 8440 5782 8452
rect 3605 8415 3663 8421
rect 3605 8381 3617 8415
rect 3651 8381 3663 8415
rect 3605 8375 3663 8381
rect 3053 8347 3111 8353
rect 3053 8313 3065 8347
rect 3099 8313 3111 8347
rect 3620 8344 3648 8375
rect 3694 8372 3700 8424
rect 3752 8412 3758 8424
rect 4433 8415 4491 8421
rect 4433 8412 4445 8415
rect 3752 8384 3797 8412
rect 3896 8384 4445 8412
rect 3752 8372 3758 8384
rect 3896 8356 3924 8384
rect 4433 8381 4445 8384
rect 4479 8381 4491 8415
rect 4433 8375 4491 8381
rect 4525 8415 4583 8421
rect 4525 8381 4537 8415
rect 4571 8381 4583 8415
rect 4525 8375 4583 8381
rect 3878 8344 3884 8356
rect 3620 8316 3884 8344
rect 3053 8307 3111 8313
rect 3878 8304 3884 8316
rect 3936 8304 3942 8356
rect 4062 8344 4068 8356
rect 3975 8316 4068 8344
rect 4062 8304 4068 8316
rect 4120 8344 4126 8356
rect 4540 8344 4568 8375
rect 5810 8372 5816 8424
rect 5868 8412 5874 8424
rect 5997 8415 6055 8421
rect 5997 8412 6009 8415
rect 5868 8384 6009 8412
rect 5868 8372 5874 8384
rect 5997 8381 6009 8384
rect 6043 8381 6055 8415
rect 5997 8375 6055 8381
rect 4120 8316 4568 8344
rect 4120 8304 4126 8316
rect 2038 8276 2044 8288
rect 1999 8248 2044 8276
rect 2038 8236 2044 8248
rect 2096 8236 2102 8288
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 4080 8276 4108 8304
rect 3016 8248 4108 8276
rect 3016 8236 3022 8248
rect 5166 8236 5172 8288
rect 5224 8276 5230 8288
rect 5813 8279 5871 8285
rect 5813 8276 5825 8279
rect 5224 8248 5825 8276
rect 5224 8236 5230 8248
rect 5813 8245 5825 8248
rect 5859 8245 5871 8279
rect 5813 8239 5871 8245
rect 5902 8236 5908 8288
rect 5960 8276 5966 8288
rect 6104 8276 6132 8452
rect 6733 8449 6745 8483
rect 6779 8449 6791 8483
rect 8036 8480 8064 8520
rect 10502 8508 10508 8520
rect 10560 8508 10566 8560
rect 10704 8520 12296 8548
rect 6733 8443 6791 8449
rect 6840 8452 8064 8480
rect 6840 8421 6868 8452
rect 8202 8440 8208 8492
rect 8260 8480 8266 8492
rect 9203 8483 9261 8489
rect 9203 8480 9215 8483
rect 8260 8452 9215 8480
rect 8260 8440 8266 8452
rect 9203 8449 9215 8452
rect 9249 8480 9261 8483
rect 9249 8452 9536 8480
rect 9249 8449 9261 8452
rect 9203 8443 9261 8449
rect 6825 8415 6883 8421
rect 6825 8381 6837 8415
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 7101 8415 7159 8421
rect 7101 8381 7113 8415
rect 7147 8412 7159 8415
rect 7190 8412 7196 8424
rect 7147 8384 7196 8412
rect 7147 8381 7159 8384
rect 7101 8375 7159 8381
rect 7190 8372 7196 8384
rect 7248 8372 7254 8424
rect 7466 8412 7472 8424
rect 7427 8384 7472 8412
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 8754 8372 8760 8424
rect 8812 8412 8818 8424
rect 9125 8415 9183 8421
rect 9125 8412 9137 8415
rect 8812 8384 9137 8412
rect 8812 8372 8818 8384
rect 9125 8381 9137 8384
rect 9171 8404 9183 8415
rect 9398 8412 9404 8424
rect 9232 8404 9404 8412
rect 9171 8384 9404 8404
rect 9171 8381 9260 8384
rect 9125 8376 9260 8381
rect 9125 8375 9183 8376
rect 9398 8372 9404 8384
rect 9456 8372 9462 8424
rect 9508 8412 9536 8452
rect 9582 8440 9588 8492
rect 9640 8480 9646 8492
rect 9677 8483 9735 8489
rect 9677 8480 9689 8483
rect 9640 8452 9689 8480
rect 9640 8440 9646 8452
rect 9677 8449 9689 8452
rect 9723 8449 9735 8483
rect 9677 8443 9735 8449
rect 9858 8440 9864 8492
rect 9916 8480 9922 8492
rect 10704 8480 10732 8520
rect 9916 8452 10732 8480
rect 11701 8483 11759 8489
rect 9916 8440 9922 8452
rect 11701 8449 11713 8483
rect 11747 8480 11759 8483
rect 11790 8480 11796 8492
rect 11747 8452 11796 8480
rect 11747 8449 11759 8452
rect 11701 8443 11759 8449
rect 11790 8440 11796 8452
rect 11848 8484 11854 8492
rect 11848 8480 11928 8484
rect 11848 8452 11941 8480
rect 11848 8440 11854 8452
rect 10594 8412 10600 8424
rect 9508 8384 10600 8412
rect 10594 8372 10600 8384
rect 10652 8372 10658 8424
rect 10689 8415 10747 8421
rect 10689 8381 10701 8415
rect 10735 8412 10747 8415
rect 11514 8412 11520 8424
rect 10735 8384 11520 8412
rect 10735 8381 10747 8384
rect 10689 8375 10747 8381
rect 11514 8372 11520 8384
rect 11572 8372 11578 8424
rect 11900 8412 11928 8452
rect 11974 8440 11980 8492
rect 12032 8480 12038 8492
rect 12268 8489 12296 8520
rect 12342 8508 12348 8560
rect 12400 8548 12406 8560
rect 14553 8551 14611 8557
rect 14553 8548 14565 8551
rect 12400 8520 12572 8548
rect 12400 8508 12406 8520
rect 12544 8489 12572 8520
rect 12820 8520 14565 8548
rect 12069 8483 12127 8489
rect 12069 8480 12081 8483
rect 12032 8452 12081 8480
rect 12032 8440 12038 8452
rect 12069 8449 12081 8452
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 12529 8483 12587 8489
rect 12529 8449 12541 8483
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 12621 8483 12679 8489
rect 12621 8449 12633 8483
rect 12667 8478 12679 8483
rect 12820 8480 12848 8520
rect 12728 8478 12848 8480
rect 12667 8452 12848 8478
rect 12667 8450 12756 8452
rect 12667 8449 12679 8450
rect 12621 8443 12679 8449
rect 12452 8412 12480 8443
rect 12894 8440 12900 8492
rect 12952 8480 12958 8492
rect 13372 8489 13400 8520
rect 14553 8517 14565 8520
rect 14599 8517 14611 8551
rect 14553 8511 14611 8517
rect 16206 8508 16212 8560
rect 16264 8508 16270 8560
rect 16942 8508 16948 8560
rect 17000 8548 17006 8560
rect 17221 8551 17279 8557
rect 17221 8548 17233 8551
rect 17000 8520 17233 8548
rect 17000 8508 17006 8520
rect 17221 8517 17233 8520
rect 17267 8517 17279 8551
rect 17221 8511 17279 8517
rect 13081 8483 13139 8489
rect 12952 8452 12997 8480
rect 12952 8440 12958 8452
rect 13081 8449 13093 8483
rect 13127 8449 13139 8483
rect 13081 8443 13139 8449
rect 13357 8483 13415 8489
rect 13357 8449 13369 8483
rect 13403 8449 13415 8483
rect 13357 8443 13415 8449
rect 13909 8483 13967 8489
rect 13909 8449 13921 8483
rect 13955 8480 13967 8483
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 13955 8452 14657 8480
rect 13955 8449 13967 8452
rect 13909 8443 13967 8449
rect 14645 8449 14657 8452
rect 14691 8480 14703 8483
rect 14918 8480 14924 8492
rect 14691 8452 14924 8480
rect 14691 8449 14703 8452
rect 14645 8443 14703 8449
rect 13096 8412 13124 8443
rect 14918 8440 14924 8452
rect 14976 8440 14982 8492
rect 18233 8483 18291 8489
rect 16500 8452 16988 8480
rect 13814 8412 13820 8424
rect 11900 8384 13124 8412
rect 13775 8384 13820 8412
rect 13814 8372 13820 8384
rect 13872 8372 13878 8424
rect 14829 8415 14887 8421
rect 14829 8381 14841 8415
rect 14875 8381 14887 8415
rect 14829 8375 14887 8381
rect 15197 8415 15255 8421
rect 15197 8381 15209 8415
rect 15243 8412 15255 8415
rect 16500 8412 16528 8452
rect 15243 8384 16528 8412
rect 15243 8381 15255 8384
rect 15197 8375 15255 8381
rect 9493 8347 9551 8353
rect 9493 8313 9505 8347
rect 9539 8344 9551 8347
rect 11146 8344 11152 8356
rect 9539 8316 11152 8344
rect 9539 8313 9551 8316
rect 9493 8307 9551 8313
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 11241 8347 11299 8353
rect 11241 8313 11253 8347
rect 11287 8344 11299 8347
rect 12342 8344 12348 8356
rect 11287 8316 12348 8344
rect 11287 8313 11299 8316
rect 11241 8307 11299 8313
rect 12342 8304 12348 8316
rect 12400 8304 12406 8356
rect 12618 8304 12624 8356
rect 12676 8344 12682 8356
rect 12676 8316 12848 8344
rect 12676 8304 12682 8316
rect 10134 8276 10140 8288
rect 5960 8248 6005 8276
rect 6104 8248 10140 8276
rect 5960 8236 5966 8248
rect 10134 8236 10140 8248
rect 10192 8236 10198 8288
rect 11422 8236 11428 8288
rect 11480 8276 11486 8288
rect 11609 8279 11667 8285
rect 11609 8276 11621 8279
rect 11480 8248 11621 8276
rect 11480 8236 11486 8248
rect 11609 8245 11621 8248
rect 11655 8245 11667 8279
rect 11609 8239 11667 8245
rect 11882 8236 11888 8288
rect 11940 8276 11946 8288
rect 12069 8279 12127 8285
rect 12069 8276 12081 8279
rect 11940 8248 12081 8276
rect 11940 8236 11946 8248
rect 12069 8245 12081 8248
rect 12115 8245 12127 8279
rect 12820 8276 12848 8316
rect 12894 8304 12900 8356
rect 12952 8344 12958 8356
rect 13998 8344 14004 8356
rect 12952 8316 14004 8344
rect 12952 8304 12958 8316
rect 13998 8304 14004 8316
rect 14056 8304 14062 8356
rect 14277 8347 14335 8353
rect 14277 8313 14289 8347
rect 14323 8344 14335 8347
rect 14642 8344 14648 8356
rect 14323 8316 14648 8344
rect 14323 8313 14335 8316
rect 14277 8307 14335 8313
rect 14642 8304 14648 8316
rect 14700 8304 14706 8356
rect 14844 8288 14872 8375
rect 16574 8372 16580 8424
rect 16632 8412 16638 8424
rect 16632 8384 16896 8412
rect 16632 8372 16638 8384
rect 16868 8353 16896 8384
rect 16853 8347 16911 8353
rect 16853 8313 16865 8347
rect 16899 8313 16911 8347
rect 16960 8344 16988 8452
rect 18233 8449 18245 8483
rect 18279 8480 18291 8483
rect 18509 8483 18567 8489
rect 18509 8480 18521 8483
rect 18279 8452 18521 8480
rect 18279 8449 18291 8452
rect 18233 8443 18291 8449
rect 18509 8449 18521 8452
rect 18555 8480 18567 8483
rect 18598 8480 18604 8492
rect 18555 8452 18604 8480
rect 18555 8449 18567 8452
rect 18509 8443 18567 8449
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 17402 8412 17408 8424
rect 17363 8384 17408 8412
rect 17402 8372 17408 8384
rect 17460 8372 17466 8424
rect 18325 8347 18383 8353
rect 18325 8344 18337 8347
rect 16960 8316 18337 8344
rect 16853 8307 16911 8313
rect 18325 8313 18337 8316
rect 18371 8313 18383 8347
rect 18325 8307 18383 8313
rect 14826 8276 14832 8288
rect 12820 8248 14832 8276
rect 12069 8239 12127 8245
rect 14826 8236 14832 8248
rect 14884 8236 14890 8288
rect 16623 8279 16681 8285
rect 16623 8245 16635 8279
rect 16669 8276 16681 8279
rect 16758 8276 16764 8288
rect 16669 8248 16764 8276
rect 16669 8245 16681 8248
rect 16623 8239 16681 8245
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 0 8186 18860 8208
rect 0 8134 3110 8186
rect 3162 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 3302 8186
rect 3354 8134 3366 8186
rect 3418 8134 6210 8186
rect 6262 8134 6274 8186
rect 6326 8134 6338 8186
rect 6390 8134 6402 8186
rect 6454 8134 6466 8186
rect 6518 8134 9310 8186
rect 9362 8134 9374 8186
rect 9426 8134 9438 8186
rect 9490 8134 9502 8186
rect 9554 8134 9566 8186
rect 9618 8134 12410 8186
rect 12462 8134 12474 8186
rect 12526 8134 12538 8186
rect 12590 8134 12602 8186
rect 12654 8134 12666 8186
rect 12718 8134 15510 8186
rect 15562 8134 15574 8186
rect 15626 8134 15638 8186
rect 15690 8134 15702 8186
rect 15754 8134 15766 8186
rect 15818 8134 18860 8186
rect 0 8112 18860 8134
rect 566 8032 572 8084
rect 624 8072 630 8084
rect 1397 8075 1455 8081
rect 1397 8072 1409 8075
rect 624 8044 1409 8072
rect 624 8032 630 8044
rect 1397 8041 1409 8044
rect 1443 8041 1455 8075
rect 1397 8035 1455 8041
rect 1489 8075 1547 8081
rect 1489 8041 1501 8075
rect 1535 8072 1547 8075
rect 2130 8072 2136 8084
rect 1535 8044 2136 8072
rect 1535 8041 1547 8044
rect 1489 8035 1547 8041
rect 2130 8032 2136 8044
rect 2188 8032 2194 8084
rect 2314 8032 2320 8084
rect 2372 8072 2378 8084
rect 2409 8075 2467 8081
rect 2409 8072 2421 8075
rect 2372 8044 2421 8072
rect 2372 8032 2378 8044
rect 2409 8041 2421 8044
rect 2455 8041 2467 8075
rect 2409 8035 2467 8041
rect 2498 8032 2504 8084
rect 2556 8072 2562 8084
rect 2556 8044 2601 8072
rect 2556 8032 2562 8044
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 9766 8072 9772 8084
rect 4304 8044 9772 8072
rect 4304 8032 4310 8044
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 11790 8072 11796 8084
rect 11751 8044 11796 8072
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 18506 8072 18512 8084
rect 11992 8044 18512 8072
rect 3694 8004 3700 8016
rect 1872 7976 3700 8004
rect 1302 7936 1308 7948
rect 1263 7908 1308 7936
rect 1302 7896 1308 7908
rect 1360 7896 1366 7948
rect 1872 7945 1900 7976
rect 3694 7964 3700 7976
rect 3752 7964 3758 8016
rect 5534 7964 5540 8016
rect 5592 8004 5598 8016
rect 5629 8007 5687 8013
rect 5629 8004 5641 8007
rect 5592 7976 5641 8004
rect 5592 7964 5598 7976
rect 5629 7973 5641 7976
rect 5675 7973 5687 8007
rect 5629 7967 5687 7973
rect 1857 7939 1915 7945
rect 1857 7905 1869 7939
rect 1903 7905 1915 7939
rect 1857 7899 1915 7905
rect 2958 7896 2964 7948
rect 3016 7936 3022 7948
rect 3053 7939 3111 7945
rect 3053 7936 3065 7939
rect 3016 7908 3065 7936
rect 3016 7896 3022 7908
rect 3053 7905 3065 7908
rect 3099 7905 3111 7939
rect 3053 7899 3111 7905
rect 6641 7939 6699 7945
rect 6641 7905 6653 7939
rect 6687 7936 6699 7939
rect 7558 7936 7564 7948
rect 6687 7908 7564 7936
rect 6687 7905 6699 7908
rect 6641 7899 6699 7905
rect 7558 7896 7564 7908
rect 7616 7896 7622 7948
rect 8846 7936 8852 7948
rect 8807 7908 8852 7936
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 11422 7936 11428 7948
rect 11383 7908 11428 7936
rect 11422 7896 11428 7908
rect 11480 7896 11486 7948
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 1946 7868 1952 7880
rect 1627 7840 1952 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 1946 7828 1952 7840
rect 2004 7868 2010 7880
rect 2869 7871 2927 7877
rect 2869 7868 2881 7871
rect 2004 7840 2881 7868
rect 2004 7828 2010 7840
rect 2869 7837 2881 7840
rect 2915 7837 2927 7871
rect 2869 7831 2927 7837
rect 3694 7828 3700 7880
rect 3752 7868 3758 7880
rect 5445 7871 5503 7877
rect 5445 7868 5457 7871
rect 3752 7840 5457 7868
rect 3752 7828 3758 7840
rect 5445 7837 5457 7840
rect 5491 7837 5503 7871
rect 5445 7831 5503 7837
rect 6086 7828 6092 7880
rect 6144 7868 6150 7880
rect 6273 7871 6331 7877
rect 6273 7868 6285 7871
rect 6144 7840 6285 7868
rect 6144 7828 6150 7840
rect 6273 7837 6285 7840
rect 6319 7837 6331 7871
rect 6273 7831 6331 7837
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 11241 7871 11299 7877
rect 11241 7868 11253 7871
rect 11204 7840 11253 7868
rect 11204 7828 11210 7840
rect 11241 7837 11253 7840
rect 11287 7837 11299 7871
rect 11698 7868 11704 7880
rect 11659 7840 11704 7868
rect 11241 7831 11299 7837
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 11882 7868 11888 7880
rect 11843 7840 11888 7868
rect 11882 7828 11888 7840
rect 11940 7828 11946 7880
rect 2041 7803 2099 7809
rect 2041 7769 2053 7803
rect 2087 7800 2099 7803
rect 2498 7800 2504 7812
rect 2087 7772 2504 7800
rect 2087 7769 2099 7772
rect 2041 7763 2099 7769
rect 2498 7760 2504 7772
rect 2556 7760 2562 7812
rect 7374 7760 7380 7812
rect 7432 7760 7438 7812
rect 11992 7809 12020 8044
rect 18506 8032 18512 8044
rect 18564 8032 18570 8084
rect 12066 7964 12072 8016
rect 12124 8004 12130 8016
rect 13357 8007 13415 8013
rect 12124 7976 13032 8004
rect 12124 7964 12130 7976
rect 13004 7945 13032 7976
rect 13357 7973 13369 8007
rect 13403 8004 13415 8007
rect 13630 8004 13636 8016
rect 13403 7976 13636 8004
rect 13403 7973 13415 7976
rect 13357 7967 13415 7973
rect 13630 7964 13636 7976
rect 13688 7964 13694 8016
rect 15749 8007 15807 8013
rect 15749 8004 15761 8007
rect 14200 7976 15761 8004
rect 12989 7939 13047 7945
rect 12406 7908 12940 7936
rect 12406 7868 12434 7908
rect 12912 7877 12940 7908
rect 12989 7905 13001 7939
rect 13035 7905 13047 7939
rect 14200 7936 14228 7976
rect 15749 7973 15761 7976
rect 15795 8004 15807 8007
rect 15930 8004 15936 8016
rect 15795 7976 15936 8004
rect 15795 7973 15807 7976
rect 15749 7967 15807 7973
rect 15930 7964 15936 7976
rect 15988 7964 15994 8016
rect 14366 7936 14372 7948
rect 12989 7899 13047 7905
rect 13188 7908 14228 7936
rect 14279 7908 14372 7936
rect 12084 7840 12434 7868
rect 12713 7871 12771 7877
rect 10597 7803 10655 7809
rect 10597 7769 10609 7803
rect 10643 7800 10655 7803
rect 11977 7803 12035 7809
rect 11977 7800 11989 7803
rect 10643 7772 11989 7800
rect 10643 7769 10655 7772
rect 10597 7763 10655 7769
rect 11977 7769 11989 7772
rect 12023 7769 12035 7803
rect 11977 7763 12035 7769
rect 1949 7735 2007 7741
rect 1949 7701 1961 7735
rect 1995 7732 2007 7735
rect 2961 7735 3019 7741
rect 2961 7732 2973 7735
rect 1995 7704 2973 7732
rect 1995 7701 2007 7704
rect 1949 7695 2007 7701
rect 2961 7701 2973 7704
rect 3007 7732 3019 7735
rect 3786 7732 3792 7744
rect 3007 7704 3792 7732
rect 3007 7701 3019 7704
rect 2961 7695 3019 7701
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 6181 7735 6239 7741
rect 6181 7701 6193 7735
rect 6227 7732 6239 7735
rect 6914 7732 6920 7744
rect 6227 7704 6920 7732
rect 6227 7701 6239 7704
rect 6181 7695 6239 7701
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 7098 7692 7104 7744
rect 7156 7732 7162 7744
rect 8067 7735 8125 7741
rect 8067 7732 8079 7735
rect 7156 7704 8079 7732
rect 7156 7692 7162 7704
rect 8067 7701 8079 7704
rect 8113 7732 8125 7735
rect 8202 7732 8208 7744
rect 8113 7704 8208 7732
rect 8113 7701 8125 7704
rect 8067 7695 8125 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 9122 7692 9128 7744
rect 9180 7732 9186 7744
rect 10873 7735 10931 7741
rect 10873 7732 10885 7735
rect 9180 7704 10885 7732
rect 9180 7692 9186 7704
rect 10873 7701 10885 7704
rect 10919 7701 10931 7735
rect 10873 7695 10931 7701
rect 11238 7692 11244 7744
rect 11296 7732 11302 7744
rect 11333 7735 11391 7741
rect 11333 7732 11345 7735
rect 11296 7704 11345 7732
rect 11296 7692 11302 7704
rect 11333 7701 11345 7704
rect 11379 7732 11391 7735
rect 12084 7732 12112 7840
rect 12713 7837 12725 7871
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7868 12955 7871
rect 13188 7868 13216 7908
rect 14366 7896 14372 7908
rect 14424 7936 14430 7948
rect 15197 7939 15255 7945
rect 15197 7936 15209 7939
rect 14424 7908 15209 7936
rect 14424 7896 14430 7908
rect 15197 7905 15209 7908
rect 15243 7905 15255 7939
rect 16574 7936 16580 7948
rect 15197 7899 15255 7905
rect 15304 7908 16580 7936
rect 12943 7840 13216 7868
rect 13909 7871 13967 7877
rect 12943 7837 12955 7840
rect 12897 7831 12955 7837
rect 13909 7837 13921 7871
rect 13955 7837 13967 7871
rect 13909 7831 13967 7837
rect 12158 7760 12164 7812
rect 12216 7800 12222 7812
rect 12728 7800 12756 7831
rect 13924 7800 13952 7831
rect 13998 7828 14004 7880
rect 14056 7868 14062 7880
rect 14461 7871 14519 7877
rect 14461 7868 14473 7871
rect 14056 7840 14473 7868
rect 14056 7828 14062 7840
rect 14461 7837 14473 7840
rect 14507 7837 14519 7871
rect 14642 7868 14648 7880
rect 14603 7840 14648 7868
rect 14461 7831 14519 7837
rect 14642 7828 14648 7840
rect 14700 7828 14706 7880
rect 14826 7828 14832 7880
rect 14884 7868 14890 7880
rect 15304 7877 15332 7908
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 16758 7896 16764 7948
rect 16816 7936 16822 7948
rect 17497 7939 17555 7945
rect 17497 7936 17509 7939
rect 16816 7908 17509 7936
rect 16816 7896 16822 7908
rect 17497 7905 17509 7908
rect 17543 7905 17555 7939
rect 17497 7899 17555 7905
rect 14921 7871 14979 7877
rect 14921 7868 14933 7871
rect 14884 7840 14933 7868
rect 14884 7828 14890 7840
rect 14921 7837 14933 7840
rect 14967 7837 14979 7871
rect 14921 7831 14979 7837
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7837 15347 7871
rect 17862 7868 17868 7880
rect 17775 7840 17868 7868
rect 15289 7831 15347 7837
rect 14734 7800 14740 7812
rect 12216 7772 14740 7800
rect 12216 7760 12222 7772
rect 14734 7760 14740 7772
rect 14792 7760 14798 7812
rect 11379 7704 12112 7732
rect 11379 7701 11391 7704
rect 11333 7695 11391 7701
rect 12250 7692 12256 7744
rect 12308 7732 12314 7744
rect 12529 7735 12587 7741
rect 12529 7732 12541 7735
rect 12308 7704 12541 7732
rect 12308 7692 12314 7704
rect 12529 7701 12541 7704
rect 12575 7701 12587 7735
rect 14936 7732 14964 7831
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 16298 7760 16304 7812
rect 16356 7800 16362 7812
rect 16356 7772 16514 7800
rect 16356 7760 16362 7772
rect 17880 7732 17908 7828
rect 14936 7704 17908 7732
rect 12529 7695 12587 7701
rect 0 7642 18860 7664
rect 0 7590 4660 7642
rect 4712 7590 4724 7642
rect 4776 7590 4788 7642
rect 4840 7590 4852 7642
rect 4904 7590 4916 7642
rect 4968 7590 7760 7642
rect 7812 7590 7824 7642
rect 7876 7590 7888 7642
rect 7940 7590 7952 7642
rect 8004 7590 8016 7642
rect 8068 7590 10860 7642
rect 10912 7590 10924 7642
rect 10976 7590 10988 7642
rect 11040 7590 11052 7642
rect 11104 7590 11116 7642
rect 11168 7590 13960 7642
rect 14012 7590 14024 7642
rect 14076 7590 14088 7642
rect 14140 7590 14152 7642
rect 14204 7590 14216 7642
rect 14268 7590 17060 7642
rect 17112 7590 17124 7642
rect 17176 7590 17188 7642
rect 17240 7590 17252 7642
rect 17304 7590 17316 7642
rect 17368 7590 18860 7642
rect 0 7568 18860 7590
rect 1302 7488 1308 7540
rect 1360 7528 1366 7540
rect 2133 7531 2191 7537
rect 2133 7528 2145 7531
rect 1360 7500 2145 7528
rect 1360 7488 1366 7500
rect 2133 7497 2145 7500
rect 2179 7497 2191 7531
rect 5537 7531 5595 7537
rect 2133 7491 2191 7497
rect 3988 7500 5396 7528
rect 1946 7460 1952 7472
rect 1907 7432 1952 7460
rect 1946 7420 1952 7432
rect 2004 7420 2010 7472
rect 3786 7420 3792 7472
rect 3844 7460 3850 7472
rect 3881 7463 3939 7469
rect 3881 7460 3893 7463
rect 3844 7432 3893 7460
rect 3844 7420 3850 7432
rect 3881 7429 3893 7432
rect 3927 7429 3939 7463
rect 3881 7423 3939 7429
rect 2038 7392 2044 7404
rect 1999 7364 2044 7392
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 2130 7352 2136 7404
rect 2188 7392 2194 7404
rect 2188 7364 2233 7392
rect 2188 7352 2194 7364
rect 2314 7352 2320 7404
rect 2372 7392 2378 7404
rect 2372 7364 2417 7392
rect 2372 7352 2378 7364
rect 2498 7352 2504 7404
rect 2556 7392 2562 7404
rect 2685 7395 2743 7401
rect 2685 7392 2697 7395
rect 2556 7364 2697 7392
rect 2556 7352 2562 7364
rect 2685 7361 2697 7364
rect 2731 7361 2743 7395
rect 3988 7392 4016 7500
rect 4062 7392 4068 7404
rect 3975 7364 4068 7392
rect 2685 7355 2743 7361
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7392 4307 7395
rect 4338 7392 4344 7404
rect 4295 7364 4344 7392
rect 4295 7361 4307 7364
rect 4249 7355 4307 7361
rect 2590 7324 2596 7336
rect 2551 7296 2596 7324
rect 2590 7284 2596 7296
rect 2648 7284 2654 7336
rect 3878 7284 3884 7336
rect 3936 7324 3942 7336
rect 4172 7324 4200 7355
rect 4338 7352 4344 7364
rect 4396 7352 4402 7404
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7361 4491 7395
rect 4890 7392 4896 7404
rect 4851 7364 4896 7392
rect 4433 7355 4491 7361
rect 4448 7324 4476 7355
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 5056 7401 5114 7407
rect 5368 7404 5396 7500
rect 5537 7497 5549 7531
rect 5583 7528 5595 7531
rect 5626 7528 5632 7540
rect 5583 7500 5632 7528
rect 5583 7497 5595 7500
rect 5537 7491 5595 7497
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 7469 7531 7527 7537
rect 7469 7528 7481 7531
rect 7340 7500 7481 7528
rect 7340 7488 7346 7500
rect 7469 7497 7481 7500
rect 7515 7497 7527 7531
rect 8478 7528 8484 7540
rect 8439 7500 8484 7528
rect 7469 7491 7527 7497
rect 8478 7488 8484 7500
rect 8536 7488 8542 7540
rect 8846 7488 8852 7540
rect 8904 7488 8910 7540
rect 8938 7488 8944 7540
rect 8996 7528 9002 7540
rect 11238 7528 11244 7540
rect 8996 7500 11244 7528
rect 8996 7488 9002 7500
rect 11238 7488 11244 7500
rect 11296 7488 11302 7540
rect 12066 7488 12072 7540
rect 12124 7528 12130 7540
rect 17037 7531 17095 7537
rect 17037 7528 17049 7531
rect 12124 7500 12664 7528
rect 12124 7488 12130 7500
rect 7377 7463 7435 7469
rect 7377 7460 7389 7463
rect 5920 7432 7389 7460
rect 5920 7404 5948 7432
rect 7377 7429 7389 7432
rect 7423 7429 7435 7463
rect 7650 7460 7656 7472
rect 7377 7423 7435 7429
rect 7484 7432 7656 7460
rect 5056 7398 5068 7401
rect 5000 7370 5068 7398
rect 3936 7296 4200 7324
rect 4264 7296 4476 7324
rect 3936 7284 3942 7296
rect 4157 7259 4215 7265
rect 4157 7225 4169 7259
rect 4203 7256 4215 7259
rect 4264 7256 4292 7296
rect 4798 7284 4804 7336
rect 4856 7324 4862 7336
rect 5000 7324 5028 7370
rect 5056 7367 5068 7370
rect 5102 7367 5114 7401
rect 5056 7361 5114 7367
rect 5166 7352 5172 7404
rect 5224 7395 5230 7404
rect 5350 7401 5356 7404
rect 5307 7395 5356 7401
rect 5224 7367 5266 7395
rect 5224 7352 5230 7367
rect 5307 7361 5319 7395
rect 5353 7361 5356 7395
rect 5307 7355 5356 7361
rect 5350 7352 5356 7355
rect 5408 7392 5414 7404
rect 5718 7392 5724 7404
rect 5408 7364 5724 7392
rect 5408 7352 5414 7364
rect 5718 7352 5724 7364
rect 5776 7352 5782 7404
rect 5902 7392 5908 7404
rect 5863 7364 5908 7392
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 6089 7395 6147 7401
rect 6089 7361 6101 7395
rect 6135 7361 6147 7395
rect 6917 7395 6975 7401
rect 6917 7392 6929 7395
rect 6089 7355 6147 7361
rect 6748 7364 6929 7392
rect 4856 7296 5028 7324
rect 4856 7284 4862 7296
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 5994 7324 6000 7336
rect 5592 7296 6000 7324
rect 5592 7284 5598 7296
rect 5994 7284 6000 7296
rect 6052 7324 6058 7336
rect 6104 7324 6132 7355
rect 6052 7296 6132 7324
rect 6457 7327 6515 7333
rect 6052 7284 6058 7296
rect 6457 7293 6469 7327
rect 6503 7324 6515 7327
rect 6546 7324 6552 7336
rect 6503 7296 6552 7324
rect 6503 7293 6515 7296
rect 6457 7287 6515 7293
rect 6546 7284 6552 7296
rect 6604 7284 6610 7336
rect 4203 7228 4292 7256
rect 6089 7259 6147 7265
rect 4203 7225 4215 7228
rect 4157 7219 4215 7225
rect 6089 7225 6101 7259
rect 6135 7256 6147 7259
rect 6748 7256 6776 7364
rect 6917 7361 6929 7364
rect 6963 7392 6975 7395
rect 7484 7392 7512 7432
rect 7650 7420 7656 7432
rect 7708 7460 7714 7472
rect 8110 7460 8116 7472
rect 7708 7432 8116 7460
rect 7708 7420 7714 7432
rect 8110 7420 8116 7432
rect 8168 7420 8174 7472
rect 8864 7460 8892 7488
rect 11333 7463 11391 7469
rect 11333 7460 11345 7463
rect 8864 7432 11345 7460
rect 11333 7429 11345 7432
rect 11379 7429 11391 7463
rect 12529 7463 12587 7469
rect 12529 7460 12541 7463
rect 11333 7423 11391 7429
rect 12360 7432 12541 7460
rect 6963 7364 7512 7392
rect 8021 7395 8079 7401
rect 6963 7361 6975 7364
rect 6917 7355 6975 7361
rect 8021 7361 8033 7395
rect 8067 7392 8079 7395
rect 8849 7395 8907 7401
rect 8067 7364 8800 7392
rect 8067 7361 8079 7364
rect 8021 7355 8079 7361
rect 6825 7327 6883 7333
rect 6825 7293 6837 7327
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 6135 7228 6776 7256
rect 6840 7256 6868 7287
rect 7006 7284 7012 7336
rect 7064 7324 7070 7336
rect 7374 7324 7380 7336
rect 7064 7296 7380 7324
rect 7064 7284 7070 7296
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8202 7324 8208 7336
rect 8159 7296 8208 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 8297 7327 8355 7333
rect 8297 7293 8309 7327
rect 8343 7293 8355 7327
rect 8297 7287 8355 7293
rect 7653 7259 7711 7265
rect 7653 7256 7665 7259
rect 6840 7228 7665 7256
rect 6135 7225 6147 7228
rect 6089 7219 6147 7225
rect 7653 7225 7665 7228
rect 7699 7225 7711 7259
rect 8312 7256 8340 7287
rect 7653 7219 7711 7225
rect 8128 7228 8340 7256
rect 8772 7256 8800 7364
rect 8849 7361 8861 7395
rect 8895 7392 8907 7395
rect 9122 7392 9128 7404
rect 8895 7364 9128 7392
rect 8895 7361 8907 7364
rect 8849 7355 8907 7361
rect 9122 7352 9128 7364
rect 9180 7352 9186 7404
rect 10413 7395 10471 7401
rect 10413 7361 10425 7395
rect 10459 7392 10471 7395
rect 10873 7395 10931 7401
rect 10873 7392 10885 7395
rect 10459 7364 10885 7392
rect 10459 7361 10471 7364
rect 10413 7355 10471 7361
rect 10873 7361 10885 7364
rect 10919 7361 10931 7395
rect 11054 7392 11060 7404
rect 11015 7364 11060 7392
rect 10873 7355 10931 7361
rect 11054 7352 11060 7364
rect 11112 7392 11118 7404
rect 11698 7392 11704 7404
rect 11112 7364 11704 7392
rect 11112 7352 11118 7364
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 12158 7392 12164 7404
rect 11808 7364 12164 7392
rect 8938 7324 8944 7336
rect 8899 7296 8944 7324
rect 8938 7284 8944 7296
rect 8996 7284 9002 7336
rect 9030 7284 9036 7336
rect 9088 7324 9094 7336
rect 10318 7324 10324 7336
rect 9088 7296 10324 7324
rect 9088 7284 9094 7296
rect 10318 7284 10324 7296
rect 10376 7284 10382 7336
rect 10505 7327 10563 7333
rect 10505 7293 10517 7327
rect 10551 7293 10563 7327
rect 10505 7287 10563 7293
rect 10689 7327 10747 7333
rect 10689 7293 10701 7327
rect 10735 7324 10747 7327
rect 11422 7324 11428 7336
rect 10735 7296 11428 7324
rect 10735 7293 10747 7296
rect 10689 7287 10747 7293
rect 10045 7259 10103 7265
rect 10045 7256 10057 7259
rect 8772 7228 10057 7256
rect 2958 7148 2964 7200
rect 3016 7188 3022 7200
rect 3053 7191 3111 7197
rect 3053 7188 3065 7191
rect 3016 7160 3065 7188
rect 3016 7148 3022 7160
rect 3053 7157 3065 7160
rect 3099 7157 3111 7191
rect 4246 7188 4252 7200
rect 4207 7160 4252 7188
rect 3053 7151 3111 7157
rect 4246 7148 4252 7160
rect 4304 7148 4310 7200
rect 7101 7191 7159 7197
rect 7101 7157 7113 7191
rect 7147 7188 7159 7191
rect 7374 7188 7380 7200
rect 7147 7160 7380 7188
rect 7147 7157 7159 7160
rect 7101 7151 7159 7157
rect 7374 7148 7380 7160
rect 7432 7148 7438 7200
rect 7558 7148 7564 7200
rect 7616 7188 7622 7200
rect 8128 7188 8156 7228
rect 10045 7225 10057 7228
rect 10091 7225 10103 7259
rect 10520 7256 10548 7287
rect 11422 7284 11428 7296
rect 11480 7284 11486 7336
rect 10778 7256 10784 7268
rect 10520 7228 10784 7256
rect 10045 7219 10103 7225
rect 10778 7216 10784 7228
rect 10836 7256 10842 7268
rect 11808 7256 11836 7364
rect 12158 7352 12164 7364
rect 12216 7352 12222 7404
rect 12360 7401 12388 7432
rect 12529 7429 12541 7432
rect 12575 7429 12587 7463
rect 12529 7423 12587 7429
rect 12636 7401 12664 7500
rect 13924 7500 17049 7528
rect 12345 7395 12403 7401
rect 12345 7361 12357 7395
rect 12391 7361 12403 7395
rect 12345 7355 12403 7361
rect 12437 7395 12495 7401
rect 12437 7361 12449 7395
rect 12483 7361 12495 7395
rect 12437 7355 12495 7361
rect 12621 7395 12679 7401
rect 12621 7361 12633 7395
rect 12667 7392 12679 7395
rect 12894 7392 12900 7404
rect 12667 7364 12900 7392
rect 12667 7361 12679 7364
rect 12621 7355 12679 7361
rect 12069 7327 12127 7333
rect 12069 7293 12081 7327
rect 12115 7324 12127 7327
rect 12250 7324 12256 7336
rect 12115 7296 12256 7324
rect 12115 7293 12127 7296
rect 12069 7287 12127 7293
rect 12250 7284 12256 7296
rect 12308 7284 12314 7336
rect 12452 7324 12480 7355
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 13541 7395 13599 7401
rect 13541 7361 13553 7395
rect 13587 7361 13599 7395
rect 13541 7355 13599 7361
rect 13725 7395 13783 7401
rect 13725 7361 13737 7395
rect 13771 7392 13783 7395
rect 13817 7395 13875 7401
rect 13817 7392 13829 7395
rect 13771 7364 13829 7392
rect 13771 7361 13783 7364
rect 13725 7355 13783 7361
rect 13817 7361 13829 7364
rect 13863 7361 13875 7395
rect 13924 7392 13952 7500
rect 17037 7497 17049 7500
rect 17083 7497 17095 7531
rect 17037 7491 17095 7497
rect 14182 7460 14188 7472
rect 14143 7432 14188 7460
rect 14182 7420 14188 7432
rect 14240 7420 14246 7472
rect 14366 7460 14372 7472
rect 14292 7432 14372 7460
rect 13998 7392 14004 7404
rect 14056 7401 14062 7404
rect 14292 7401 14320 7432
rect 14366 7420 14372 7432
rect 14424 7420 14430 7472
rect 14056 7395 14078 7401
rect 13924 7364 14004 7392
rect 13817 7355 13875 7361
rect 12802 7324 12808 7336
rect 12452 7296 12808 7324
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 10836 7228 11836 7256
rect 13556 7256 13584 7355
rect 13998 7352 14004 7364
rect 14066 7392 14078 7395
rect 14277 7395 14335 7401
rect 14066 7364 14149 7392
rect 14066 7361 14078 7364
rect 14056 7355 14078 7361
rect 14277 7361 14289 7395
rect 14323 7361 14335 7395
rect 14458 7392 14464 7404
rect 14419 7364 14464 7392
rect 14277 7355 14335 7361
rect 14056 7352 14062 7355
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 13633 7327 13691 7333
rect 13633 7293 13645 7327
rect 13679 7324 13691 7327
rect 14829 7327 14887 7333
rect 14829 7324 14841 7327
rect 13679 7296 14841 7324
rect 13679 7293 13691 7296
rect 13633 7287 13691 7293
rect 14829 7293 14841 7296
rect 14875 7293 14887 7327
rect 15856 7324 15884 7446
rect 16255 7395 16313 7401
rect 16255 7361 16267 7395
rect 16301 7392 16313 7395
rect 16942 7392 16948 7404
rect 16301 7364 16948 7392
rect 16301 7361 16313 7364
rect 16255 7355 16313 7361
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 15856 7296 16344 7324
rect 14829 7287 14887 7293
rect 14090 7256 14096 7268
rect 13556 7228 14096 7256
rect 10836 7216 10842 7228
rect 14090 7216 14096 7228
rect 14148 7216 14154 7268
rect 16316 7200 16344 7296
rect 9030 7188 9036 7200
rect 7616 7160 9036 7188
rect 7616 7148 7622 7160
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 11422 7188 11428 7200
rect 11383 7160 11428 7188
rect 11422 7148 11428 7160
rect 11480 7148 11486 7200
rect 12158 7188 12164 7200
rect 12119 7160 12164 7188
rect 12158 7148 12164 7160
rect 12216 7148 12222 7200
rect 12250 7148 12256 7200
rect 12308 7188 12314 7200
rect 12308 7160 12353 7188
rect 12308 7148 12314 7160
rect 16298 7148 16304 7200
rect 16356 7188 16362 7200
rect 16393 7191 16451 7197
rect 16393 7188 16405 7191
rect 16356 7160 16405 7188
rect 16356 7148 16362 7160
rect 16393 7157 16405 7160
rect 16439 7157 16451 7191
rect 16393 7151 16451 7157
rect 0 7098 18860 7120
rect 0 7046 3110 7098
rect 3162 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 3302 7098
rect 3354 7046 3366 7098
rect 3418 7046 6210 7098
rect 6262 7046 6274 7098
rect 6326 7046 6338 7098
rect 6390 7046 6402 7098
rect 6454 7046 6466 7098
rect 6518 7046 9310 7098
rect 9362 7046 9374 7098
rect 9426 7046 9438 7098
rect 9490 7046 9502 7098
rect 9554 7046 9566 7098
rect 9618 7046 12410 7098
rect 12462 7046 12474 7098
rect 12526 7046 12538 7098
rect 12590 7046 12602 7098
rect 12654 7046 12666 7098
rect 12718 7046 15510 7098
rect 15562 7046 15574 7098
rect 15626 7046 15638 7098
rect 15690 7046 15702 7098
rect 15754 7046 15766 7098
rect 15818 7046 18860 7098
rect 0 7024 18860 7046
rect 3878 6944 3884 6996
rect 3936 6944 3942 6996
rect 6365 6987 6423 6993
rect 6365 6953 6377 6987
rect 6411 6984 6423 6987
rect 6546 6984 6552 6996
rect 6411 6956 6552 6984
rect 6411 6953 6423 6956
rect 6365 6947 6423 6953
rect 6546 6944 6552 6956
rect 6604 6944 6610 6996
rect 7374 6944 7380 6996
rect 7432 6984 7438 6996
rect 8033 6987 8091 6993
rect 8033 6984 8045 6987
rect 7432 6956 8045 6984
rect 7432 6944 7438 6956
rect 8033 6953 8045 6956
rect 8079 6953 8091 6987
rect 8033 6947 8091 6953
rect 8202 6944 8208 6996
rect 8260 6984 8266 6996
rect 10778 6984 10784 6996
rect 8260 6956 10784 6984
rect 8260 6944 8266 6956
rect 10778 6944 10784 6956
rect 10836 6944 10842 6996
rect 12250 6944 12256 6996
rect 12308 6984 12314 6996
rect 12345 6987 12403 6993
rect 12345 6984 12357 6987
rect 12308 6956 12357 6984
rect 12308 6944 12314 6956
rect 12345 6953 12357 6956
rect 12391 6953 12403 6987
rect 14090 6984 14096 6996
rect 14051 6956 14096 6984
rect 12345 6947 12403 6953
rect 14090 6944 14096 6956
rect 14148 6944 14154 6996
rect 3896 6916 3924 6944
rect 4430 6916 4436 6928
rect 3896 6888 4436 6916
rect 4430 6876 4436 6888
rect 4488 6916 4494 6928
rect 5166 6916 5172 6928
rect 4488 6888 5172 6916
rect 4488 6876 4494 6888
rect 2225 6851 2283 6857
rect 2225 6817 2237 6851
rect 2271 6848 2283 6851
rect 2498 6848 2504 6860
rect 2271 6820 2504 6848
rect 2271 6817 2283 6820
rect 2225 6811 2283 6817
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 3329 6851 3387 6857
rect 3329 6817 3341 6851
rect 3375 6848 3387 6851
rect 3694 6848 3700 6860
rect 3375 6820 3700 6848
rect 3375 6817 3387 6820
rect 3329 6811 3387 6817
rect 3694 6808 3700 6820
rect 3752 6808 3758 6860
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 3970 6848 3976 6860
rect 3927 6820 3976 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 3970 6808 3976 6820
rect 4028 6808 4034 6860
rect 4890 6848 4896 6860
rect 4172 6820 4896 6848
rect 937 6783 995 6789
rect 937 6749 949 6783
rect 983 6749 995 6783
rect 937 6743 995 6749
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6780 2007 6783
rect 2406 6780 2412 6792
rect 1995 6752 2412 6780
rect 1995 6749 2007 6752
rect 1949 6743 2007 6749
rect 566 6604 572 6656
rect 624 6644 630 6656
rect 753 6647 811 6653
rect 753 6644 765 6647
rect 624 6616 765 6644
rect 624 6604 630 6616
rect 753 6613 765 6616
rect 799 6613 811 6647
rect 952 6644 980 6743
rect 2406 6740 2412 6752
rect 2464 6740 2470 6792
rect 2593 6783 2651 6789
rect 2593 6749 2605 6783
rect 2639 6780 2651 6783
rect 2866 6780 2872 6792
rect 2639 6752 2872 6780
rect 2639 6749 2651 6752
rect 2593 6743 2651 6749
rect 2866 6740 2872 6752
rect 2924 6740 2930 6792
rect 4172 6789 4200 6820
rect 4890 6808 4896 6820
rect 4948 6808 4954 6860
rect 5000 6789 5028 6888
rect 5166 6876 5172 6888
rect 5224 6876 5230 6928
rect 5905 6919 5963 6925
rect 5905 6885 5917 6919
rect 5951 6916 5963 6919
rect 7006 6916 7012 6928
rect 5951 6888 7012 6916
rect 5951 6885 5963 6888
rect 5905 6879 5963 6885
rect 7006 6876 7012 6888
rect 7064 6876 7070 6928
rect 14274 6916 14280 6928
rect 14108 6888 14280 6916
rect 7282 6848 7288 6860
rect 6380 6820 7288 6848
rect 4157 6783 4215 6789
rect 4157 6780 4169 6783
rect 3068 6752 4169 6780
rect 2501 6715 2559 6721
rect 2501 6681 2513 6715
rect 2547 6712 2559 6715
rect 3068 6712 3096 6752
rect 4157 6749 4169 6752
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6780 5319 6783
rect 5350 6780 5356 6792
rect 5307 6752 5356 6780
rect 5307 6749 5319 6752
rect 5261 6743 5319 6749
rect 2547 6684 3096 6712
rect 3145 6715 3203 6721
rect 2547 6681 2559 6684
rect 2501 6675 2559 6681
rect 3145 6681 3157 6715
rect 3191 6712 3203 6715
rect 4338 6712 4344 6724
rect 3191 6684 4344 6712
rect 3191 6681 3203 6684
rect 3145 6675 3203 6681
rect 4338 6672 4344 6684
rect 4396 6672 4402 6724
rect 4522 6672 4528 6724
rect 4580 6712 4586 6724
rect 4632 6712 4660 6743
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 5994 6740 6000 6792
rect 6052 6780 6058 6792
rect 6380 6789 6408 6820
rect 7282 6808 7288 6820
rect 7340 6808 7346 6860
rect 10873 6851 10931 6857
rect 10873 6848 10885 6851
rect 8588 6820 10885 6848
rect 8588 6789 8616 6820
rect 10873 6817 10885 6820
rect 10919 6817 10931 6851
rect 12802 6848 12808 6860
rect 10873 6811 10931 6817
rect 12544 6820 12808 6848
rect 6273 6783 6331 6789
rect 6273 6780 6285 6783
rect 6052 6752 6285 6780
rect 6052 6740 6058 6752
rect 6273 6749 6285 6752
rect 6319 6749 6331 6783
rect 6273 6743 6331 6749
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 8297 6783 8355 6789
rect 8297 6749 8309 6783
rect 8343 6780 8355 6783
rect 8573 6783 8631 6789
rect 8573 6780 8585 6783
rect 8343 6752 8585 6780
rect 8343 6749 8355 6752
rect 8297 6743 8355 6749
rect 8573 6749 8585 6752
rect 8619 6749 8631 6783
rect 8573 6743 8631 6749
rect 10318 6740 10324 6792
rect 10376 6780 10382 6792
rect 10597 6783 10655 6789
rect 10597 6780 10609 6783
rect 10376 6752 10609 6780
rect 10376 6740 10382 6752
rect 10597 6749 10609 6752
rect 10643 6749 10655 6783
rect 10888 6780 10916 6811
rect 11422 6780 11428 6792
rect 10888 6752 11428 6780
rect 10597 6743 10655 6749
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 12544 6789 12572 6820
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 12529 6783 12587 6789
rect 12529 6749 12541 6783
rect 12575 6749 12587 6783
rect 12529 6743 12587 6749
rect 12713 6783 12771 6789
rect 12713 6749 12725 6783
rect 12759 6780 12771 6783
rect 12894 6780 12900 6792
rect 12759 6752 12900 6780
rect 12759 6749 12771 6752
rect 12713 6743 12771 6749
rect 4798 6712 4804 6724
rect 4580 6684 4804 6712
rect 4580 6672 4586 6684
rect 4798 6672 4804 6684
rect 4856 6712 4862 6724
rect 5718 6712 5724 6724
rect 4856 6684 5724 6712
rect 4856 6672 4862 6684
rect 5718 6672 5724 6684
rect 5776 6672 5782 6724
rect 6089 6715 6147 6721
rect 6089 6681 6101 6715
rect 6135 6712 6147 6715
rect 6135 6684 6592 6712
rect 6135 6681 6147 6684
rect 6089 6675 6147 6681
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 952 6616 1593 6644
rect 753 6607 811 6613
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 2041 6647 2099 6653
rect 2041 6613 2053 6647
rect 2087 6644 2099 6647
rect 2685 6647 2743 6653
rect 2685 6644 2697 6647
rect 2087 6616 2697 6644
rect 2087 6613 2099 6616
rect 2041 6607 2099 6613
rect 2685 6613 2697 6616
rect 2731 6613 2743 6647
rect 2685 6607 2743 6613
rect 2958 6604 2964 6656
rect 3016 6644 3022 6656
rect 6564 6653 6592 6684
rect 7006 6672 7012 6724
rect 7064 6672 7070 6724
rect 8846 6712 8852 6724
rect 8807 6684 8852 6712
rect 8846 6672 8852 6684
rect 8904 6672 8910 6724
rect 10686 6712 10692 6724
rect 10074 6684 10692 6712
rect 10686 6672 10692 6684
rect 10744 6672 10750 6724
rect 10962 6712 10968 6724
rect 10796 6684 10968 6712
rect 3053 6647 3111 6653
rect 3053 6644 3065 6647
rect 3016 6616 3065 6644
rect 3016 6604 3022 6616
rect 3053 6613 3065 6616
rect 3099 6613 3111 6647
rect 3053 6607 3111 6613
rect 6549 6647 6607 6653
rect 6549 6613 6561 6647
rect 6595 6644 6607 6647
rect 8754 6644 8760 6656
rect 6595 6616 8760 6644
rect 6595 6613 6607 6616
rect 6549 6607 6607 6613
rect 8754 6604 8760 6616
rect 8812 6644 8818 6656
rect 10796 6644 10824 6684
rect 10962 6672 10968 6684
rect 11020 6672 11026 6724
rect 11140 6715 11198 6721
rect 11140 6681 11152 6715
rect 11186 6712 11198 6715
rect 12728 6712 12756 6743
rect 12894 6740 12900 6752
rect 12952 6780 12958 6792
rect 13538 6780 13544 6792
rect 12952 6752 13544 6780
rect 12952 6740 12958 6752
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 14108 6789 14136 6888
rect 14274 6876 14280 6888
rect 14332 6916 14338 6928
rect 14332 6888 14504 6916
rect 14332 6876 14338 6888
rect 14366 6808 14372 6860
rect 14424 6808 14430 6860
rect 14476 6848 14504 6888
rect 15381 6851 15439 6857
rect 15381 6848 15393 6851
rect 14476 6820 15393 6848
rect 15381 6817 15393 6820
rect 15427 6848 15439 6851
rect 16942 6848 16948 6860
rect 15427 6820 16948 6848
rect 15427 6817 15439 6820
rect 15381 6811 15439 6817
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 17862 6848 17868 6860
rect 17823 6820 17868 6848
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 14093 6783 14151 6789
rect 14093 6749 14105 6783
rect 14139 6749 14151 6783
rect 14093 6743 14151 6749
rect 14185 6783 14243 6789
rect 14185 6749 14197 6783
rect 14231 6780 14243 6783
rect 14384 6780 14412 6808
rect 15749 6783 15807 6789
rect 15749 6780 15761 6783
rect 14231 6752 14412 6780
rect 15396 6752 15761 6780
rect 14231 6749 14243 6752
rect 14185 6743 14243 6749
rect 11186 6684 12756 6712
rect 11186 6681 11198 6684
rect 11140 6675 11198 6681
rect 13998 6672 14004 6724
rect 14056 6712 14062 6724
rect 14369 6715 14427 6721
rect 14369 6712 14381 6715
rect 14056 6684 14381 6712
rect 14056 6672 14062 6684
rect 14369 6681 14381 6684
rect 14415 6681 14427 6715
rect 14369 6675 14427 6681
rect 14461 6715 14519 6721
rect 14461 6681 14473 6715
rect 14507 6712 14519 6715
rect 15396 6712 15424 6752
rect 15749 6749 15761 6752
rect 15795 6780 15807 6783
rect 18233 6783 18291 6789
rect 15795 6752 16344 6780
rect 15795 6749 15807 6752
rect 15749 6743 15807 6749
rect 16316 6724 16344 6752
rect 18233 6749 18245 6783
rect 18279 6780 18291 6783
rect 18506 6780 18512 6792
rect 18279 6752 18512 6780
rect 18279 6749 18291 6752
rect 18233 6743 18291 6749
rect 18506 6740 18512 6752
rect 18564 6740 18570 6792
rect 15838 6712 15844 6724
rect 14507 6684 15424 6712
rect 15799 6684 15844 6712
rect 14507 6681 14519 6684
rect 14461 6675 14519 6681
rect 15838 6672 15844 6684
rect 15896 6672 15902 6724
rect 16298 6672 16304 6724
rect 16356 6712 16362 6724
rect 16356 6684 16422 6712
rect 16356 6672 16362 6684
rect 17494 6672 17500 6724
rect 17552 6712 17558 6724
rect 17589 6715 17647 6721
rect 17589 6712 17601 6715
rect 17552 6684 17601 6712
rect 17552 6672 17558 6684
rect 17589 6681 17601 6684
rect 17635 6681 17647 6715
rect 17589 6675 17647 6681
rect 8812 6616 10824 6644
rect 12253 6647 12311 6653
rect 8812 6604 8818 6616
rect 12253 6613 12265 6647
rect 12299 6644 12311 6647
rect 12802 6644 12808 6656
rect 12299 6616 12808 6644
rect 12299 6613 12311 6616
rect 12253 6607 12311 6613
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 14550 6604 14556 6656
rect 14608 6644 14614 6656
rect 14737 6647 14795 6653
rect 14737 6644 14749 6647
rect 14608 6616 14749 6644
rect 14608 6604 14614 6616
rect 14737 6613 14749 6616
rect 14783 6613 14795 6647
rect 15102 6644 15108 6656
rect 15063 6616 15108 6644
rect 14737 6607 14795 6613
rect 15102 6604 15108 6616
rect 15160 6604 15166 6656
rect 15197 6647 15255 6653
rect 15197 6613 15209 6647
rect 15243 6644 15255 6647
rect 15930 6644 15936 6656
rect 15243 6616 15936 6644
rect 15243 6613 15255 6616
rect 15197 6607 15255 6613
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 18322 6644 18328 6656
rect 18283 6616 18328 6644
rect 18322 6604 18328 6616
rect 18380 6604 18386 6656
rect 0 6554 18860 6576
rect 0 6502 4660 6554
rect 4712 6502 4724 6554
rect 4776 6502 4788 6554
rect 4840 6502 4852 6554
rect 4904 6502 4916 6554
rect 4968 6502 7760 6554
rect 7812 6502 7824 6554
rect 7876 6502 7888 6554
rect 7940 6502 7952 6554
rect 8004 6502 8016 6554
rect 8068 6502 10860 6554
rect 10912 6502 10924 6554
rect 10976 6502 10988 6554
rect 11040 6502 11052 6554
rect 11104 6502 11116 6554
rect 11168 6502 13960 6554
rect 14012 6502 14024 6554
rect 14076 6502 14088 6554
rect 14140 6502 14152 6554
rect 14204 6502 14216 6554
rect 14268 6502 17060 6554
rect 17112 6502 17124 6554
rect 17176 6502 17188 6554
rect 17240 6502 17252 6554
rect 17304 6502 17316 6554
rect 17368 6502 18860 6554
rect 0 6480 18860 6502
rect 2041 6443 2099 6449
rect 2041 6409 2053 6443
rect 2087 6440 2099 6443
rect 2406 6440 2412 6452
rect 2087 6412 2412 6440
rect 2087 6409 2099 6412
rect 2041 6403 2099 6409
rect 2406 6400 2412 6412
rect 2464 6400 2470 6452
rect 2590 6440 2596 6452
rect 2551 6412 2596 6440
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 3513 6443 3571 6449
rect 3513 6409 3525 6443
rect 3559 6440 3571 6443
rect 4246 6440 4252 6452
rect 3559 6412 4252 6440
rect 3559 6409 3571 6412
rect 3513 6403 3571 6409
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 7469 6443 7527 6449
rect 7469 6409 7481 6443
rect 7515 6440 7527 6443
rect 8846 6440 8852 6452
rect 7515 6412 8852 6440
rect 7515 6409 7527 6412
rect 7469 6403 7527 6409
rect 8846 6400 8852 6412
rect 8904 6400 8910 6452
rect 12713 6443 12771 6449
rect 12713 6409 12725 6443
rect 12759 6440 12771 6443
rect 13449 6443 13507 6449
rect 13449 6440 13461 6443
rect 12759 6412 13461 6440
rect 12759 6409 12771 6412
rect 12713 6403 12771 6409
rect 13449 6409 13461 6412
rect 13495 6409 13507 6443
rect 13449 6403 13507 6409
rect 13538 6400 13544 6452
rect 13596 6440 13602 6452
rect 13909 6443 13967 6449
rect 13909 6440 13921 6443
rect 13596 6412 13921 6440
rect 13596 6400 13602 6412
rect 13909 6409 13921 6412
rect 13955 6409 13967 6443
rect 13909 6403 13967 6409
rect 14737 6443 14795 6449
rect 14737 6409 14749 6443
rect 14783 6440 14795 6443
rect 15102 6440 15108 6452
rect 14783 6412 15108 6440
rect 14783 6409 14795 6412
rect 14737 6403 14795 6409
rect 15102 6400 15108 6412
rect 15160 6400 15166 6452
rect 16206 6440 16212 6452
rect 15212 6412 16212 6440
rect 566 6372 572 6384
rect 527 6344 572 6372
rect 566 6332 572 6344
rect 624 6332 630 6384
rect 2222 6372 2228 6384
rect 1794 6344 2228 6372
rect 2222 6332 2228 6344
rect 2280 6332 2286 6384
rect 3973 6375 4031 6381
rect 3973 6341 3985 6375
rect 4019 6372 4031 6375
rect 4338 6372 4344 6384
rect 4019 6344 4344 6372
rect 4019 6341 4031 6344
rect 3973 6335 4031 6341
rect 4338 6332 4344 6344
rect 4396 6332 4402 6384
rect 5629 6375 5687 6381
rect 5629 6341 5641 6375
rect 5675 6372 5687 6375
rect 12158 6372 12164 6384
rect 5675 6344 7696 6372
rect 5675 6341 5687 6344
rect 5629 6335 5687 6341
rect 7668 6316 7696 6344
rect 7852 6344 12164 6372
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6273 2559 6307
rect 2682 6304 2688 6316
rect 2643 6276 2688 6304
rect 2501 6267 2559 6273
rect 290 6236 296 6248
rect 251 6208 296 6236
rect 290 6196 296 6208
rect 348 6196 354 6248
rect 2516 6236 2544 6267
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3421 6307 3479 6313
rect 3421 6304 3433 6307
rect 2832 6276 3433 6304
rect 2832 6264 2838 6276
rect 3421 6273 3433 6276
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 4157 6307 4215 6313
rect 4157 6304 4169 6307
rect 4120 6276 4169 6304
rect 4120 6264 4126 6276
rect 4157 6273 4169 6276
rect 4203 6273 4215 6307
rect 5721 6307 5779 6313
rect 5721 6304 5733 6307
rect 4157 6267 4215 6273
rect 4356 6276 5733 6304
rect 2866 6236 2872 6248
rect 2516 6208 2872 6236
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 3694 6236 3700 6248
rect 3655 6208 3700 6236
rect 3694 6196 3700 6208
rect 3752 6236 3758 6248
rect 4356 6236 4384 6276
rect 5721 6273 5733 6276
rect 5767 6304 5779 6307
rect 5767 6276 5948 6304
rect 5767 6273 5779 6276
rect 5721 6267 5779 6273
rect 3752 6208 4384 6236
rect 4433 6239 4491 6245
rect 3752 6196 3758 6208
rect 4433 6205 4445 6239
rect 4479 6236 4491 6239
rect 4522 6236 4528 6248
rect 4479 6208 4528 6236
rect 4479 6205 4491 6208
rect 4433 6199 4491 6205
rect 4522 6196 4528 6208
rect 4580 6196 4586 6248
rect 5813 6239 5871 6245
rect 5813 6205 5825 6239
rect 5859 6205 5871 6239
rect 5813 6199 5871 6205
rect 2498 6128 2504 6180
rect 2556 6168 2562 6180
rect 5261 6171 5319 6177
rect 5261 6168 5273 6171
rect 2556 6140 5273 6168
rect 2556 6128 2562 6140
rect 5261 6137 5273 6140
rect 5307 6168 5319 6171
rect 5442 6168 5448 6180
rect 5307 6140 5448 6168
rect 5307 6137 5319 6140
rect 5261 6131 5319 6137
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 5626 6128 5632 6180
rect 5684 6168 5690 6180
rect 5828 6168 5856 6199
rect 5684 6140 5856 6168
rect 5920 6168 5948 6276
rect 5994 6264 6000 6316
rect 6052 6304 6058 6316
rect 6457 6307 6515 6313
rect 6457 6304 6469 6307
rect 6052 6276 6469 6304
rect 6052 6264 6058 6276
rect 6457 6273 6469 6276
rect 6503 6273 6515 6307
rect 7650 6304 7656 6316
rect 7611 6276 7656 6304
rect 6457 6267 6515 6273
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 7852 6313 7880 6344
rect 12158 6332 12164 6344
rect 12216 6332 12222 6384
rect 15212 6372 15240 6412
rect 16206 6400 16212 6412
rect 16264 6400 16270 6452
rect 16942 6440 16948 6452
rect 16903 6412 16948 6440
rect 16942 6400 16948 6412
rect 17000 6400 17006 6452
rect 14752 6344 15240 6372
rect 7837 6307 7895 6313
rect 7837 6273 7849 6307
rect 7883 6273 7895 6307
rect 8018 6304 8024 6316
rect 7979 6276 8024 6304
rect 7837 6267 7895 6273
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6273 8631 6307
rect 8573 6267 8631 6273
rect 11885 6307 11943 6313
rect 11885 6273 11897 6307
rect 11931 6304 11943 6307
rect 13814 6304 13820 6316
rect 11931 6276 12388 6304
rect 13775 6276 13820 6304
rect 11931 6273 11943 6276
rect 11885 6267 11943 6273
rect 6546 6236 6552 6248
rect 6507 6208 6552 6236
rect 6546 6196 6552 6208
rect 6604 6196 6610 6248
rect 6641 6239 6699 6245
rect 6641 6205 6653 6239
rect 6687 6236 6699 6239
rect 7558 6236 7564 6248
rect 6687 6208 7564 6236
rect 6687 6205 6699 6208
rect 6641 6199 6699 6205
rect 6656 6168 6684 6199
rect 7558 6196 7564 6208
rect 7616 6196 7622 6248
rect 7929 6239 7987 6245
rect 7929 6205 7941 6239
rect 7975 6236 7987 6239
rect 8386 6236 8392 6248
rect 7975 6208 8392 6236
rect 7975 6205 7987 6208
rect 7929 6199 7987 6205
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 8588 6168 8616 6267
rect 8938 6168 8944 6180
rect 5920 6140 6684 6168
rect 8312 6140 8616 6168
rect 8680 6140 8944 6168
rect 5684 6128 5690 6140
rect 8312 6112 8340 6140
rect 8680 6112 8708 6140
rect 8938 6128 8944 6140
rect 8996 6128 9002 6180
rect 12360 6177 12388 6276
rect 13814 6264 13820 6276
rect 13872 6264 13878 6316
rect 14642 6264 14648 6316
rect 14700 6304 14706 6316
rect 14752 6313 14780 6344
rect 14737 6307 14795 6313
rect 14737 6304 14749 6307
rect 14700 6276 14749 6304
rect 14700 6264 14706 6276
rect 14737 6273 14749 6276
rect 14783 6273 14795 6307
rect 14737 6267 14795 6273
rect 16298 6264 16304 6316
rect 16356 6264 16362 6316
rect 16482 6264 16488 6316
rect 16540 6304 16546 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16540 6276 16865 6304
rect 16540 6264 16546 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 17313 6307 17371 6313
rect 17313 6273 17325 6307
rect 17359 6273 17371 6307
rect 17313 6267 17371 6273
rect 17681 6307 17739 6313
rect 17681 6273 17693 6307
rect 17727 6273 17739 6307
rect 17681 6267 17739 6273
rect 12802 6236 12808 6248
rect 12763 6208 12808 6236
rect 12802 6196 12808 6208
rect 12860 6196 12866 6248
rect 12989 6239 13047 6245
rect 12989 6205 13001 6239
rect 13035 6205 13047 6239
rect 12989 6199 13047 6205
rect 14093 6239 14151 6245
rect 14093 6205 14105 6239
rect 14139 6236 14151 6239
rect 14366 6236 14372 6248
rect 14139 6208 14372 6236
rect 14139 6205 14151 6208
rect 14093 6199 14151 6205
rect 12345 6171 12403 6177
rect 12345 6137 12357 6171
rect 12391 6137 12403 6171
rect 13004 6168 13032 6199
rect 14366 6196 14372 6208
rect 14424 6196 14430 6248
rect 14458 6196 14464 6248
rect 14516 6236 14522 6248
rect 14921 6239 14979 6245
rect 14921 6236 14933 6239
rect 14516 6208 14933 6236
rect 14516 6196 14522 6208
rect 14921 6205 14933 6208
rect 14967 6205 14979 6239
rect 14921 6199 14979 6205
rect 15197 6239 15255 6245
rect 15197 6205 15209 6239
rect 15243 6236 15255 6239
rect 16574 6236 16580 6248
rect 15243 6208 16580 6236
rect 15243 6205 15255 6208
rect 15197 6199 15255 6205
rect 16574 6196 16580 6208
rect 16632 6196 16638 6248
rect 16669 6239 16727 6245
rect 16669 6205 16681 6239
rect 16715 6236 16727 6239
rect 17328 6236 17356 6267
rect 17402 6236 17408 6248
rect 16715 6208 17408 6236
rect 16715 6205 16727 6208
rect 16669 6199 16727 6205
rect 17402 6196 17408 6208
rect 17460 6196 17466 6248
rect 13004 6140 14320 6168
rect 12345 6131 12403 6137
rect 14292 6112 14320 6140
rect 16206 6128 16212 6180
rect 16264 6168 16270 6180
rect 17696 6168 17724 6267
rect 16264 6140 17724 6168
rect 16264 6128 16270 6140
rect 2222 6100 2228 6112
rect 2183 6072 2228 6100
rect 2222 6060 2228 6072
rect 2280 6060 2286 6112
rect 2958 6060 2964 6112
rect 3016 6100 3022 6112
rect 3053 6103 3111 6109
rect 3053 6100 3065 6103
rect 3016 6072 3065 6100
rect 3016 6060 3022 6072
rect 3053 6069 3065 6072
rect 3099 6069 3111 6103
rect 3053 6063 3111 6069
rect 4341 6103 4399 6109
rect 4341 6069 4353 6103
rect 4387 6100 4399 6103
rect 4430 6100 4436 6112
rect 4387 6072 4436 6100
rect 4387 6069 4399 6072
rect 4341 6063 4399 6069
rect 4430 6060 4436 6072
rect 4488 6060 4494 6112
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 6089 6103 6147 6109
rect 6089 6100 6101 6103
rect 5592 6072 6101 6100
rect 5592 6060 5598 6072
rect 6089 6069 6101 6072
rect 6135 6069 6147 6103
rect 8294 6100 8300 6112
rect 8207 6072 8300 6100
rect 6089 6063 6147 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 8481 6103 8539 6109
rect 8481 6069 8493 6103
rect 8527 6100 8539 6103
rect 8570 6100 8576 6112
rect 8527 6072 8576 6100
rect 8527 6069 8539 6072
rect 8481 6063 8539 6069
rect 8570 6060 8576 6072
rect 8628 6060 8634 6112
rect 8662 6060 8668 6112
rect 8720 6100 8726 6112
rect 9030 6100 9036 6112
rect 8720 6072 8765 6100
rect 8991 6072 9036 6100
rect 8720 6060 8726 6072
rect 9030 6060 9036 6072
rect 9088 6060 9094 6112
rect 9217 6103 9275 6109
rect 9217 6069 9229 6103
rect 9263 6100 9275 6103
rect 10686 6100 10692 6112
rect 9263 6072 10692 6100
rect 9263 6069 9275 6072
rect 9217 6063 9275 6069
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 11698 6100 11704 6112
rect 11659 6072 11704 6100
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 14274 6060 14280 6112
rect 14332 6100 14338 6112
rect 14734 6100 14740 6112
rect 14332 6072 14740 6100
rect 14332 6060 14338 6072
rect 14734 6060 14740 6072
rect 14792 6100 14798 6112
rect 15838 6100 15844 6112
rect 14792 6072 15844 6100
rect 14792 6060 14798 6072
rect 15838 6060 15844 6072
rect 15896 6060 15902 6112
rect 0 6010 18860 6032
rect 0 5958 3110 6010
rect 3162 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 3302 6010
rect 3354 5958 3366 6010
rect 3418 5958 6210 6010
rect 6262 5958 6274 6010
rect 6326 5958 6338 6010
rect 6390 5958 6402 6010
rect 6454 5958 6466 6010
rect 6518 5958 9310 6010
rect 9362 5958 9374 6010
rect 9426 5958 9438 6010
rect 9490 5958 9502 6010
rect 9554 5958 9566 6010
rect 9618 5958 12410 6010
rect 12462 5958 12474 6010
rect 12526 5958 12538 6010
rect 12590 5958 12602 6010
rect 12654 5958 12666 6010
rect 12718 5958 15510 6010
rect 15562 5958 15574 6010
rect 15626 5958 15638 6010
rect 15690 5958 15702 6010
rect 15754 5958 15766 6010
rect 15818 5958 18860 6010
rect 0 5936 18860 5958
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 3099 5899 3157 5905
rect 3099 5896 3111 5899
rect 2924 5868 3111 5896
rect 2924 5856 2930 5868
rect 3099 5865 3111 5868
rect 3145 5865 3157 5899
rect 3099 5859 3157 5865
rect 4430 5856 4436 5908
rect 4488 5896 4494 5908
rect 6546 5896 6552 5908
rect 4488 5868 6224 5896
rect 6507 5868 6552 5896
rect 4488 5856 4494 5868
rect 290 5720 296 5772
rect 348 5760 354 5772
rect 4157 5763 4215 5769
rect 4157 5760 4169 5763
rect 348 5732 4169 5760
rect 348 5720 354 5732
rect 1044 5701 1072 5732
rect 4157 5729 4169 5732
rect 4203 5760 4215 5763
rect 6086 5760 6092 5772
rect 4203 5732 6092 5760
rect 4203 5729 4215 5732
rect 4157 5723 4215 5729
rect 6086 5720 6092 5732
rect 6144 5720 6150 5772
rect 6196 5769 6224 5868
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 8294 5896 8300 5908
rect 8255 5868 8300 5896
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 10597 5899 10655 5905
rect 10597 5865 10609 5899
rect 10643 5896 10655 5899
rect 15378 5896 15384 5908
rect 10643 5868 15384 5896
rect 10643 5865 10655 5868
rect 10597 5859 10655 5865
rect 6270 5788 6276 5840
rect 6328 5828 6334 5840
rect 6328 5800 6960 5828
rect 6328 5788 6334 5800
rect 6932 5769 6960 5800
rect 6181 5763 6239 5769
rect 6181 5729 6193 5763
rect 6227 5760 6239 5763
rect 6917 5763 6975 5769
rect 6227 5732 6408 5760
rect 6227 5729 6239 5732
rect 6181 5723 6239 5729
rect 1029 5695 1087 5701
rect 1029 5661 1041 5695
rect 1075 5661 1087 5695
rect 1029 5655 1087 5661
rect 1121 5695 1179 5701
rect 1121 5661 1133 5695
rect 1167 5692 1179 5695
rect 1305 5695 1363 5701
rect 1305 5692 1317 5695
rect 1167 5664 1317 5692
rect 1167 5661 1179 5664
rect 1121 5655 1179 5661
rect 1305 5661 1317 5664
rect 1351 5661 1363 5695
rect 1673 5695 1731 5701
rect 1673 5692 1685 5695
rect 1305 5655 1363 5661
rect 1412 5664 1685 5692
rect 1210 5584 1216 5636
rect 1268 5624 1274 5636
rect 1412 5624 1440 5664
rect 1673 5661 1685 5664
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 5718 5652 5724 5704
rect 5776 5692 5782 5704
rect 6273 5695 6331 5701
rect 6273 5692 6285 5695
rect 5776 5664 6285 5692
rect 5776 5652 5782 5664
rect 6273 5661 6285 5664
rect 6319 5661 6331 5695
rect 6380 5692 6408 5732
rect 6917 5729 6929 5763
rect 6963 5729 6975 5763
rect 6917 5723 6975 5729
rect 7173 5695 7231 5701
rect 7173 5692 7185 5695
rect 6380 5664 7185 5692
rect 6273 5655 6331 5661
rect 7173 5661 7185 5664
rect 7219 5692 7231 5695
rect 8018 5692 8024 5704
rect 7219 5664 8024 5692
rect 7219 5661 7231 5664
rect 7173 5655 7231 5661
rect 4430 5624 4436 5636
rect 1268 5596 1440 5624
rect 1268 5584 1274 5596
rect 2222 5516 2228 5568
rect 2280 5556 2286 5568
rect 2700 5556 2728 5610
rect 4391 5596 4436 5624
rect 4430 5584 4436 5596
rect 4488 5584 4494 5636
rect 6288 5624 6316 5655
rect 8018 5652 8024 5664
rect 8076 5692 8082 5704
rect 8662 5692 8668 5704
rect 8076 5664 8668 5692
rect 8076 5652 8082 5664
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 10413 5695 10471 5701
rect 10413 5661 10425 5695
rect 10459 5692 10471 5695
rect 10612 5692 10640 5859
rect 15378 5856 15384 5868
rect 15436 5856 15442 5908
rect 16025 5899 16083 5905
rect 16025 5865 16037 5899
rect 16071 5896 16083 5899
rect 16942 5896 16948 5908
rect 16071 5868 16948 5896
rect 16071 5865 16083 5868
rect 16025 5859 16083 5865
rect 16942 5856 16948 5868
rect 17000 5856 17006 5908
rect 14458 5828 14464 5840
rect 13280 5800 14464 5828
rect 11149 5763 11207 5769
rect 11149 5729 11161 5763
rect 11195 5760 11207 5763
rect 11422 5760 11428 5772
rect 11195 5732 11428 5760
rect 11195 5729 11207 5732
rect 11149 5723 11207 5729
rect 11422 5720 11428 5732
rect 11480 5760 11486 5772
rect 13280 5760 13308 5800
rect 14458 5788 14464 5800
rect 14516 5788 14522 5840
rect 16482 5828 16488 5840
rect 15764 5800 16488 5828
rect 11480 5732 13308 5760
rect 13541 5763 13599 5769
rect 11480 5720 11486 5732
rect 13541 5729 13553 5763
rect 13587 5760 13599 5763
rect 13909 5763 13967 5769
rect 13909 5760 13921 5763
rect 13587 5732 13921 5760
rect 13587 5729 13599 5732
rect 13541 5723 13599 5729
rect 13909 5729 13921 5732
rect 13955 5729 13967 5763
rect 14274 5760 14280 5772
rect 14235 5732 14280 5760
rect 13909 5723 13967 5729
rect 14274 5720 14280 5732
rect 14332 5720 14338 5772
rect 15764 5769 15792 5800
rect 16482 5788 16488 5800
rect 16540 5788 16546 5840
rect 15749 5763 15807 5769
rect 15749 5760 15761 5763
rect 14384 5732 15761 5760
rect 10459 5664 10640 5692
rect 13449 5695 13507 5701
rect 10459 5661 10471 5664
rect 10413 5655 10471 5661
rect 13449 5661 13461 5695
rect 13495 5692 13507 5695
rect 14384 5692 14412 5732
rect 15749 5729 15761 5732
rect 15795 5729 15807 5763
rect 15749 5723 15807 5729
rect 15838 5720 15844 5772
rect 15896 5760 15902 5772
rect 15933 5763 15991 5769
rect 15933 5760 15945 5763
rect 15896 5732 15945 5760
rect 15896 5720 15902 5732
rect 15933 5729 15945 5732
rect 15979 5729 15991 5763
rect 15933 5723 15991 5729
rect 16117 5763 16175 5769
rect 16117 5729 16129 5763
rect 16163 5760 16175 5763
rect 17494 5760 17500 5772
rect 16163 5732 17500 5760
rect 16163 5729 16175 5732
rect 16117 5723 16175 5729
rect 17494 5720 17500 5732
rect 17552 5720 17558 5772
rect 17589 5763 17647 5769
rect 17589 5729 17601 5763
rect 17635 5760 17647 5763
rect 18322 5760 18328 5772
rect 17635 5732 18328 5760
rect 17635 5729 17647 5732
rect 17589 5723 17647 5729
rect 18322 5720 18328 5732
rect 18380 5720 18386 5772
rect 14550 5692 14556 5704
rect 13495 5664 14412 5692
rect 14511 5664 14556 5692
rect 13495 5661 13507 5664
rect 13449 5655 13507 5661
rect 8202 5624 8208 5636
rect 3329 5559 3387 5565
rect 3329 5556 3341 5559
rect 2280 5528 3341 5556
rect 2280 5516 2286 5528
rect 3329 5525 3341 5528
rect 3375 5556 3387 5559
rect 3510 5556 3516 5568
rect 3375 5528 3516 5556
rect 3375 5525 3387 5528
rect 3329 5519 3387 5525
rect 3510 5516 3516 5528
rect 3568 5556 3574 5568
rect 3973 5559 4031 5565
rect 3973 5556 3985 5559
rect 3568 5528 3985 5556
rect 3568 5516 3574 5528
rect 3973 5525 3985 5528
rect 4019 5556 4031 5559
rect 4908 5556 4936 5610
rect 6288 5596 8208 5624
rect 8202 5584 8208 5596
rect 8260 5584 8266 5636
rect 11425 5627 11483 5633
rect 11425 5593 11437 5627
rect 11471 5624 11483 5627
rect 11698 5624 11704 5636
rect 11471 5596 11704 5624
rect 11471 5593 11483 5596
rect 11425 5587 11483 5593
rect 11698 5584 11704 5596
rect 11756 5584 11762 5636
rect 12360 5568 12388 5610
rect 5902 5556 5908 5568
rect 4019 5528 4936 5556
rect 5863 5528 5908 5556
rect 4019 5525 4031 5528
rect 3973 5519 4031 5525
rect 5902 5516 5908 5528
rect 5960 5516 5966 5568
rect 9125 5559 9183 5565
rect 9125 5525 9137 5559
rect 9171 5556 9183 5559
rect 9306 5556 9312 5568
rect 9171 5528 9312 5556
rect 9171 5525 9183 5528
rect 9125 5519 9183 5525
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 10686 5516 10692 5568
rect 10744 5556 10750 5568
rect 11057 5559 11115 5565
rect 11057 5556 11069 5559
rect 10744 5528 11069 5556
rect 10744 5516 10750 5528
rect 11057 5525 11069 5528
rect 11103 5556 11115 5559
rect 12342 5556 12348 5568
rect 11103 5528 12348 5556
rect 11103 5525 11115 5528
rect 11057 5519 11115 5525
rect 12342 5516 12348 5528
rect 12400 5516 12406 5568
rect 12802 5516 12808 5568
rect 12860 5556 12866 5568
rect 12897 5559 12955 5565
rect 12897 5556 12909 5559
rect 12860 5528 12909 5556
rect 12860 5516 12866 5528
rect 12897 5525 12909 5528
rect 12943 5556 12955 5559
rect 13464 5556 13492 5655
rect 14550 5652 14556 5664
rect 14608 5652 14614 5704
rect 15197 5695 15255 5701
rect 15197 5692 15209 5695
rect 14844 5664 15209 5692
rect 13909 5627 13967 5633
rect 13909 5593 13921 5627
rect 13955 5624 13967 5627
rect 14461 5627 14519 5633
rect 14461 5624 14473 5627
rect 13955 5596 14473 5624
rect 13955 5593 13967 5596
rect 13909 5587 13967 5593
rect 14461 5593 14473 5596
rect 14507 5624 14519 5627
rect 14642 5624 14648 5636
rect 14507 5596 14648 5624
rect 14507 5593 14519 5596
rect 14461 5587 14519 5593
rect 14642 5584 14648 5596
rect 14700 5584 14706 5636
rect 13814 5556 13820 5568
rect 12943 5528 13492 5556
rect 13775 5528 13820 5556
rect 12943 5525 12955 5528
rect 12897 5519 12955 5525
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 14093 5559 14151 5565
rect 14093 5525 14105 5559
rect 14139 5556 14151 5559
rect 14366 5556 14372 5568
rect 14139 5528 14372 5556
rect 14139 5525 14151 5528
rect 14093 5519 14151 5525
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 14844 5556 14872 5664
rect 15197 5661 15209 5664
rect 15243 5661 15255 5695
rect 15197 5655 15255 5661
rect 16025 5695 16083 5701
rect 16025 5661 16037 5695
rect 16071 5692 16083 5695
rect 16206 5692 16212 5704
rect 16071 5664 16212 5692
rect 16071 5661 16083 5664
rect 16025 5655 16083 5661
rect 16206 5652 16212 5664
rect 16264 5652 16270 5704
rect 17862 5652 17868 5704
rect 17920 5692 17926 5704
rect 18233 5695 18291 5701
rect 17920 5664 17965 5692
rect 17920 5652 17926 5664
rect 18233 5661 18245 5695
rect 18279 5692 18291 5695
rect 18506 5692 18512 5704
rect 18279 5664 18512 5692
rect 18279 5661 18291 5664
rect 18233 5655 18291 5661
rect 18506 5652 18512 5664
rect 18564 5652 18570 5704
rect 16114 5584 16120 5636
rect 16172 5624 16178 5636
rect 16172 5596 16422 5624
rect 16172 5584 16178 5596
rect 14921 5559 14979 5565
rect 14921 5556 14933 5559
rect 14844 5528 14933 5556
rect 14921 5525 14933 5528
rect 14967 5525 14979 5559
rect 14921 5519 14979 5525
rect 15010 5516 15016 5568
rect 15068 5556 15074 5568
rect 15473 5559 15531 5565
rect 15068 5528 15113 5556
rect 15068 5516 15074 5528
rect 15473 5525 15485 5559
rect 15519 5556 15531 5559
rect 16132 5556 16160 5584
rect 15519 5528 16160 5556
rect 15519 5525 15531 5528
rect 15473 5519 15531 5525
rect 18046 5516 18052 5568
rect 18104 5556 18110 5568
rect 18325 5559 18383 5565
rect 18325 5556 18337 5559
rect 18104 5528 18337 5556
rect 18104 5516 18110 5528
rect 18325 5525 18337 5528
rect 18371 5525 18383 5559
rect 18325 5519 18383 5525
rect 0 5466 18860 5488
rect 0 5414 4660 5466
rect 4712 5414 4724 5466
rect 4776 5414 4788 5466
rect 4840 5414 4852 5466
rect 4904 5414 4916 5466
rect 4968 5414 7760 5466
rect 7812 5414 7824 5466
rect 7876 5414 7888 5466
rect 7940 5414 7952 5466
rect 8004 5414 8016 5466
rect 8068 5414 10860 5466
rect 10912 5414 10924 5466
rect 10976 5414 10988 5466
rect 11040 5414 11052 5466
rect 11104 5414 11116 5466
rect 11168 5414 13960 5466
rect 14012 5414 14024 5466
rect 14076 5414 14088 5466
rect 14140 5414 14152 5466
rect 14204 5414 14216 5466
rect 14268 5414 17060 5466
rect 17112 5414 17124 5466
rect 17176 5414 17188 5466
rect 17240 5414 17252 5466
rect 17304 5414 17316 5466
rect 17368 5414 18860 5466
rect 0 5392 18860 5414
rect 1210 5352 1216 5364
rect 1171 5324 1216 5352
rect 1210 5312 1216 5324
rect 1268 5312 1274 5364
rect 2317 5355 2375 5361
rect 2317 5321 2329 5355
rect 2363 5352 2375 5355
rect 2774 5352 2780 5364
rect 2363 5324 2780 5352
rect 2363 5321 2375 5324
rect 2317 5315 2375 5321
rect 2774 5312 2780 5324
rect 2832 5312 2838 5364
rect 2958 5352 2964 5364
rect 2919 5324 2964 5352
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 4430 5312 4436 5364
rect 4488 5352 4494 5364
rect 4525 5355 4583 5361
rect 4525 5352 4537 5355
rect 4488 5324 4537 5352
rect 4488 5312 4494 5324
rect 4525 5321 4537 5324
rect 4571 5321 4583 5355
rect 4525 5315 4583 5321
rect 4893 5355 4951 5361
rect 4893 5321 4905 5355
rect 4939 5321 4951 5355
rect 4893 5315 4951 5321
rect 5353 5355 5411 5361
rect 5353 5321 5365 5355
rect 5399 5352 5411 5355
rect 5534 5352 5540 5364
rect 5399 5324 5540 5352
rect 5399 5321 5411 5324
rect 5353 5315 5411 5321
rect 2498 5244 2504 5296
rect 2556 5284 2562 5296
rect 2556 5256 3096 5284
rect 2556 5244 2562 5256
rect 1029 5219 1087 5225
rect 1029 5185 1041 5219
rect 1075 5185 1087 5219
rect 1029 5179 1087 5185
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5216 2007 5219
rect 2866 5216 2872 5228
rect 1995 5188 2872 5216
rect 1995 5185 2007 5188
rect 1949 5179 2007 5185
rect 1044 5080 1072 5179
rect 2866 5176 2872 5188
rect 2924 5176 2930 5228
rect 2041 5151 2099 5157
rect 2041 5117 2053 5151
rect 2087 5148 2099 5151
rect 2682 5148 2688 5160
rect 2087 5120 2688 5148
rect 2087 5117 2099 5120
rect 2041 5111 2099 5117
rect 2682 5108 2688 5120
rect 2740 5108 2746 5160
rect 3068 5157 3096 5256
rect 3513 5219 3571 5225
rect 3513 5185 3525 5219
rect 3559 5216 3571 5219
rect 3602 5216 3608 5228
rect 3559 5188 3608 5216
rect 3559 5185 3571 5188
rect 3513 5179 3571 5185
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4709 5219 4767 5225
rect 4709 5185 4721 5219
rect 4755 5216 4767 5219
rect 4908 5216 4936 5315
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 6086 5312 6092 5364
rect 6144 5352 6150 5364
rect 6825 5355 6883 5361
rect 6825 5352 6837 5355
rect 6144 5324 6837 5352
rect 6144 5312 6150 5324
rect 6825 5321 6837 5324
rect 6871 5352 6883 5355
rect 7466 5352 7472 5364
rect 6871 5324 7472 5352
rect 6871 5321 6883 5324
rect 6825 5315 6883 5321
rect 7466 5312 7472 5324
rect 7524 5352 7530 5364
rect 8478 5352 8484 5364
rect 7524 5324 8484 5352
rect 7524 5312 7530 5324
rect 8478 5312 8484 5324
rect 8536 5312 8542 5364
rect 9214 5312 9220 5364
rect 9272 5352 9278 5364
rect 11330 5352 11336 5364
rect 9272 5324 11336 5352
rect 9272 5312 9278 5324
rect 11330 5312 11336 5324
rect 11388 5312 11394 5364
rect 11514 5312 11520 5364
rect 11572 5352 11578 5364
rect 12069 5355 12127 5361
rect 12069 5352 12081 5355
rect 11572 5324 12081 5352
rect 11572 5312 11578 5324
rect 12069 5321 12081 5324
rect 12115 5321 12127 5355
rect 12069 5315 12127 5321
rect 12526 5312 12532 5364
rect 12584 5352 12590 5364
rect 13446 5352 13452 5364
rect 12584 5324 13452 5352
rect 12584 5312 12590 5324
rect 5994 5244 6000 5296
rect 6052 5284 6058 5296
rect 6181 5287 6239 5293
rect 6181 5284 6193 5287
rect 6052 5256 6193 5284
rect 6052 5244 6058 5256
rect 6181 5253 6193 5256
rect 6227 5253 6239 5287
rect 6181 5247 6239 5253
rect 6917 5287 6975 5293
rect 6917 5253 6929 5287
rect 6963 5284 6975 5287
rect 9306 5284 9312 5296
rect 6963 5256 9312 5284
rect 6963 5253 6975 5256
rect 6917 5247 6975 5253
rect 9306 5244 9312 5256
rect 9364 5284 9370 5296
rect 11241 5287 11299 5293
rect 11241 5284 11253 5287
rect 9364 5256 11253 5284
rect 9364 5244 9370 5256
rect 11241 5253 11253 5256
rect 11287 5253 11299 5287
rect 13096 5270 13124 5324
rect 13446 5312 13452 5324
rect 13504 5312 13510 5364
rect 17954 5352 17960 5364
rect 14568 5324 17960 5352
rect 11241 5247 11299 5253
rect 13262 5244 13268 5296
rect 13320 5284 13326 5296
rect 13320 5256 13860 5284
rect 13320 5244 13326 5256
rect 4755 5188 4936 5216
rect 5261 5219 5319 5225
rect 4755 5185 4767 5188
rect 4709 5179 4767 5185
rect 5261 5185 5273 5219
rect 5307 5216 5319 5219
rect 5902 5216 5908 5228
rect 5307 5188 5908 5216
rect 5307 5185 5319 5188
rect 5261 5179 5319 5185
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5117 3111 5151
rect 3053 5111 3111 5117
rect 3421 5151 3479 5157
rect 3421 5117 3433 5151
rect 3467 5148 3479 5151
rect 3878 5148 3884 5160
rect 3467 5120 3884 5148
rect 3467 5117 3479 5120
rect 3421 5111 3479 5117
rect 3878 5108 3884 5120
rect 3936 5108 3942 5160
rect 2501 5083 2559 5089
rect 2501 5080 2513 5083
rect 1044 5052 2513 5080
rect 2501 5049 2513 5052
rect 2547 5049 2559 5083
rect 2700 5080 2728 5108
rect 5276 5080 5304 5179
rect 5902 5176 5908 5188
rect 5960 5176 5966 5228
rect 8481 5219 8539 5225
rect 8481 5185 8493 5219
rect 8527 5216 8539 5219
rect 8846 5216 8852 5228
rect 8527 5188 8852 5216
rect 8527 5185 8539 5188
rect 8481 5179 8539 5185
rect 8846 5176 8852 5188
rect 8904 5176 8910 5228
rect 9030 5176 9036 5228
rect 9088 5216 9094 5228
rect 9125 5219 9183 5225
rect 9125 5216 9137 5219
rect 9088 5188 9137 5216
rect 9088 5176 9094 5188
rect 9125 5185 9137 5188
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 9217 5219 9275 5225
rect 9217 5185 9229 5219
rect 9263 5185 9275 5219
rect 9217 5179 9275 5185
rect 9401 5219 9459 5225
rect 9401 5185 9413 5219
rect 9447 5216 9459 5219
rect 9447 5188 9720 5216
rect 9447 5185 9459 5188
rect 9401 5179 9459 5185
rect 5442 5148 5448 5160
rect 5403 5120 5448 5148
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 8202 5108 8208 5160
rect 8260 5148 8266 5160
rect 8389 5151 8447 5157
rect 8389 5148 8401 5151
rect 8260 5120 8401 5148
rect 8260 5108 8266 5120
rect 8389 5117 8401 5120
rect 8435 5117 8447 5151
rect 8389 5111 8447 5117
rect 8570 5108 8576 5160
rect 8628 5148 8634 5160
rect 9232 5148 9260 5179
rect 8628 5120 9260 5148
rect 8628 5108 8634 5120
rect 2700 5052 5304 5080
rect 8849 5083 8907 5089
rect 2501 5043 2559 5049
rect 8849 5049 8861 5083
rect 8895 5080 8907 5083
rect 9214 5080 9220 5092
rect 8895 5052 9220 5080
rect 8895 5049 8907 5052
rect 8849 5043 8907 5049
rect 9214 5040 9220 5052
rect 9272 5040 9278 5092
rect 9692 5089 9720 5188
rect 10778 5176 10784 5228
rect 10836 5225 10842 5228
rect 10836 5216 10848 5225
rect 11057 5219 11115 5225
rect 10836 5188 10881 5216
rect 10836 5179 10848 5188
rect 11057 5185 11069 5219
rect 11103 5216 11115 5219
rect 11422 5216 11428 5228
rect 11103 5188 11428 5216
rect 11103 5185 11115 5188
rect 11057 5179 11115 5185
rect 10836 5176 10842 5179
rect 11422 5176 11428 5188
rect 11480 5176 11486 5228
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5185 11575 5219
rect 11698 5216 11704 5228
rect 11659 5188 11704 5216
rect 11517 5179 11575 5185
rect 11532 5148 11560 5179
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 13832 5225 13860 5256
rect 13817 5219 13875 5225
rect 13817 5185 13829 5219
rect 13863 5185 13875 5219
rect 14458 5216 14464 5228
rect 14419 5188 14464 5216
rect 13817 5179 13875 5185
rect 14458 5176 14464 5188
rect 14516 5176 14522 5228
rect 13541 5151 13599 5157
rect 11532 5120 11836 5148
rect 9677 5083 9735 5089
rect 9677 5049 9689 5083
rect 9723 5049 9735 5083
rect 9677 5043 9735 5049
rect 11808 5024 11836 5120
rect 13541 5117 13553 5151
rect 13587 5148 13599 5151
rect 14568 5148 14596 5324
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 16114 5284 16120 5296
rect 15870 5256 16120 5284
rect 16114 5244 16120 5256
rect 16172 5244 16178 5296
rect 16206 5244 16212 5296
rect 16264 5293 16270 5296
rect 16264 5287 16313 5293
rect 16264 5253 16267 5287
rect 16301 5253 16313 5287
rect 16264 5247 16313 5253
rect 16264 5244 16270 5247
rect 16577 5219 16635 5225
rect 16577 5185 16589 5219
rect 16623 5185 16635 5219
rect 16577 5179 16635 5185
rect 17221 5219 17279 5225
rect 17221 5185 17233 5219
rect 17267 5216 17279 5219
rect 17402 5216 17408 5228
rect 17267 5188 17408 5216
rect 17267 5185 17279 5188
rect 17221 5179 17279 5185
rect 13587 5120 14596 5148
rect 14829 5151 14887 5157
rect 13587 5117 13599 5120
rect 13541 5111 13599 5117
rect 14829 5117 14841 5151
rect 14875 5148 14887 5151
rect 15010 5148 15016 5160
rect 14875 5120 15016 5148
rect 14875 5117 14887 5120
rect 14829 5111 14887 5117
rect 15010 5108 15016 5120
rect 15068 5108 15074 5160
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 16592 5148 16620 5179
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 15436 5120 16620 5148
rect 15436 5108 15442 5120
rect 16942 5108 16948 5160
rect 17000 5148 17006 5160
rect 17129 5151 17187 5157
rect 17129 5148 17141 5151
rect 17000 5120 17141 5148
rect 17000 5108 17006 5120
rect 17129 5117 17141 5120
rect 17175 5117 17187 5151
rect 17129 5111 17187 5117
rect 16393 5083 16451 5089
rect 16393 5080 16405 5083
rect 15580 5052 16405 5080
rect 3789 5015 3847 5021
rect 3789 4981 3801 5015
rect 3835 5012 3847 5015
rect 4062 5012 4068 5024
rect 3835 4984 4068 5012
rect 3835 4981 3847 4984
rect 3789 4975 3847 4981
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 8386 4972 8392 5024
rect 8444 5012 8450 5024
rect 9125 5015 9183 5021
rect 9125 5012 9137 5015
rect 8444 4984 9137 5012
rect 8444 4972 8450 4984
rect 9125 4981 9137 4984
rect 9171 4981 9183 5015
rect 11514 5012 11520 5024
rect 11475 4984 11520 5012
rect 9125 4975 9183 4981
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 11790 5012 11796 5024
rect 11751 4984 11796 5012
rect 11790 4972 11796 4984
rect 11848 4972 11854 5024
rect 14277 5015 14335 5021
rect 14277 4981 14289 5015
rect 14323 5012 14335 5015
rect 14366 5012 14372 5024
rect 14323 4984 14372 5012
rect 14323 4981 14335 4984
rect 14277 4975 14335 4981
rect 14366 4972 14372 4984
rect 14424 5012 14430 5024
rect 15194 5012 15200 5024
rect 14424 4984 15200 5012
rect 14424 4972 14430 4984
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 15286 4972 15292 5024
rect 15344 5012 15350 5024
rect 15580 5012 15608 5052
rect 16393 5049 16405 5052
rect 16439 5049 16451 5083
rect 16393 5043 16451 5049
rect 16574 5040 16580 5092
rect 16632 5080 16638 5092
rect 16853 5083 16911 5089
rect 16853 5080 16865 5083
rect 16632 5052 16865 5080
rect 16632 5040 16638 5052
rect 16853 5049 16865 5052
rect 16899 5049 16911 5083
rect 16853 5043 16911 5049
rect 15344 4984 15608 5012
rect 15344 4972 15350 4984
rect 0 4922 18860 4944
rect 0 4870 3110 4922
rect 3162 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 3302 4922
rect 3354 4870 3366 4922
rect 3418 4870 6210 4922
rect 6262 4870 6274 4922
rect 6326 4870 6338 4922
rect 6390 4870 6402 4922
rect 6454 4870 6466 4922
rect 6518 4870 9310 4922
rect 9362 4870 9374 4922
rect 9426 4870 9438 4922
rect 9490 4870 9502 4922
rect 9554 4870 9566 4922
rect 9618 4870 12410 4922
rect 12462 4870 12474 4922
rect 12526 4870 12538 4922
rect 12590 4870 12602 4922
rect 12654 4870 12666 4922
rect 12718 4870 15510 4922
rect 15562 4870 15574 4922
rect 15626 4870 15638 4922
rect 15690 4870 15702 4922
rect 15754 4870 15766 4922
rect 15818 4870 18860 4922
rect 0 4848 18860 4870
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 8202 4808 8208 4820
rect 5592 4780 7972 4808
rect 8163 4780 8208 4808
rect 5592 4768 5598 4780
rect 5810 4740 5816 4752
rect 4632 4712 5816 4740
rect 3970 4632 3976 4684
rect 4028 4672 4034 4684
rect 4341 4675 4399 4681
rect 4341 4672 4353 4675
rect 4028 4644 4353 4672
rect 4028 4632 4034 4644
rect 4341 4641 4353 4644
rect 4387 4672 4399 4675
rect 4525 4675 4583 4681
rect 4525 4672 4537 4675
rect 4387 4644 4537 4672
rect 4387 4641 4399 4644
rect 4341 4635 4399 4641
rect 4525 4641 4537 4644
rect 4571 4641 4583 4675
rect 4525 4635 4583 4641
rect 845 4607 903 4613
rect 845 4573 857 4607
rect 891 4604 903 4607
rect 1118 4604 1124 4616
rect 891 4576 1124 4604
rect 891 4573 903 4576
rect 845 4567 903 4573
rect 1118 4564 1124 4576
rect 1176 4564 1182 4616
rect 1302 4604 1308 4616
rect 1263 4576 1308 4604
rect 1302 4564 1308 4576
rect 1360 4564 1366 4616
rect 4062 4604 4068 4616
rect 4023 4576 4068 4604
rect 4062 4564 4068 4576
rect 4120 4564 4126 4616
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4604 4215 4607
rect 4632 4604 4660 4712
rect 5810 4700 5816 4712
rect 5868 4700 5874 4752
rect 5905 4743 5963 4749
rect 5905 4709 5917 4743
rect 5951 4740 5963 4743
rect 5951 4712 6224 4740
rect 5951 4709 5963 4712
rect 5905 4703 5963 4709
rect 4801 4675 4859 4681
rect 4801 4641 4813 4675
rect 4847 4672 4859 4675
rect 5626 4672 5632 4684
rect 4847 4644 5488 4672
rect 5587 4644 5632 4672
rect 4847 4641 4859 4644
rect 4801 4635 4859 4641
rect 4203 4576 4660 4604
rect 4709 4607 4767 4613
rect 4203 4573 4215 4576
rect 4157 4567 4215 4573
rect 4709 4573 4721 4607
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4604 4951 4607
rect 5460 4604 5488 4644
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 6086 4672 6092 4684
rect 6047 4644 6092 4672
rect 6086 4632 6092 4644
rect 6144 4632 6150 4684
rect 6196 4672 6224 4712
rect 6365 4675 6423 4681
rect 6365 4672 6377 4675
rect 6196 4644 6377 4672
rect 6365 4641 6377 4644
rect 6411 4641 6423 4675
rect 6365 4635 6423 4641
rect 7944 4613 7972 4780
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 8846 4768 8852 4820
rect 8904 4808 8910 4820
rect 10643 4811 10701 4817
rect 10643 4808 10655 4811
rect 8904 4780 10655 4808
rect 8904 4768 8910 4780
rect 10643 4777 10655 4780
rect 10689 4808 10701 4811
rect 10689 4780 10824 4808
rect 10689 4777 10701 4780
rect 10643 4771 10701 4777
rect 8849 4675 8907 4681
rect 8849 4641 8861 4675
rect 8895 4672 8907 4675
rect 9122 4672 9128 4684
rect 8895 4644 9128 4672
rect 8895 4641 8907 4644
rect 8849 4635 8907 4641
rect 9122 4632 9128 4644
rect 9180 4632 9186 4684
rect 9214 4632 9220 4684
rect 9272 4672 9278 4684
rect 9272 4644 9317 4672
rect 9272 4632 9278 4644
rect 5537 4607 5595 4613
rect 5537 4604 5549 4607
rect 4939 4576 5120 4604
rect 5460 4576 5549 4604
rect 4939 4573 4951 4576
rect 4893 4567 4951 4573
rect 1581 4539 1639 4545
rect 1581 4536 1593 4539
rect 1044 4508 1593 4536
rect 1044 4477 1072 4508
rect 1581 4505 1593 4508
rect 1627 4505 1639 4539
rect 1581 4499 1639 4505
rect 1854 4496 1860 4548
rect 1912 4536 1918 4548
rect 3237 4539 3295 4545
rect 3237 4536 3249 4539
rect 1912 4522 2070 4536
rect 1912 4508 2084 4522
rect 1912 4496 1918 4508
rect 1029 4471 1087 4477
rect 1029 4437 1041 4471
rect 1075 4437 1087 4471
rect 2056 4468 2084 4508
rect 2884 4508 3249 4536
rect 2884 4468 2912 4508
rect 3237 4505 3249 4508
rect 3283 4536 3295 4539
rect 3510 4536 3516 4548
rect 3283 4508 3516 4536
rect 3283 4505 3295 4508
rect 3237 4499 3295 4505
rect 3510 4496 3516 4508
rect 3568 4496 3574 4548
rect 4724 4536 4752 4567
rect 4982 4536 4988 4548
rect 4724 4508 4988 4536
rect 4982 4496 4988 4508
rect 5040 4496 5046 4548
rect 5092 4536 5120 4576
rect 5537 4573 5549 4576
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4573 7987 4607
rect 8202 4604 8208 4616
rect 8163 4576 8208 4604
rect 7929 4567 7987 4573
rect 5442 4536 5448 4548
rect 5092 4508 5448 4536
rect 5442 4496 5448 4508
rect 5500 4496 5506 4548
rect 3050 4468 3056 4480
rect 2056 4440 2912 4468
rect 3011 4440 3056 4468
rect 1029 4431 1087 4437
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 3694 4468 3700 4480
rect 3655 4440 3700 4468
rect 3694 4428 3700 4440
rect 3752 4428 3758 4480
rect 5552 4468 5580 4567
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 10796 4604 10824 4780
rect 11330 4672 11336 4684
rect 11291 4644 11336 4672
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 11514 4672 11520 4684
rect 11475 4644 11520 4672
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 13078 4632 13084 4684
rect 13136 4672 13142 4684
rect 13449 4675 13507 4681
rect 13449 4672 13461 4675
rect 13136 4644 13461 4672
rect 13136 4632 13142 4644
rect 13449 4641 13461 4644
rect 13495 4641 13507 4675
rect 13449 4635 13507 4641
rect 16117 4675 16175 4681
rect 16117 4641 16129 4675
rect 16163 4672 16175 4675
rect 16574 4672 16580 4684
rect 16163 4644 16580 4672
rect 16163 4641 16175 4644
rect 16117 4635 16175 4641
rect 16574 4632 16580 4644
rect 16632 4632 16638 4684
rect 17494 4672 17500 4684
rect 17455 4644 17500 4672
rect 17494 4632 17500 4644
rect 17552 4632 17558 4684
rect 11241 4607 11299 4613
rect 11241 4604 11253 4607
rect 10796 4576 11253 4604
rect 11241 4573 11253 4576
rect 11287 4573 11299 4607
rect 11348 4604 11376 4632
rect 13262 4604 13268 4616
rect 11348 4576 13268 4604
rect 11241 4567 11299 4573
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 15010 4564 15016 4616
rect 15068 4604 15074 4616
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 15068 4576 15761 4604
rect 15068 4564 15074 4576
rect 15749 4573 15761 4576
rect 15795 4604 15807 4607
rect 15838 4604 15844 4616
rect 15795 4576 15844 4604
rect 15795 4573 15807 4576
rect 15749 4567 15807 4573
rect 15838 4564 15844 4576
rect 15896 4564 15902 4616
rect 17512 4604 17540 4632
rect 18141 4607 18199 4613
rect 18141 4604 18153 4607
rect 17512 4576 18153 4604
rect 18141 4573 18153 4576
rect 18187 4573 18199 4607
rect 18141 4567 18199 4573
rect 7006 4496 7012 4548
rect 7064 4496 7070 4548
rect 8113 4539 8171 4545
rect 8113 4505 8125 4539
rect 8159 4536 8171 4539
rect 8938 4536 8944 4548
rect 8159 4508 8944 4536
rect 8159 4505 8171 4508
rect 8113 4499 8171 4505
rect 8938 4496 8944 4508
rect 8996 4496 9002 4548
rect 11885 4539 11943 4545
rect 11885 4536 11897 4539
rect 10258 4522 11897 4536
rect 10244 4508 11897 4522
rect 7374 4468 7380 4480
rect 5552 4440 7380 4468
rect 7374 4428 7380 4440
rect 7432 4468 7438 4480
rect 7837 4471 7895 4477
rect 7837 4468 7849 4471
rect 7432 4440 7849 4468
rect 7432 4428 7438 4440
rect 7837 4437 7849 4440
rect 7883 4437 7895 4471
rect 7837 4431 7895 4437
rect 8757 4471 8815 4477
rect 8757 4437 8769 4471
rect 8803 4468 8815 4471
rect 9122 4468 9128 4480
rect 8803 4440 9128 4468
rect 8803 4437 8815 4440
rect 8757 4431 8815 4437
rect 9122 4428 9128 4440
rect 9180 4468 9186 4480
rect 10244 4468 10272 4508
rect 11885 4505 11897 4508
rect 11931 4505 11943 4539
rect 13722 4536 13728 4548
rect 13683 4508 13728 4536
rect 11885 4499 11943 4505
rect 9180 4440 10272 4468
rect 9180 4428 9186 4440
rect 10778 4428 10784 4480
rect 10836 4468 10842 4480
rect 10873 4471 10931 4477
rect 10873 4468 10885 4471
rect 10836 4440 10885 4468
rect 10836 4428 10842 4440
rect 10873 4437 10885 4440
rect 10919 4437 10931 4471
rect 11900 4468 11928 4499
rect 13722 4496 13728 4508
rect 13780 4496 13786 4548
rect 12434 4468 12440 4480
rect 11900 4440 12440 4468
rect 10873 4431 10931 4437
rect 12434 4428 12440 4440
rect 12492 4468 12498 4480
rect 13357 4471 13415 4477
rect 13357 4468 13369 4471
rect 12492 4440 13369 4468
rect 12492 4428 12498 4440
rect 13357 4437 13369 4440
rect 13403 4468 13415 4471
rect 13446 4468 13452 4480
rect 13403 4440 13452 4468
rect 13403 4437 13415 4440
rect 13357 4431 13415 4437
rect 13446 4428 13452 4440
rect 13504 4468 13510 4480
rect 14936 4468 14964 4522
rect 15378 4496 15384 4548
rect 15436 4536 15442 4548
rect 15473 4539 15531 4545
rect 15473 4536 15485 4539
rect 15436 4508 15485 4536
rect 15436 4496 15442 4508
rect 15473 4505 15485 4508
rect 15519 4505 15531 4539
rect 15473 4499 15531 4505
rect 15194 4468 15200 4480
rect 13504 4440 15200 4468
rect 13504 4428 13510 4440
rect 15194 4428 15200 4440
rect 15252 4468 15258 4480
rect 16114 4468 16120 4480
rect 15252 4440 16120 4468
rect 15252 4428 15258 4440
rect 16114 4428 16120 4440
rect 16172 4468 16178 4480
rect 16500 4468 16528 4522
rect 16172 4440 16528 4468
rect 16172 4428 16178 4440
rect 17770 4428 17776 4480
rect 17828 4468 17834 4480
rect 18233 4471 18291 4477
rect 18233 4468 18245 4471
rect 17828 4440 18245 4468
rect 17828 4428 17834 4440
rect 18233 4437 18245 4440
rect 18279 4437 18291 4471
rect 18233 4431 18291 4437
rect 0 4378 18860 4400
rect 0 4326 4660 4378
rect 4712 4326 4724 4378
rect 4776 4326 4788 4378
rect 4840 4326 4852 4378
rect 4904 4326 4916 4378
rect 4968 4326 7760 4378
rect 7812 4326 7824 4378
rect 7876 4326 7888 4378
rect 7940 4326 7952 4378
rect 8004 4326 8016 4378
rect 8068 4326 10860 4378
rect 10912 4326 10924 4378
rect 10976 4326 10988 4378
rect 11040 4326 11052 4378
rect 11104 4326 11116 4378
rect 11168 4326 13960 4378
rect 14012 4326 14024 4378
rect 14076 4326 14088 4378
rect 14140 4326 14152 4378
rect 14204 4326 14216 4378
rect 14268 4326 17060 4378
rect 17112 4326 17124 4378
rect 17176 4326 17188 4378
rect 17240 4326 17252 4378
rect 17304 4326 17316 4378
rect 17368 4326 18860 4378
rect 0 4304 18860 4326
rect 2961 4267 3019 4273
rect 2961 4233 2973 4267
rect 3007 4264 3019 4267
rect 3694 4264 3700 4276
rect 3007 4236 3700 4264
rect 3007 4233 3019 4236
rect 2961 4227 3019 4233
rect 3694 4224 3700 4236
rect 3752 4224 3758 4276
rect 5626 4264 5632 4276
rect 5587 4236 5632 4264
rect 5626 4224 5632 4236
rect 5684 4224 5690 4276
rect 6089 4267 6147 4273
rect 6089 4233 6101 4267
rect 6135 4264 6147 4267
rect 7006 4264 7012 4276
rect 6135 4236 7012 4264
rect 6135 4233 6147 4236
rect 6089 4227 6147 4233
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 7377 4267 7435 4273
rect 7377 4233 7389 4267
rect 7423 4264 7435 4267
rect 8202 4264 8208 4276
rect 7423 4236 8208 4264
rect 7423 4233 7435 4236
rect 7377 4227 7435 4233
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 12437 4267 12495 4273
rect 12437 4233 12449 4267
rect 12483 4264 12495 4267
rect 13722 4264 13728 4276
rect 12483 4236 13728 4264
rect 12483 4233 12495 4236
rect 12437 4227 12495 4233
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 17954 4264 17960 4276
rect 17915 4236 17960 4264
rect 17954 4224 17960 4236
rect 18012 4224 18018 4276
rect 1860 4208 1912 4214
rect 3050 4196 3056 4208
rect 2963 4168 3056 4196
rect 3050 4156 3056 4168
rect 3108 4196 3114 4208
rect 3602 4196 3608 4208
rect 3108 4168 3608 4196
rect 3108 4156 3114 4168
rect 3602 4156 3608 4168
rect 3660 4196 3666 4208
rect 4982 4196 4988 4208
rect 3660 4168 4988 4196
rect 3660 4156 3666 4168
rect 4982 4156 4988 4168
rect 5040 4196 5046 4208
rect 11790 4196 11796 4208
rect 5040 4168 5764 4196
rect 5040 4156 5046 4168
rect 1860 4150 1912 4156
rect 477 4131 535 4137
rect 477 4097 489 4131
rect 523 4128 535 4131
rect 2317 4131 2375 4137
rect 523 4100 980 4128
rect 523 4097 535 4100
rect 477 4091 535 4097
rect 842 4060 848 4072
rect 803 4032 848 4060
rect 842 4020 848 4032
rect 900 4020 906 4072
rect 952 4060 980 4100
rect 2317 4097 2329 4131
rect 2363 4128 2375 4131
rect 3786 4128 3792 4140
rect 2363 4100 3648 4128
rect 3747 4100 3792 4128
rect 2363 4097 2375 4100
rect 2317 4091 2375 4097
rect 1302 4060 1308 4072
rect 952 4032 1308 4060
rect 1302 4020 1308 4032
rect 1360 4020 1366 4072
rect 3237 4063 3295 4069
rect 3237 4029 3249 4063
rect 3283 4029 3295 4063
rect 3620 4060 3648 4100
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 3878 4088 3884 4140
rect 3936 4128 3942 4140
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 3936 4100 4537 4128
rect 3936 4088 3942 4100
rect 4525 4097 4537 4100
rect 4571 4128 4583 4131
rect 5534 4128 5540 4140
rect 4571 4100 5540 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 5534 4088 5540 4100
rect 5592 4128 5598 4140
rect 5736 4137 5764 4168
rect 8680 4168 11796 4196
rect 5629 4131 5687 4137
rect 5629 4128 5641 4131
rect 5592 4100 5641 4128
rect 5592 4088 5598 4100
rect 5629 4097 5641 4100
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4128 5779 4131
rect 7285 4131 7343 4137
rect 7285 4128 7297 4131
rect 5767 4100 7297 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 7285 4097 7297 4100
rect 7331 4097 7343 4131
rect 7285 4091 7343 4097
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 7469 4131 7527 4137
rect 7469 4128 7481 4131
rect 7432 4100 7481 4128
rect 7432 4088 7438 4100
rect 7469 4097 7481 4100
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 8202 4088 8208 4140
rect 8260 4128 8266 4140
rect 8680 4128 8708 4168
rect 11790 4156 11796 4168
rect 11848 4196 11854 4208
rect 12250 4196 12256 4208
rect 11848 4168 12256 4196
rect 11848 4156 11854 4168
rect 12250 4156 12256 4168
rect 12308 4156 12314 4208
rect 13446 4156 13452 4208
rect 13504 4156 13510 4208
rect 13814 4156 13820 4208
rect 13872 4196 13878 4208
rect 13872 4168 14228 4196
rect 13872 4156 13878 4168
rect 8846 4128 8852 4140
rect 8260 4100 8708 4128
rect 8807 4100 8852 4128
rect 8260 4088 8266 4100
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 10597 4131 10655 4137
rect 10597 4097 10609 4131
rect 10643 4128 10655 4131
rect 10778 4128 10784 4140
rect 10643 4100 10784 4128
rect 10643 4097 10655 4100
rect 10597 4091 10655 4097
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 11238 4128 11244 4140
rect 11199 4100 11244 4128
rect 11238 4088 11244 4100
rect 11296 4088 11302 4140
rect 12345 4131 12403 4137
rect 12345 4097 12357 4131
rect 12391 4128 12403 4131
rect 12434 4128 12440 4140
rect 12391 4100 12440 4128
rect 12391 4097 12403 4100
rect 12345 4091 12403 4097
rect 12434 4088 12440 4100
rect 12492 4088 12498 4140
rect 14200 4137 14228 4168
rect 16114 4156 16120 4208
rect 16172 4156 16178 4208
rect 14185 4131 14243 4137
rect 14185 4097 14197 4131
rect 14231 4097 14243 4131
rect 14185 4091 14243 4097
rect 14461 4131 14519 4137
rect 14461 4097 14473 4131
rect 14507 4128 14519 4131
rect 14550 4128 14556 4140
rect 14507 4100 14556 4128
rect 14507 4097 14519 4100
rect 14461 4091 14519 4097
rect 3896 4060 3924 4088
rect 3620 4032 3924 4060
rect 3973 4063 4031 4069
rect 3237 4023 3295 4029
rect 3973 4029 3985 4063
rect 4019 4029 4031 4063
rect 3973 4023 4031 4029
rect 2593 3995 2651 4001
rect 2593 3992 2605 3995
rect 1780 3964 2605 3992
rect 1118 3884 1124 3936
rect 1176 3924 1182 3936
rect 1780 3924 1808 3964
rect 2593 3961 2605 3964
rect 2639 3961 2651 3995
rect 3252 3992 3280 4023
rect 3988 3992 4016 4023
rect 4890 4020 4896 4072
rect 4948 4060 4954 4072
rect 5350 4060 5356 4072
rect 4948 4032 5356 4060
rect 4948 4020 4954 4032
rect 5350 4020 5356 4032
rect 5408 4060 5414 4072
rect 5905 4063 5963 4069
rect 5905 4060 5917 4063
rect 5408 4032 5917 4060
rect 5408 4020 5414 4032
rect 5905 4029 5917 4032
rect 5951 4029 5963 4063
rect 8938 4060 8944 4072
rect 8851 4032 8944 4060
rect 5905 4023 5963 4029
rect 8938 4020 8944 4032
rect 8996 4060 9002 4072
rect 10413 4063 10471 4069
rect 10413 4060 10425 4063
rect 8996 4032 10425 4060
rect 8996 4020 9002 4032
rect 10413 4029 10425 4032
rect 10459 4029 10471 4063
rect 11330 4060 11336 4072
rect 11291 4032 11336 4060
rect 10413 4023 10471 4029
rect 11330 4020 11336 4032
rect 11388 4020 11394 4072
rect 13170 4060 13176 4072
rect 11716 4032 13176 4060
rect 3252 3964 4016 3992
rect 11149 3995 11207 4001
rect 2593 3955 2651 3961
rect 3896 3936 3924 3964
rect 11149 3961 11161 3995
rect 11195 3992 11207 3995
rect 11716 3992 11744 4032
rect 13170 4020 13176 4032
rect 13228 4060 13234 4072
rect 13814 4060 13820 4072
rect 13228 4032 13820 4060
rect 13228 4020 13234 4032
rect 13814 4020 13820 4032
rect 13872 4020 13878 4072
rect 13909 4063 13967 4069
rect 13909 4029 13921 4063
rect 13955 4060 13967 4063
rect 14200 4060 14228 4091
rect 14550 4088 14556 4100
rect 14608 4128 14614 4140
rect 15286 4128 15292 4140
rect 14608 4100 15292 4128
rect 14608 4088 14614 4100
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 14829 4063 14887 4069
rect 14829 4060 14841 4063
rect 13955 4032 14136 4060
rect 14200 4032 14841 4060
rect 13955 4029 13967 4032
rect 13909 4023 13967 4029
rect 12894 3992 12900 4004
rect 11195 3964 11744 3992
rect 12406 3964 12900 3992
rect 11195 3961 11207 3964
rect 11149 3955 11207 3961
rect 1176 3896 1808 3924
rect 1176 3884 1182 3896
rect 2682 3884 2688 3936
rect 2740 3924 2746 3936
rect 3421 3927 3479 3933
rect 3421 3924 3433 3927
rect 2740 3896 3433 3924
rect 2740 3884 2746 3896
rect 3421 3893 3433 3896
rect 3467 3893 3479 3927
rect 3421 3887 3479 3893
rect 3878 3884 3884 3936
rect 3936 3884 3942 3936
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 4341 3927 4399 3933
rect 4341 3924 4353 3927
rect 4120 3896 4353 3924
rect 4120 3884 4126 3896
rect 4341 3893 4353 3896
rect 4387 3893 4399 3927
rect 4341 3887 4399 3893
rect 6822 3884 6828 3936
rect 6880 3924 6886 3936
rect 11698 3924 11704 3936
rect 6880 3896 11704 3924
rect 6880 3884 6886 3896
rect 11698 3884 11704 3896
rect 11756 3924 11762 3936
rect 12406 3924 12434 3964
rect 12894 3952 12900 3964
rect 12952 3952 12958 4004
rect 14108 3992 14136 4032
rect 14829 4029 14841 4032
rect 14875 4060 14887 4063
rect 15010 4060 15016 4072
rect 14875 4032 15016 4060
rect 14875 4029 14887 4032
rect 14829 4023 14887 4029
rect 15010 4020 15016 4032
rect 15068 4020 15074 4072
rect 15194 4060 15200 4072
rect 15155 4032 15200 4060
rect 15194 4020 15200 4032
rect 15252 4020 15258 4072
rect 15930 4020 15936 4072
rect 15988 4060 15994 4072
rect 16132 4060 16160 4156
rect 16574 4088 16580 4140
rect 16632 4137 16638 4140
rect 16632 4131 16681 4137
rect 16632 4097 16635 4131
rect 16669 4097 16681 4131
rect 16632 4091 16681 4097
rect 18233 4131 18291 4137
rect 18233 4097 18245 4131
rect 18279 4128 18291 4131
rect 18322 4128 18328 4140
rect 18279 4100 18328 4128
rect 18279 4097 18291 4100
rect 18233 4091 18291 4097
rect 16632 4088 16638 4091
rect 18322 4088 18328 4100
rect 18380 4088 18386 4140
rect 16390 4060 16396 4072
rect 15988 4032 16396 4060
rect 15988 4020 15994 4032
rect 16390 4020 16396 4032
rect 16448 4060 16454 4072
rect 16853 4063 16911 4069
rect 16853 4060 16865 4063
rect 16448 4032 16865 4060
rect 16448 4020 16454 4032
rect 16853 4029 16865 4032
rect 16899 4060 16911 4063
rect 17037 4063 17095 4069
rect 17037 4060 17049 4063
rect 16899 4032 17049 4060
rect 16899 4029 16911 4032
rect 16853 4023 16911 4029
rect 17037 4029 17049 4032
rect 17083 4029 17095 4063
rect 17037 4023 17095 4029
rect 18046 3992 18052 4004
rect 14108 3964 14872 3992
rect 11756 3896 12434 3924
rect 12912 3924 12940 3952
rect 14645 3927 14703 3933
rect 14645 3924 14657 3927
rect 12912 3896 14657 3924
rect 11756 3884 11762 3896
rect 14645 3893 14657 3896
rect 14691 3924 14703 3927
rect 14734 3924 14740 3936
rect 14691 3896 14740 3924
rect 14691 3893 14703 3896
rect 14645 3887 14703 3893
rect 14734 3884 14740 3896
rect 14792 3884 14798 3936
rect 14844 3924 14872 3964
rect 16132 3964 18052 3992
rect 16132 3924 16160 3964
rect 18046 3952 18052 3964
rect 18104 3952 18110 4004
rect 14844 3896 16160 3924
rect 0 3834 18860 3856
rect 0 3782 3110 3834
rect 3162 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 3302 3834
rect 3354 3782 3366 3834
rect 3418 3782 6210 3834
rect 6262 3782 6274 3834
rect 6326 3782 6338 3834
rect 6390 3782 6402 3834
rect 6454 3782 6466 3834
rect 6518 3782 9310 3834
rect 9362 3782 9374 3834
rect 9426 3782 9438 3834
rect 9490 3782 9502 3834
rect 9554 3782 9566 3834
rect 9618 3782 12410 3834
rect 12462 3782 12474 3834
rect 12526 3782 12538 3834
rect 12590 3782 12602 3834
rect 12654 3782 12666 3834
rect 12718 3782 15510 3834
rect 15562 3782 15574 3834
rect 15626 3782 15638 3834
rect 15690 3782 15702 3834
rect 15754 3782 15766 3834
rect 15818 3782 18860 3834
rect 0 3760 18860 3782
rect 842 3680 848 3732
rect 900 3720 906 3732
rect 1305 3723 1363 3729
rect 1305 3720 1317 3723
rect 900 3692 1317 3720
rect 900 3680 906 3692
rect 1305 3689 1317 3692
rect 1351 3689 1363 3723
rect 1305 3683 1363 3689
rect 3697 3723 3755 3729
rect 3697 3689 3709 3723
rect 3743 3720 3755 3723
rect 3786 3720 3792 3732
rect 3743 3692 3792 3720
rect 3743 3689 3755 3692
rect 3697 3683 3755 3689
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 5721 3723 5779 3729
rect 5721 3689 5733 3723
rect 5767 3720 5779 3723
rect 11146 3720 11152 3732
rect 5767 3692 11152 3720
rect 5767 3689 5779 3692
rect 5721 3683 5779 3689
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 11238 3680 11244 3732
rect 11296 3720 11302 3732
rect 11333 3723 11391 3729
rect 11333 3720 11345 3723
rect 11296 3692 11345 3720
rect 11296 3680 11302 3692
rect 11333 3689 11345 3692
rect 11379 3689 11391 3723
rect 11333 3683 11391 3689
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 14829 3723 14887 3729
rect 14829 3720 14841 3723
rect 12308 3692 14841 3720
rect 12308 3680 12314 3692
rect 14829 3689 14841 3692
rect 14875 3689 14887 3723
rect 14829 3683 14887 3689
rect 4522 3612 4528 3664
rect 4580 3652 4586 3664
rect 4709 3655 4767 3661
rect 4709 3652 4721 3655
rect 4580 3624 4721 3652
rect 4580 3612 4586 3624
rect 4709 3621 4721 3624
rect 4755 3621 4767 3655
rect 8202 3652 8208 3664
rect 4709 3615 4767 3621
rect 6564 3624 8208 3652
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 2924 3556 3372 3584
rect 2924 3544 2930 3556
rect 1489 3519 1547 3525
rect 1489 3485 1501 3519
rect 1535 3516 1547 3519
rect 2682 3516 2688 3528
rect 1535 3488 2688 3516
rect 1535 3485 1547 3488
rect 1489 3479 1547 3485
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 3344 3525 3372 3556
rect 3970 3544 3976 3596
rect 4028 3584 4034 3596
rect 4249 3587 4307 3593
rect 4249 3584 4261 3587
rect 4028 3556 4261 3584
rect 4028 3544 4034 3556
rect 4249 3553 4261 3556
rect 4295 3553 4307 3587
rect 6564 3584 6592 3624
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 8297 3655 8355 3661
rect 8297 3621 8309 3655
rect 8343 3652 8355 3655
rect 14844 3652 14872 3683
rect 15194 3680 15200 3732
rect 15252 3720 15258 3732
rect 18325 3723 18383 3729
rect 18325 3720 18337 3723
rect 15252 3692 18337 3720
rect 15252 3680 15258 3692
rect 18325 3689 18337 3692
rect 18371 3689 18383 3723
rect 18325 3683 18383 3689
rect 15289 3655 15347 3661
rect 15289 3652 15301 3655
rect 8343 3624 8524 3652
rect 14844 3624 15301 3652
rect 8343 3621 8355 3624
rect 8297 3615 8355 3621
rect 4249 3547 4307 3553
rect 4540 3556 6592 3584
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3485 3203 3519
rect 3145 3479 3203 3485
rect 3329 3519 3387 3525
rect 3329 3485 3341 3519
rect 3375 3485 3387 3519
rect 4062 3516 4068 3528
rect 4023 3488 4068 3516
rect 3329 3479 3387 3485
rect 2501 3383 2559 3389
rect 2501 3349 2513 3383
rect 2547 3380 2559 3383
rect 2590 3380 2596 3392
rect 2547 3352 2596 3380
rect 2547 3349 2559 3352
rect 2501 3343 2559 3349
rect 2590 3340 2596 3352
rect 2648 3340 2654 3392
rect 2682 3340 2688 3392
rect 2740 3380 2746 3392
rect 3160 3380 3188 3479
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 4540 3525 4568 3556
rect 6638 3544 6644 3596
rect 6696 3584 6702 3596
rect 6917 3587 6975 3593
rect 6917 3584 6929 3587
rect 6696 3556 6929 3584
rect 6696 3544 6702 3556
rect 6917 3553 6929 3556
rect 6963 3553 6975 3587
rect 6917 3547 6975 3553
rect 7006 3544 7012 3596
rect 7064 3584 7070 3596
rect 7837 3587 7895 3593
rect 7837 3584 7849 3587
rect 7064 3556 7849 3584
rect 7064 3544 7070 3556
rect 7837 3553 7849 3556
rect 7883 3553 7895 3587
rect 8496 3584 8524 3624
rect 15289 3621 15301 3624
rect 15335 3652 15347 3655
rect 15473 3655 15531 3661
rect 15473 3652 15485 3655
rect 15335 3624 15485 3652
rect 15335 3621 15347 3624
rect 15289 3615 15347 3621
rect 15473 3621 15485 3624
rect 15519 3621 15531 3655
rect 15473 3615 15531 3621
rect 8849 3587 8907 3593
rect 8849 3584 8861 3587
rect 8496 3556 8861 3584
rect 7837 3547 7895 3553
rect 8849 3553 8861 3556
rect 8895 3553 8907 3587
rect 8849 3547 8907 3553
rect 11149 3587 11207 3593
rect 11149 3553 11161 3587
rect 11195 3584 11207 3587
rect 11790 3584 11796 3596
rect 11195 3556 11796 3584
rect 11195 3553 11207 3556
rect 11149 3547 11207 3553
rect 11790 3544 11796 3556
rect 11848 3544 11854 3596
rect 13262 3584 13268 3596
rect 12544 3556 13268 3584
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3516 4215 3519
rect 4525 3519 4583 3525
rect 4525 3516 4537 3519
rect 4203 3488 4537 3516
rect 4203 3485 4215 3488
rect 4157 3479 4215 3485
rect 4525 3485 4537 3488
rect 4571 3485 4583 3519
rect 4890 3516 4896 3528
rect 4851 3488 4896 3516
rect 4525 3479 4583 3485
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 5258 3516 5264 3528
rect 5219 3488 5264 3516
rect 5258 3476 5264 3488
rect 5316 3476 5322 3528
rect 5810 3476 5816 3528
rect 5868 3516 5874 3528
rect 6822 3516 6828 3528
rect 5868 3488 6828 3516
rect 5868 3476 5874 3488
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 8297 3519 8355 3525
rect 8297 3485 8309 3519
rect 8343 3516 8355 3519
rect 8386 3516 8392 3528
rect 8343 3488 8392 3516
rect 8343 3485 8355 3488
rect 8297 3479 8355 3485
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 8536 3488 8581 3516
rect 8536 3476 8542 3488
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 12544 3525 12572 3556
rect 13262 3544 13268 3556
rect 13320 3544 13326 3596
rect 14734 3584 14740 3596
rect 14695 3556 14740 3584
rect 14734 3544 14740 3556
rect 14792 3544 14798 3596
rect 10275 3519 10333 3525
rect 10275 3516 10287 3519
rect 10100 3488 10287 3516
rect 10100 3476 10106 3488
rect 10275 3485 10287 3488
rect 10321 3516 10333 3519
rect 11057 3519 11115 3525
rect 11057 3516 11069 3519
rect 10321 3488 11069 3516
rect 10321 3485 10333 3488
rect 10275 3479 10333 3485
rect 11057 3485 11069 3488
rect 11103 3485 11115 3519
rect 11057 3479 11115 3485
rect 12529 3519 12587 3525
rect 12529 3485 12541 3519
rect 12575 3485 12587 3519
rect 12894 3516 12900 3528
rect 12855 3488 12900 3516
rect 12529 3479 12587 3485
rect 12894 3476 12900 3488
rect 12952 3476 12958 3528
rect 13081 3519 13139 3525
rect 13081 3485 13093 3519
rect 13127 3516 13139 3519
rect 13127 3488 14136 3516
rect 13127 3485 13139 3488
rect 13081 3479 13139 3485
rect 3237 3451 3295 3457
rect 3237 3417 3249 3451
rect 3283 3448 3295 3451
rect 4430 3448 4436 3460
rect 3283 3420 4436 3448
rect 3283 3417 3295 3420
rect 3237 3411 3295 3417
rect 4430 3408 4436 3420
rect 4488 3408 4494 3460
rect 5077 3451 5135 3457
rect 5077 3417 5089 3451
rect 5123 3448 5135 3451
rect 7006 3448 7012 3460
rect 5123 3420 7012 3448
rect 5123 3417 5135 3420
rect 5077 3411 5135 3417
rect 7006 3408 7012 3420
rect 7064 3408 7070 3460
rect 7558 3408 7564 3460
rect 7616 3448 7622 3460
rect 8021 3451 8079 3457
rect 7616 3420 7972 3448
rect 7616 3408 7622 3420
rect 2740 3352 3188 3380
rect 6365 3383 6423 3389
rect 2740 3340 2746 3352
rect 6365 3349 6377 3383
rect 6411 3380 6423 3383
rect 6546 3380 6552 3392
rect 6411 3352 6552 3380
rect 6411 3349 6423 3352
rect 6365 3343 6423 3349
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 6730 3380 6736 3392
rect 6691 3352 6736 3380
rect 6730 3340 6736 3352
rect 6788 3340 6794 3392
rect 7944 3380 7972 3420
rect 8021 3417 8033 3451
rect 8067 3448 8079 3451
rect 8110 3448 8116 3460
rect 8067 3420 8116 3448
rect 8067 3417 8079 3420
rect 8021 3411 8079 3417
rect 8110 3408 8116 3420
rect 8168 3408 8174 3460
rect 8205 3451 8263 3457
rect 8205 3417 8217 3451
rect 8251 3417 8263 3451
rect 8205 3411 8263 3417
rect 8220 3380 8248 3411
rect 9214 3408 9220 3460
rect 9272 3408 9278 3460
rect 12912 3448 12940 3476
rect 13510 3451 13568 3457
rect 13510 3448 13522 3451
rect 12912 3420 13522 3448
rect 13510 3417 13522 3420
rect 13556 3417 13568 3451
rect 13510 3411 13568 3417
rect 11698 3380 11704 3392
rect 7944 3352 11704 3380
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 12066 3340 12072 3392
rect 12124 3380 12130 3392
rect 12253 3383 12311 3389
rect 12253 3380 12265 3383
rect 12124 3352 12265 3380
rect 12124 3340 12130 3352
rect 12253 3349 12265 3352
rect 12299 3349 12311 3383
rect 12253 3343 12311 3349
rect 12989 3383 13047 3389
rect 12989 3349 13001 3383
rect 13035 3380 13047 3383
rect 13814 3380 13820 3392
rect 13035 3352 13820 3380
rect 13035 3349 13047 3352
rect 12989 3343 13047 3349
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 14108 3380 14136 3488
rect 14918 3476 14924 3528
rect 14976 3516 14982 3528
rect 15013 3519 15071 3525
rect 15013 3516 15025 3519
rect 14976 3488 15025 3516
rect 14976 3476 14982 3488
rect 15013 3485 15025 3488
rect 15059 3485 15071 3519
rect 15838 3516 15844 3528
rect 15799 3488 15844 3516
rect 15013 3479 15071 3485
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 18233 3519 18291 3525
rect 18233 3485 18245 3519
rect 18279 3516 18291 3519
rect 18506 3516 18512 3528
rect 18279 3488 18512 3516
rect 18279 3485 18291 3488
rect 18233 3479 18291 3485
rect 18506 3476 18512 3488
rect 18564 3476 18570 3528
rect 15473 3451 15531 3457
rect 15473 3417 15485 3451
rect 15519 3448 15531 3451
rect 16114 3448 16120 3460
rect 15519 3420 15976 3448
rect 16075 3420 16120 3448
rect 15519 3417 15531 3420
rect 15473 3411 15531 3417
rect 14642 3380 14648 3392
rect 14108 3352 14648 3380
rect 14642 3340 14648 3352
rect 14700 3340 14706 3392
rect 14734 3340 14740 3392
rect 14792 3380 14798 3392
rect 15197 3383 15255 3389
rect 15197 3380 15209 3383
rect 14792 3352 15209 3380
rect 14792 3340 14798 3352
rect 15197 3349 15209 3352
rect 15243 3349 15255 3383
rect 15197 3343 15255 3349
rect 15749 3383 15807 3389
rect 15749 3349 15761 3383
rect 15795 3380 15807 3383
rect 15838 3380 15844 3392
rect 15795 3352 15844 3380
rect 15795 3349 15807 3352
rect 15749 3343 15807 3349
rect 15838 3340 15844 3352
rect 15896 3340 15902 3392
rect 15948 3380 15976 3420
rect 16114 3408 16120 3420
rect 16172 3408 16178 3460
rect 16390 3408 16396 3460
rect 16448 3448 16454 3460
rect 16448 3420 16606 3448
rect 16448 3408 16454 3420
rect 17402 3408 17408 3460
rect 17460 3448 17466 3460
rect 17865 3451 17923 3457
rect 17865 3448 17877 3451
rect 17460 3420 17877 3448
rect 17460 3408 17466 3420
rect 17865 3417 17877 3420
rect 17911 3417 17923 3451
rect 17865 3411 17923 3417
rect 16850 3380 16856 3392
rect 15948 3352 16856 3380
rect 16850 3340 16856 3352
rect 16908 3340 16914 3392
rect 0 3290 18860 3312
rect 0 3238 4660 3290
rect 4712 3238 4724 3290
rect 4776 3238 4788 3290
rect 4840 3238 4852 3290
rect 4904 3238 4916 3290
rect 4968 3238 7760 3290
rect 7812 3238 7824 3290
rect 7876 3238 7888 3290
rect 7940 3238 7952 3290
rect 8004 3238 8016 3290
rect 8068 3238 10860 3290
rect 10912 3238 10924 3290
rect 10976 3238 10988 3290
rect 11040 3238 11052 3290
rect 11104 3238 11116 3290
rect 11168 3238 13960 3290
rect 14012 3238 14024 3290
rect 14076 3238 14088 3290
rect 14140 3238 14152 3290
rect 14204 3238 14216 3290
rect 14268 3238 17060 3290
rect 17112 3238 17124 3290
rect 17176 3238 17188 3290
rect 17240 3238 17252 3290
rect 17304 3238 17316 3290
rect 17368 3238 18860 3290
rect 0 3216 18860 3238
rect 1302 3176 1308 3188
rect 308 3148 1308 3176
rect 308 3049 336 3148
rect 1302 3136 1308 3148
rect 1360 3176 1366 3188
rect 6086 3176 6092 3188
rect 1360 3148 6092 3176
rect 1360 3136 1366 3148
rect 1854 3108 1860 3120
rect 1767 3080 1860 3108
rect 1854 3068 1860 3080
rect 1912 3108 1918 3120
rect 2317 3111 2375 3117
rect 2317 3108 2329 3111
rect 1912 3080 2329 3108
rect 1912 3068 1918 3080
rect 2317 3077 2329 3080
rect 2363 3077 2375 3111
rect 2317 3071 2375 3077
rect 2682 3068 2688 3120
rect 2740 3108 2746 3120
rect 2869 3111 2927 3117
rect 2869 3108 2881 3111
rect 2740 3080 2881 3108
rect 2740 3068 2746 3080
rect 2869 3077 2881 3080
rect 2915 3077 2927 3111
rect 2869 3071 2927 3077
rect 293 3043 351 3049
rect 293 3009 305 3043
rect 339 3009 351 3043
rect 293 3003 351 3009
rect 566 2972 572 2984
rect 527 2944 572 2972
rect 566 2932 572 2944
rect 624 2932 630 2984
rect 2038 2972 2044 2984
rect 1951 2944 2044 2972
rect 2038 2932 2044 2944
rect 2096 2972 2102 2984
rect 2700 2972 2728 3068
rect 5184 3052 5212 3148
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8297 3179 8355 3185
rect 8297 3176 8309 3179
rect 8168 3148 8309 3176
rect 8168 3136 8174 3148
rect 8297 3145 8309 3148
rect 8343 3145 8355 3179
rect 8297 3139 8355 3145
rect 8386 3136 8392 3188
rect 8444 3176 8450 3188
rect 8573 3179 8631 3185
rect 8573 3176 8585 3179
rect 8444 3148 8585 3176
rect 8444 3136 8450 3148
rect 8573 3145 8585 3148
rect 8619 3145 8631 3179
rect 15010 3176 15016 3188
rect 8573 3139 8631 3145
rect 8864 3148 14320 3176
rect 7006 3108 7012 3120
rect 6670 3080 7012 3108
rect 7006 3068 7012 3080
rect 7064 3068 7070 3120
rect 7300 3080 8064 3108
rect 3694 3040 3700 3052
rect 3655 3012 3700 3040
rect 3694 3000 3700 3012
rect 3752 3000 3758 3052
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 4154 3040 4160 3052
rect 3835 3012 4160 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 4338 3040 4344 3052
rect 4299 3012 4344 3040
rect 4338 3000 4344 3012
rect 4396 3000 4402 3052
rect 4522 3000 4528 3052
rect 4580 3040 4586 3052
rect 4617 3043 4675 3049
rect 4617 3040 4629 3043
rect 4580 3012 4629 3040
rect 4580 3000 4586 3012
rect 4617 3009 4629 3012
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3009 4951 3043
rect 5166 3040 5172 3052
rect 5079 3012 5172 3040
rect 4893 3003 4951 3009
rect 2096 2944 2728 2972
rect 2961 2975 3019 2981
rect 2096 2932 2102 2944
rect 2961 2941 2973 2975
rect 3007 2941 3019 2975
rect 2961 2935 3019 2941
rect 3145 2975 3203 2981
rect 3145 2941 3157 2975
rect 3191 2972 3203 2975
rect 3602 2972 3608 2984
rect 3191 2944 3608 2972
rect 3191 2941 3203 2944
rect 3145 2935 3203 2941
rect 2501 2907 2559 2913
rect 2501 2904 2513 2907
rect 1596 2876 2513 2904
rect 934 2796 940 2848
rect 992 2836 998 2848
rect 1596 2836 1624 2876
rect 2501 2873 2513 2876
rect 2547 2873 2559 2907
rect 2976 2904 3004 2935
rect 3602 2932 3608 2944
rect 3660 2932 3666 2984
rect 3970 2972 3976 2984
rect 3931 2944 3976 2972
rect 3970 2932 3976 2944
rect 4028 2932 4034 2984
rect 4908 2972 4936 3003
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 7300 3049 7328 3080
rect 8036 3052 8064 3080
rect 7285 3043 7343 3049
rect 7285 3009 7297 3043
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3009 7435 3043
rect 7558 3040 7564 3052
rect 7519 3012 7564 3040
rect 7377 3003 7435 3009
rect 5445 2975 5503 2981
rect 4908 2944 5304 2972
rect 3329 2907 3387 2913
rect 3329 2904 3341 2907
rect 2976 2876 3341 2904
rect 2501 2867 2559 2873
rect 3329 2873 3341 2876
rect 3375 2873 3387 2907
rect 3329 2867 3387 2873
rect 992 2808 1624 2836
rect 2225 2839 2283 2845
rect 992 2796 998 2808
rect 2225 2805 2237 2839
rect 2271 2836 2283 2839
rect 2317 2839 2375 2845
rect 2317 2836 2329 2839
rect 2271 2808 2329 2836
rect 2271 2805 2283 2808
rect 2225 2799 2283 2805
rect 2317 2805 2329 2808
rect 2363 2836 2375 2839
rect 2590 2836 2596 2848
rect 2363 2808 2596 2836
rect 2363 2805 2375 2808
rect 2317 2799 2375 2805
rect 2590 2796 2596 2808
rect 2648 2796 2654 2848
rect 4522 2836 4528 2848
rect 4483 2808 4528 2836
rect 4522 2796 4528 2808
rect 4580 2796 4586 2848
rect 5074 2836 5080 2848
rect 5035 2808 5080 2836
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 5276 2836 5304 2944
rect 5445 2941 5457 2975
rect 5491 2972 5503 2975
rect 6086 2972 6092 2984
rect 5491 2944 6092 2972
rect 5491 2941 5503 2944
rect 5445 2935 5503 2941
rect 6086 2932 6092 2944
rect 6144 2932 6150 2984
rect 6914 2972 6920 2984
rect 6827 2944 6920 2972
rect 6914 2932 6920 2944
rect 6972 2972 6978 2984
rect 7392 2972 7420 3003
rect 7558 3000 7564 3012
rect 7616 3000 7622 3052
rect 8018 3040 8024 3052
rect 7979 3012 8024 3040
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3040 8263 3043
rect 8662 3040 8668 3052
rect 8251 3012 8668 3040
rect 8251 3009 8263 3012
rect 8205 3003 8263 3009
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 8864 3049 8892 3148
rect 11885 3111 11943 3117
rect 11885 3077 11897 3111
rect 11931 3108 11943 3111
rect 11931 3080 12204 3108
rect 11931 3077 11943 3080
rect 11885 3071 11943 3077
rect 8757 3043 8815 3049
rect 8757 3009 8769 3043
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 8849 3043 8907 3049
rect 8849 3009 8861 3043
rect 8895 3009 8907 3043
rect 8849 3003 8907 3009
rect 6972 2944 7420 2972
rect 8481 2975 8539 2981
rect 6972 2932 6978 2944
rect 8481 2941 8493 2975
rect 8527 2972 8539 2975
rect 8772 2972 8800 3003
rect 8938 3000 8944 3052
rect 8996 3040 9002 3052
rect 9861 3043 9919 3049
rect 8996 3012 9041 3040
rect 8996 3000 9002 3012
rect 9861 3009 9873 3043
rect 9907 3040 9919 3043
rect 10042 3040 10048 3052
rect 9907 3012 10048 3040
rect 9907 3009 9919 3012
rect 9861 3003 9919 3009
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 12066 3040 12072 3052
rect 12027 3012 12072 3040
rect 12066 3000 12072 3012
rect 12124 3000 12130 3052
rect 12176 3040 12204 3080
rect 13446 3068 13452 3120
rect 13504 3068 13510 3120
rect 12526 3040 12532 3052
rect 12176 3012 12532 3040
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 9769 2975 9827 2981
rect 9769 2972 9781 2975
rect 8527 2944 9781 2972
rect 8527 2941 8539 2944
rect 8481 2935 8539 2941
rect 9769 2941 9781 2944
rect 9815 2941 9827 2975
rect 9769 2935 9827 2941
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 12802 2972 12808 2984
rect 12483 2944 12808 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 12802 2932 12808 2944
rect 12860 2932 12866 2984
rect 12986 2932 12992 2984
rect 13044 2972 13050 2984
rect 13464 2972 13492 3068
rect 13814 3000 13820 3052
rect 13872 3040 13878 3052
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 13872 3012 14013 3040
rect 13872 3000 13878 3012
rect 14001 3009 14013 3012
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 14292 2981 14320 3148
rect 14936 3148 15016 3176
rect 14642 3040 14648 3052
rect 14603 3012 14648 3040
rect 14642 3000 14648 3012
rect 14700 3000 14706 3052
rect 14826 3040 14832 3052
rect 14787 3012 14832 3040
rect 14826 3000 14832 3012
rect 14884 3000 14890 3052
rect 14936 3049 14964 3148
rect 15010 3136 15016 3148
rect 15068 3136 15074 3188
rect 16114 3136 16120 3188
rect 16172 3176 16178 3188
rect 16669 3179 16727 3185
rect 16669 3176 16681 3179
rect 16172 3148 16681 3176
rect 16172 3136 16178 3148
rect 16669 3145 16681 3148
rect 16715 3145 16727 3179
rect 16669 3139 16727 3145
rect 15838 3068 15844 3120
rect 15896 3068 15902 3120
rect 14921 3043 14979 3049
rect 14921 3009 14933 3043
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 16850 3000 16856 3052
rect 16908 3040 16914 3052
rect 17037 3043 17095 3049
rect 17037 3040 17049 3043
rect 16908 3012 17049 3040
rect 16908 3000 16914 3012
rect 17037 3009 17049 3012
rect 17083 3040 17095 3043
rect 17589 3043 17647 3049
rect 17589 3040 17601 3043
rect 17083 3012 17601 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 17589 3009 17601 3012
rect 17635 3040 17647 3043
rect 17770 3040 17776 3052
rect 17635 3012 17776 3040
rect 17635 3009 17647 3012
rect 17589 3003 17647 3009
rect 17770 3000 17776 3012
rect 17828 3000 17834 3052
rect 13044 2944 13492 2972
rect 14277 2975 14335 2981
rect 13044 2932 13050 2944
rect 14277 2941 14289 2975
rect 14323 2972 14335 2975
rect 14734 2972 14740 2984
rect 14323 2944 14740 2972
rect 14323 2941 14335 2944
rect 14277 2935 14335 2941
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 15197 2975 15255 2981
rect 15197 2941 15209 2975
rect 15243 2972 15255 2975
rect 17678 2972 17684 2984
rect 15243 2944 17684 2972
rect 15243 2941 15255 2944
rect 15197 2935 15255 2941
rect 17678 2932 17684 2944
rect 17736 2932 17742 2984
rect 6822 2864 6828 2916
rect 6880 2904 6886 2916
rect 7285 2907 7343 2913
rect 7285 2904 7297 2907
rect 6880 2876 7297 2904
rect 6880 2864 6886 2876
rect 7285 2873 7297 2876
rect 7331 2873 7343 2907
rect 7285 2867 7343 2873
rect 8662 2864 8668 2916
rect 8720 2904 8726 2916
rect 8938 2904 8944 2916
rect 8720 2876 8944 2904
rect 8720 2864 8726 2876
rect 8938 2864 8944 2876
rect 8996 2864 9002 2916
rect 14093 2907 14151 2913
rect 14093 2873 14105 2907
rect 14139 2904 14151 2907
rect 14461 2907 14519 2913
rect 14461 2904 14473 2907
rect 14139 2876 14473 2904
rect 14139 2873 14151 2876
rect 14093 2867 14151 2873
rect 14461 2873 14473 2876
rect 14507 2873 14519 2907
rect 14461 2867 14519 2873
rect 16390 2864 16396 2916
rect 16448 2904 16454 2916
rect 16853 2907 16911 2913
rect 16853 2904 16865 2907
rect 16448 2876 16865 2904
rect 16448 2864 16454 2876
rect 16853 2873 16865 2876
rect 16899 2873 16911 2907
rect 16853 2867 16911 2873
rect 17497 2907 17555 2913
rect 17497 2873 17509 2907
rect 17543 2904 17555 2907
rect 18138 2904 18144 2916
rect 17543 2876 18144 2904
rect 17543 2873 17555 2876
rect 17497 2867 17555 2873
rect 18138 2864 18144 2876
rect 18196 2864 18202 2916
rect 7190 2836 7196 2848
rect 5276 2808 7196 2836
rect 7190 2796 7196 2808
rect 7248 2796 7254 2848
rect 11790 2796 11796 2848
rect 11848 2836 11854 2848
rect 11974 2836 11980 2848
rect 11848 2808 11980 2836
rect 11848 2796 11854 2808
rect 11974 2796 11980 2808
rect 12032 2836 12038 2848
rect 13863 2839 13921 2845
rect 13863 2836 13875 2839
rect 12032 2808 13875 2836
rect 12032 2796 12038 2808
rect 13863 2805 13875 2808
rect 13909 2805 13921 2839
rect 13863 2799 13921 2805
rect 14185 2839 14243 2845
rect 14185 2805 14197 2839
rect 14231 2836 14243 2839
rect 14366 2836 14372 2848
rect 14231 2808 14372 2836
rect 14231 2805 14243 2808
rect 14185 2799 14243 2805
rect 14366 2796 14372 2808
rect 14424 2796 14430 2848
rect 17126 2836 17132 2848
rect 17087 2808 17132 2836
rect 17126 2796 17132 2808
rect 17184 2796 17190 2848
rect 17862 2796 17868 2848
rect 17920 2836 17926 2848
rect 17957 2839 18015 2845
rect 17957 2836 17969 2839
rect 17920 2808 17969 2836
rect 17920 2796 17926 2808
rect 17957 2805 17969 2808
rect 18003 2805 18015 2839
rect 17957 2799 18015 2805
rect 0 2746 18860 2768
rect 0 2694 3110 2746
rect 3162 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 3302 2746
rect 3354 2694 3366 2746
rect 3418 2694 6210 2746
rect 6262 2694 6274 2746
rect 6326 2694 6338 2746
rect 6390 2694 6402 2746
rect 6454 2694 6466 2746
rect 6518 2694 9310 2746
rect 9362 2694 9374 2746
rect 9426 2694 9438 2746
rect 9490 2694 9502 2746
rect 9554 2694 9566 2746
rect 9618 2694 12410 2746
rect 12462 2694 12474 2746
rect 12526 2694 12538 2746
rect 12590 2694 12602 2746
rect 12654 2694 12666 2746
rect 12718 2694 15510 2746
rect 15562 2694 15574 2746
rect 15626 2694 15638 2746
rect 15690 2694 15702 2746
rect 15754 2694 15766 2746
rect 15818 2694 18860 2746
rect 0 2672 18860 2694
rect 566 2592 572 2644
rect 624 2632 630 2644
rect 753 2635 811 2641
rect 753 2632 765 2635
rect 624 2604 765 2632
rect 624 2592 630 2604
rect 753 2601 765 2604
rect 799 2601 811 2635
rect 753 2595 811 2601
rect 2409 2635 2467 2641
rect 2409 2601 2421 2635
rect 2455 2632 2467 2635
rect 3694 2632 3700 2644
rect 2455 2604 3700 2632
rect 2455 2601 2467 2604
rect 2409 2595 2467 2601
rect 3694 2592 3700 2604
rect 3752 2592 3758 2644
rect 3789 2635 3847 2641
rect 3789 2601 3801 2635
rect 3835 2632 3847 2635
rect 3878 2632 3884 2644
rect 3835 2604 3884 2632
rect 3835 2601 3847 2604
rect 3789 2595 3847 2601
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 4522 2592 4528 2644
rect 4580 2592 4586 2644
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 5350 2632 5356 2644
rect 4764 2604 5356 2632
rect 4764 2592 4770 2604
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 6086 2632 6092 2644
rect 6047 2604 6092 2632
rect 6086 2592 6092 2604
rect 6144 2592 6150 2644
rect 6730 2592 6736 2644
rect 6788 2632 6794 2644
rect 6825 2635 6883 2641
rect 6825 2632 6837 2635
rect 6788 2604 6837 2632
rect 6788 2592 6794 2604
rect 6825 2601 6837 2604
rect 6871 2601 6883 2635
rect 8481 2635 8539 2641
rect 8481 2632 8493 2635
rect 6825 2595 6883 2601
rect 6932 2604 8493 2632
rect 3510 2524 3516 2576
rect 3568 2564 3574 2576
rect 4540 2564 4568 2592
rect 6932 2564 6960 2604
rect 8481 2601 8493 2604
rect 8527 2601 8539 2635
rect 8481 2595 8539 2601
rect 8846 2592 8852 2644
rect 8904 2632 8910 2644
rect 9585 2635 9643 2641
rect 9585 2632 9597 2635
rect 8904 2604 9597 2632
rect 8904 2592 8910 2604
rect 9585 2601 9597 2604
rect 9631 2601 9643 2635
rect 9585 2595 9643 2601
rect 10042 2592 10048 2644
rect 10100 2632 10106 2644
rect 11330 2632 11336 2644
rect 10100 2604 11336 2632
rect 10100 2592 10106 2604
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 11609 2635 11667 2641
rect 11609 2601 11621 2635
rect 11655 2632 11667 2635
rect 12802 2632 12808 2644
rect 11655 2604 12808 2632
rect 11655 2601 11667 2604
rect 11609 2595 11667 2601
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 12986 2592 12992 2644
rect 13044 2632 13050 2644
rect 13357 2635 13415 2641
rect 13357 2632 13369 2635
rect 13044 2604 13369 2632
rect 13044 2592 13050 2604
rect 13357 2601 13369 2604
rect 13403 2632 13415 2635
rect 15102 2632 15108 2644
rect 13403 2604 15108 2632
rect 13403 2601 13415 2604
rect 13357 2595 13415 2601
rect 15102 2592 15108 2604
rect 15160 2592 15166 2644
rect 17037 2635 17095 2641
rect 17037 2601 17049 2635
rect 17083 2632 17095 2635
rect 17126 2632 17132 2644
rect 17083 2604 17132 2632
rect 17083 2601 17095 2604
rect 17037 2595 17095 2601
rect 17126 2592 17132 2604
rect 17184 2592 17190 2644
rect 17221 2635 17279 2641
rect 17221 2601 17233 2635
rect 17267 2601 17279 2635
rect 17678 2632 17684 2644
rect 17639 2604 17684 2632
rect 17221 2595 17279 2601
rect 3568 2536 4568 2564
rect 4908 2536 6960 2564
rect 3568 2524 3574 2536
rect 2133 2499 2191 2505
rect 2133 2465 2145 2499
rect 2179 2496 2191 2499
rect 2222 2496 2228 2508
rect 2179 2468 2228 2496
rect 2179 2465 2191 2468
rect 2133 2459 2191 2465
rect 2222 2456 2228 2468
rect 2280 2456 2286 2508
rect 2774 2456 2780 2508
rect 2832 2496 2838 2508
rect 3421 2499 3479 2505
rect 2832 2468 2877 2496
rect 2832 2456 2838 2468
rect 3421 2465 3433 2499
rect 3467 2496 3479 2499
rect 4338 2496 4344 2508
rect 3467 2468 4344 2496
rect 3467 2465 3479 2468
rect 3421 2459 3479 2465
rect 4338 2456 4344 2468
rect 4396 2496 4402 2508
rect 4908 2496 4936 2536
rect 7650 2524 7656 2576
rect 7708 2564 7714 2576
rect 8018 2564 8024 2576
rect 7708 2536 8024 2564
rect 7708 2524 7714 2536
rect 8018 2524 8024 2536
rect 8076 2564 8082 2576
rect 10060 2564 10088 2592
rect 13170 2564 13176 2576
rect 8076 2536 10088 2564
rect 10152 2536 13176 2564
rect 8076 2524 8082 2536
rect 4396 2468 4936 2496
rect 4396 2456 4402 2468
rect 934 2428 940 2440
rect 895 2400 940 2428
rect 934 2388 940 2400
rect 992 2388 998 2440
rect 2038 2428 2044 2440
rect 1999 2400 2044 2428
rect 2038 2388 2044 2400
rect 2096 2388 2102 2440
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2428 2743 2431
rect 2866 2428 2872 2440
rect 2731 2400 2872 2428
rect 2731 2397 2743 2400
rect 2685 2391 2743 2397
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 3510 2428 3516 2440
rect 3471 2400 3516 2428
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2397 4307 2431
rect 4522 2428 4528 2440
rect 4483 2400 4528 2428
rect 4249 2391 4307 2397
rect 2958 2320 2964 2372
rect 3016 2360 3022 2372
rect 3237 2363 3295 2369
rect 3237 2360 3249 2363
rect 3016 2332 3249 2360
rect 3016 2320 3022 2332
rect 3237 2329 3249 2332
rect 3283 2360 3295 2363
rect 4264 2360 4292 2391
rect 4522 2388 4528 2400
rect 4580 2388 4586 2440
rect 4706 2428 4712 2440
rect 4667 2400 4712 2428
rect 4706 2388 4712 2400
rect 4764 2388 4770 2440
rect 4908 2437 4936 2468
rect 6365 2499 6423 2505
rect 6365 2465 6377 2499
rect 6411 2496 6423 2499
rect 6546 2496 6552 2508
rect 6411 2468 6552 2496
rect 6411 2465 6423 2468
rect 6365 2459 6423 2465
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 6822 2496 6828 2508
rect 6779 2468 6828 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 6822 2456 6828 2468
rect 6880 2456 6886 2508
rect 7469 2499 7527 2505
rect 7116 2468 7420 2496
rect 4801 2431 4859 2437
rect 4801 2397 4813 2431
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 4614 2360 4620 2372
rect 3283 2332 4620 2360
rect 3283 2329 3295 2332
rect 3237 2323 3295 2329
rect 4614 2320 4620 2332
rect 4672 2320 4678 2372
rect 4816 2360 4844 2391
rect 5920 2360 5948 2391
rect 5994 2388 6000 2440
rect 6052 2428 6058 2440
rect 6273 2431 6331 2437
rect 6273 2428 6285 2431
rect 6052 2400 6285 2428
rect 6052 2388 6058 2400
rect 6273 2397 6285 2400
rect 6319 2428 6331 2431
rect 7116 2428 7144 2468
rect 6319 2400 7144 2428
rect 6319 2397 6331 2400
rect 6273 2391 6331 2397
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 7285 2431 7343 2437
rect 7285 2428 7297 2431
rect 7248 2400 7297 2428
rect 7248 2388 7254 2400
rect 7285 2397 7297 2400
rect 7331 2397 7343 2431
rect 7392 2428 7420 2468
rect 7469 2465 7481 2499
rect 7515 2496 7527 2499
rect 8573 2499 8631 2505
rect 8573 2496 8585 2499
rect 7515 2468 8585 2496
rect 7515 2465 7527 2468
rect 7469 2459 7527 2465
rect 8573 2465 8585 2468
rect 8619 2496 8631 2499
rect 9030 2496 9036 2508
rect 8619 2468 9036 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 9030 2456 9036 2468
rect 9088 2456 9094 2508
rect 9214 2456 9220 2508
rect 9272 2496 9278 2508
rect 10152 2496 10180 2536
rect 13170 2524 13176 2536
rect 13228 2524 13234 2576
rect 17236 2564 17264 2595
rect 17678 2592 17684 2604
rect 17736 2592 17742 2644
rect 17770 2564 17776 2576
rect 16960 2536 17776 2564
rect 9272 2468 10180 2496
rect 10980 2468 11468 2496
rect 9272 2456 9278 2468
rect 8110 2428 8116 2440
rect 7392 2400 8116 2428
rect 7285 2391 7343 2397
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 8662 2428 8668 2440
rect 8623 2400 8668 2428
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 9490 2388 9496 2440
rect 9548 2428 9554 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9548 2400 9781 2428
rect 9548 2388 9554 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 9306 2360 9312 2372
rect 4816 2332 9312 2360
rect 3053 2295 3111 2301
rect 3053 2261 3065 2295
rect 3099 2292 3111 2295
rect 3418 2292 3424 2304
rect 3099 2264 3424 2292
rect 3099 2261 3111 2264
rect 3053 2255 3111 2261
rect 3418 2252 3424 2264
rect 3476 2252 3482 2304
rect 3513 2295 3571 2301
rect 3513 2261 3525 2295
rect 3559 2292 3571 2295
rect 4338 2292 4344 2304
rect 3559 2264 4344 2292
rect 3559 2261 3571 2264
rect 3513 2255 3571 2261
rect 4338 2252 4344 2264
rect 4396 2252 4402 2304
rect 4430 2252 4436 2304
rect 4488 2292 4494 2304
rect 4816 2292 4844 2332
rect 9306 2320 9312 2332
rect 9364 2320 9370 2372
rect 10980 2360 11008 2468
rect 11057 2431 11115 2437
rect 11057 2397 11069 2431
rect 11103 2428 11115 2431
rect 11238 2428 11244 2440
rect 11103 2400 11244 2428
rect 11103 2397 11115 2400
rect 11057 2391 11115 2397
rect 11238 2388 11244 2400
rect 11296 2388 11302 2440
rect 11440 2437 11468 2468
rect 13262 2456 13268 2508
rect 13320 2496 13326 2508
rect 13449 2499 13507 2505
rect 13449 2496 13461 2499
rect 13320 2468 13461 2496
rect 13320 2456 13326 2468
rect 13449 2465 13461 2468
rect 13495 2496 13507 2499
rect 13722 2496 13728 2508
rect 13495 2468 13728 2496
rect 13495 2465 13507 2468
rect 13449 2459 13507 2465
rect 13722 2456 13728 2468
rect 13780 2496 13786 2508
rect 15657 2499 15715 2505
rect 15657 2496 15669 2499
rect 13780 2468 15669 2496
rect 13780 2456 13786 2468
rect 15657 2465 15669 2468
rect 15703 2465 15715 2499
rect 15657 2459 15715 2465
rect 11425 2431 11483 2437
rect 11425 2397 11437 2431
rect 11471 2397 11483 2431
rect 11974 2428 11980 2440
rect 11935 2400 11980 2428
rect 11425 2391 11483 2397
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 15102 2428 15108 2440
rect 14858 2400 15108 2428
rect 15102 2388 15108 2400
rect 15160 2388 15166 2440
rect 15924 2431 15982 2437
rect 15924 2397 15936 2431
rect 15970 2428 15982 2431
rect 16960 2428 16988 2536
rect 17770 2524 17776 2536
rect 17828 2564 17834 2576
rect 18417 2567 18475 2573
rect 18417 2564 18429 2567
rect 17828 2536 18429 2564
rect 17828 2524 17834 2536
rect 18417 2533 18429 2536
rect 18463 2533 18475 2567
rect 18417 2527 18475 2533
rect 17589 2499 17647 2505
rect 17589 2465 17601 2499
rect 17635 2496 17647 2499
rect 17635 2468 18092 2496
rect 17635 2465 17647 2468
rect 17589 2459 17647 2465
rect 17126 2428 17132 2440
rect 15970 2400 16988 2428
rect 17087 2400 17132 2428
rect 15970 2397 15982 2400
rect 15924 2391 15982 2397
rect 17126 2388 17132 2400
rect 17184 2388 17190 2440
rect 17862 2428 17868 2440
rect 17823 2400 17868 2428
rect 17862 2388 17868 2400
rect 17920 2388 17926 2440
rect 18064 2437 18092 2468
rect 18049 2431 18107 2437
rect 18049 2397 18061 2431
rect 18095 2397 18107 2431
rect 18049 2391 18107 2397
rect 18138 2388 18144 2440
rect 18196 2428 18202 2440
rect 18196 2400 18241 2428
rect 18196 2388 18202 2400
rect 11149 2363 11207 2369
rect 10980 2332 11100 2360
rect 4488 2264 4844 2292
rect 5169 2295 5227 2301
rect 4488 2252 4494 2264
rect 5169 2261 5181 2295
rect 5215 2292 5227 2295
rect 5258 2292 5264 2304
rect 5215 2264 5264 2292
rect 5215 2261 5227 2264
rect 5169 2255 5227 2261
rect 5258 2252 5264 2264
rect 5316 2252 5322 2304
rect 5442 2292 5448 2304
rect 5403 2264 5448 2292
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 7006 2252 7012 2304
rect 7064 2292 7070 2304
rect 7193 2295 7251 2301
rect 7193 2292 7205 2295
rect 7064 2264 7205 2292
rect 7064 2252 7070 2264
rect 7193 2261 7205 2264
rect 7239 2261 7251 2295
rect 7193 2255 7251 2261
rect 8481 2295 8539 2301
rect 8481 2261 8493 2295
rect 8527 2292 8539 2295
rect 9214 2292 9220 2304
rect 8527 2264 9220 2292
rect 8527 2261 8539 2264
rect 8481 2255 8539 2261
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 11072 2301 11100 2332
rect 11149 2329 11161 2363
rect 11195 2329 11207 2363
rect 11330 2360 11336 2372
rect 11291 2332 11336 2360
rect 11149 2323 11207 2329
rect 11057 2295 11115 2301
rect 11057 2261 11069 2295
rect 11103 2261 11115 2295
rect 11164 2292 11192 2323
rect 11330 2320 11336 2332
rect 11388 2320 11394 2372
rect 11517 2363 11575 2369
rect 11517 2329 11529 2363
rect 11563 2360 11575 2363
rect 11606 2360 11612 2372
rect 11563 2332 11612 2360
rect 11563 2329 11575 2332
rect 11517 2323 11575 2329
rect 11606 2320 11612 2332
rect 11664 2320 11670 2372
rect 11698 2320 11704 2372
rect 11756 2360 11762 2372
rect 13725 2363 13783 2369
rect 11756 2332 11801 2360
rect 11756 2320 11762 2332
rect 13725 2329 13737 2363
rect 13771 2360 13783 2363
rect 13814 2360 13820 2372
rect 13771 2332 13820 2360
rect 13771 2329 13783 2332
rect 13725 2323 13783 2329
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 15470 2360 15476 2372
rect 15431 2332 15476 2360
rect 15470 2320 15476 2332
rect 15528 2320 15534 2372
rect 18230 2320 18236 2372
rect 18288 2360 18294 2372
rect 18325 2363 18383 2369
rect 18325 2360 18337 2363
rect 18288 2332 18337 2360
rect 18288 2320 18294 2332
rect 18325 2329 18337 2332
rect 18371 2329 18383 2363
rect 18325 2323 18383 2329
rect 11422 2292 11428 2304
rect 11164 2264 11428 2292
rect 11057 2255 11115 2261
rect 11422 2252 11428 2264
rect 11480 2292 11486 2304
rect 11885 2295 11943 2301
rect 11885 2292 11897 2295
rect 11480 2264 11897 2292
rect 11480 2252 11486 2264
rect 11885 2261 11897 2264
rect 11931 2261 11943 2295
rect 11885 2255 11943 2261
rect 14458 2252 14464 2304
rect 14516 2292 14522 2304
rect 18049 2295 18107 2301
rect 18049 2292 18061 2295
rect 14516 2264 18061 2292
rect 14516 2252 14522 2264
rect 18049 2261 18061 2264
rect 18095 2261 18107 2295
rect 18049 2255 18107 2261
rect 0 2202 18860 2224
rect 0 2150 4660 2202
rect 4712 2150 4724 2202
rect 4776 2150 4788 2202
rect 4840 2150 4852 2202
rect 4904 2150 4916 2202
rect 4968 2150 7760 2202
rect 7812 2150 7824 2202
rect 7876 2150 7888 2202
rect 7940 2150 7952 2202
rect 8004 2150 8016 2202
rect 8068 2150 10860 2202
rect 10912 2150 10924 2202
rect 10976 2150 10988 2202
rect 11040 2150 11052 2202
rect 11104 2150 11116 2202
rect 11168 2150 13960 2202
rect 14012 2150 14024 2202
rect 14076 2150 14088 2202
rect 14140 2150 14152 2202
rect 14204 2150 14216 2202
rect 14268 2150 17060 2202
rect 17112 2150 17124 2202
rect 17176 2150 17188 2202
rect 17240 2150 17252 2202
rect 17304 2150 17316 2202
rect 17368 2150 18860 2202
rect 0 2128 18860 2150
rect 2222 2088 2228 2100
rect 2183 2060 2228 2088
rect 2222 2048 2228 2060
rect 2280 2048 2286 2100
rect 2501 2091 2559 2097
rect 2501 2057 2513 2091
rect 2547 2057 2559 2091
rect 2866 2088 2872 2100
rect 2827 2060 2872 2088
rect 2501 2051 2559 2057
rect 2516 2020 2544 2051
rect 2866 2048 2872 2060
rect 2924 2048 2930 2100
rect 2961 2091 3019 2097
rect 2961 2057 2973 2091
rect 3007 2088 3019 2091
rect 3329 2091 3387 2097
rect 3329 2088 3341 2091
rect 3007 2060 3341 2088
rect 3007 2057 3019 2060
rect 2961 2051 3019 2057
rect 3329 2057 3341 2060
rect 3375 2057 3387 2091
rect 3329 2051 3387 2057
rect 3418 2048 3424 2100
rect 3476 2088 3482 2100
rect 3697 2091 3755 2097
rect 3697 2088 3709 2091
rect 3476 2060 3709 2088
rect 3476 2048 3482 2060
rect 3697 2057 3709 2060
rect 3743 2057 3755 2091
rect 3697 2051 3755 2057
rect 7098 2048 7104 2100
rect 7156 2088 7162 2100
rect 7745 2091 7803 2097
rect 7745 2088 7757 2091
rect 7156 2060 7757 2088
rect 7156 2048 7162 2060
rect 7745 2057 7757 2060
rect 7791 2088 7803 2091
rect 8202 2088 8208 2100
rect 7791 2060 8208 2088
rect 7791 2057 7803 2060
rect 7745 2051 7803 2057
rect 8202 2048 8208 2060
rect 8260 2048 8266 2100
rect 8573 2091 8631 2097
rect 8573 2057 8585 2091
rect 8619 2088 8631 2091
rect 8662 2088 8668 2100
rect 8619 2060 8668 2088
rect 8619 2057 8631 2060
rect 8573 2051 8631 2057
rect 8662 2048 8668 2060
rect 8720 2048 8726 2100
rect 9306 2088 9312 2100
rect 9219 2060 9312 2088
rect 9306 2048 9312 2060
rect 9364 2088 9370 2100
rect 11238 2088 11244 2100
rect 9364 2060 11244 2088
rect 9364 2048 9370 2060
rect 11238 2048 11244 2060
rect 11296 2048 11302 2100
rect 11606 2088 11612 2100
rect 11567 2060 11612 2088
rect 11606 2048 11612 2060
rect 11664 2048 11670 2100
rect 13170 2088 13176 2100
rect 13083 2060 13176 2088
rect 13170 2048 13176 2060
rect 13228 2088 13234 2100
rect 13814 2088 13820 2100
rect 13228 2060 13676 2088
rect 13775 2060 13820 2088
rect 13228 2048 13234 2060
rect 1044 1992 2544 2020
rect 3789 2023 3847 2029
rect 1044 1961 1072 1992
rect 3789 1989 3801 2023
rect 3835 2020 3847 2023
rect 4249 2023 4307 2029
rect 4249 2020 4261 2023
rect 3835 1992 4261 2020
rect 3835 1989 3847 1992
rect 3789 1983 3847 1989
rect 4249 1989 4261 1992
rect 4295 1989 4307 2023
rect 4249 1983 4307 1989
rect 4522 1980 4528 2032
rect 4580 2020 4586 2032
rect 6914 2020 6920 2032
rect 4580 1992 6040 2020
rect 4580 1980 4586 1992
rect 1029 1955 1087 1961
rect 1029 1921 1041 1955
rect 1075 1921 1087 1955
rect 1029 1915 1087 1921
rect 2139 1955 2197 1961
rect 2139 1921 2151 1955
rect 2185 1952 2197 1955
rect 2317 1955 2375 1961
rect 2185 1924 2268 1952
rect 2185 1921 2197 1924
rect 2139 1915 2197 1921
rect 2240 1896 2268 1924
rect 2317 1921 2329 1955
rect 2363 1952 2375 1955
rect 2774 1952 2780 1964
rect 2363 1924 2780 1952
rect 2363 1921 2375 1924
rect 2317 1915 2375 1921
rect 2774 1912 2780 1924
rect 2832 1912 2838 1964
rect 4154 1952 4160 1964
rect 4115 1924 4160 1952
rect 4154 1912 4160 1924
rect 4212 1912 4218 1964
rect 4338 1952 4344 1964
rect 4299 1924 4344 1952
rect 4338 1912 4344 1924
rect 4396 1912 4402 1964
rect 4430 1912 4436 1964
rect 4488 1952 4494 1964
rect 4617 1955 4675 1961
rect 4617 1952 4629 1955
rect 4488 1924 4629 1952
rect 4488 1912 4494 1924
rect 4617 1921 4629 1924
rect 4663 1921 4675 1955
rect 5074 1952 5080 1964
rect 5035 1924 5080 1952
rect 4617 1915 4675 1921
rect 5074 1912 5080 1924
rect 5132 1912 5138 1964
rect 5442 1952 5448 1964
rect 5403 1924 5448 1952
rect 5442 1912 5448 1924
rect 5500 1912 5506 1964
rect 6012 1961 6040 1992
rect 6656 1992 6920 2020
rect 6656 1961 6684 1992
rect 6914 1980 6920 1992
rect 6972 2020 6978 2032
rect 8297 2023 8355 2029
rect 6972 1992 8248 2020
rect 6972 1980 6978 1992
rect 5997 1955 6055 1961
rect 5997 1921 6009 1955
rect 6043 1921 6055 1955
rect 5997 1915 6055 1921
rect 6641 1955 6699 1961
rect 6641 1921 6653 1955
rect 6687 1921 6699 1955
rect 7282 1952 7288 1964
rect 7243 1924 7288 1952
rect 6641 1915 6699 1921
rect 7282 1912 7288 1924
rect 7340 1912 7346 1964
rect 7377 1955 7435 1961
rect 7377 1921 7389 1955
rect 7423 1921 7435 1955
rect 7377 1915 7435 1921
rect 7561 1955 7619 1961
rect 7561 1921 7573 1955
rect 7607 1921 7619 1955
rect 7561 1915 7619 1921
rect 2222 1844 2228 1896
rect 2280 1884 2286 1896
rect 2866 1884 2872 1896
rect 2280 1856 2872 1884
rect 2280 1844 2286 1856
rect 2866 1844 2872 1856
rect 2924 1844 2930 1896
rect 3145 1887 3203 1893
rect 3145 1853 3157 1887
rect 3191 1884 3203 1887
rect 3602 1884 3608 1896
rect 3191 1856 3608 1884
rect 3191 1853 3203 1856
rect 3145 1847 3203 1853
rect 3602 1844 3608 1856
rect 3660 1844 3666 1896
rect 3970 1884 3976 1896
rect 3931 1856 3976 1884
rect 3970 1844 3976 1856
rect 4028 1844 4034 1896
rect 5810 1884 5816 1896
rect 5771 1856 5816 1884
rect 5810 1844 5816 1856
rect 5868 1844 5874 1896
rect 5902 1844 5908 1896
rect 5960 1884 5966 1896
rect 6549 1887 6607 1893
rect 6549 1884 6561 1887
rect 5960 1856 6561 1884
rect 5960 1844 5966 1856
rect 6549 1853 6561 1856
rect 6595 1853 6607 1887
rect 7006 1884 7012 1896
rect 6967 1856 7012 1884
rect 6549 1847 6607 1853
rect 7006 1844 7012 1856
rect 7064 1844 7070 1896
rect 3510 1776 3516 1828
rect 3568 1816 3574 1828
rect 4433 1819 4491 1825
rect 4433 1816 4445 1819
rect 3568 1788 4445 1816
rect 3568 1776 3574 1788
rect 4433 1785 4445 1788
rect 4479 1785 4491 1819
rect 4433 1779 4491 1785
rect 6365 1819 6423 1825
rect 6365 1785 6377 1819
rect 6411 1816 6423 1819
rect 6914 1816 6920 1828
rect 6411 1788 6920 1816
rect 6411 1785 6423 1788
rect 6365 1779 6423 1785
rect 6914 1776 6920 1788
rect 6972 1776 6978 1828
rect 7392 1816 7420 1915
rect 7576 1884 7604 1915
rect 7650 1912 7656 1964
rect 7708 1952 7714 1964
rect 7837 1955 7895 1961
rect 7837 1952 7849 1955
rect 7708 1924 7849 1952
rect 7708 1912 7714 1924
rect 7837 1921 7849 1924
rect 7883 1921 7895 1955
rect 7837 1915 7895 1921
rect 7926 1912 7932 1964
rect 7984 1952 7990 1964
rect 8220 1961 8248 1992
rect 8297 1989 8309 2023
rect 8343 2020 8355 2023
rect 8343 1992 8524 2020
rect 8343 1989 8355 1992
rect 8297 1983 8355 1989
rect 8496 1961 8524 1992
rect 8113 1955 8171 1961
rect 7984 1924 8029 1952
rect 7984 1912 7990 1924
rect 8113 1921 8125 1955
rect 8159 1921 8171 1955
rect 8113 1915 8171 1921
rect 8205 1955 8263 1961
rect 8205 1921 8217 1955
rect 8251 1921 8263 1955
rect 8389 1955 8447 1961
rect 8389 1952 8401 1955
rect 8205 1915 8263 1921
rect 8312 1924 8401 1952
rect 8018 1884 8024 1896
rect 7576 1856 8024 1884
rect 8018 1844 8024 1856
rect 8076 1884 8082 1896
rect 8128 1884 8156 1915
rect 8076 1856 8156 1884
rect 8076 1844 8082 1856
rect 7466 1816 7472 1828
rect 7379 1788 7472 1816
rect 7466 1776 7472 1788
rect 7524 1816 7530 1828
rect 8312 1816 8340 1924
rect 8389 1921 8401 1924
rect 8435 1921 8447 1955
rect 8389 1915 8447 1921
rect 8481 1955 8539 1961
rect 8481 1921 8493 1955
rect 8527 1921 8539 1955
rect 8481 1915 8539 1921
rect 8665 1955 8723 1961
rect 8665 1921 8677 1955
rect 8711 1952 8723 1955
rect 8754 1952 8760 1964
rect 8711 1924 8760 1952
rect 8711 1921 8723 1924
rect 8665 1915 8723 1921
rect 8754 1912 8760 1924
rect 8812 1912 8818 1964
rect 9214 1952 9220 1964
rect 9175 1924 9220 1952
rect 9214 1912 9220 1924
rect 9272 1912 9278 1964
rect 9324 1961 9352 2048
rect 9398 1980 9404 2032
rect 9456 2020 9462 2032
rect 9677 2023 9735 2029
rect 9677 2020 9689 2023
rect 9456 1992 9689 2020
rect 9456 1980 9462 1992
rect 9677 1989 9689 1992
rect 9723 2020 9735 2023
rect 10318 2020 10324 2032
rect 9723 1992 10324 2020
rect 9723 1989 9735 1992
rect 9677 1983 9735 1989
rect 10318 1980 10324 1992
rect 10376 2020 10382 2032
rect 10376 1992 11100 2020
rect 10376 1980 10382 1992
rect 9309 1955 9367 1961
rect 9309 1921 9321 1955
rect 9355 1921 9367 1955
rect 9309 1915 9367 1921
rect 9766 1912 9772 1964
rect 9824 1952 9830 1964
rect 10137 1955 10195 1961
rect 10137 1952 10149 1955
rect 9824 1924 10149 1952
rect 9824 1912 9830 1924
rect 10137 1921 10149 1924
rect 10183 1952 10195 1955
rect 10686 1952 10692 1964
rect 10183 1924 10692 1952
rect 10183 1921 10195 1924
rect 10137 1915 10195 1921
rect 10686 1912 10692 1924
rect 10744 1912 10750 1964
rect 11072 1961 11100 1992
rect 11330 1980 11336 2032
rect 11388 2020 11394 2032
rect 12986 2020 12992 2032
rect 11388 1992 12992 2020
rect 11388 1980 11394 1992
rect 12986 1980 12992 1992
rect 13044 2020 13050 2032
rect 13648 2020 13676 2060
rect 13814 2048 13820 2060
rect 13872 2048 13878 2100
rect 14734 2048 14740 2100
rect 14792 2088 14798 2100
rect 14921 2091 14979 2097
rect 14921 2088 14933 2091
rect 14792 2060 14933 2088
rect 14792 2048 14798 2060
rect 14921 2057 14933 2060
rect 14967 2088 14979 2091
rect 15102 2088 15108 2100
rect 14967 2060 15108 2088
rect 14967 2057 14979 2060
rect 14921 2051 14979 2057
rect 15102 2048 15108 2060
rect 15160 2088 15166 2100
rect 17494 2088 17500 2100
rect 15160 2060 17500 2088
rect 15160 2048 15166 2060
rect 17494 2048 17500 2060
rect 17552 2048 17558 2100
rect 18230 2088 18236 2100
rect 18191 2060 18236 2088
rect 18230 2048 18236 2060
rect 18288 2048 18294 2100
rect 15378 2020 15384 2032
rect 13044 1992 13216 2020
rect 13648 1992 15384 2020
rect 13044 1980 13050 1992
rect 10873 1955 10931 1961
rect 10873 1952 10885 1955
rect 10805 1924 10885 1952
rect 9490 1844 9496 1896
rect 9548 1884 9554 1896
rect 10805 1884 10833 1924
rect 10873 1921 10885 1924
rect 10919 1921 10931 1955
rect 10873 1915 10931 1921
rect 11057 1955 11115 1961
rect 11057 1921 11069 1955
rect 11103 1921 11115 1955
rect 11057 1915 11115 1921
rect 11146 1912 11152 1964
rect 11204 1952 11210 1964
rect 11422 1952 11428 1964
rect 11204 1924 11249 1952
rect 11383 1924 11428 1952
rect 11204 1912 11210 1924
rect 11422 1912 11428 1924
rect 11480 1912 11486 1964
rect 11606 1912 11612 1964
rect 11664 1952 11670 1964
rect 11701 1955 11759 1961
rect 11701 1952 11713 1955
rect 11664 1924 11713 1952
rect 11664 1912 11670 1924
rect 11701 1921 11713 1924
rect 11747 1921 11759 1955
rect 11701 1915 11759 1921
rect 11885 1955 11943 1961
rect 11885 1921 11897 1955
rect 11931 1952 11943 1955
rect 12894 1952 12900 1964
rect 11931 1924 12900 1952
rect 11931 1921 11943 1924
rect 11885 1915 11943 1921
rect 12894 1912 12900 1924
rect 12952 1912 12958 1964
rect 13078 1952 13084 1964
rect 13039 1924 13084 1952
rect 13078 1912 13084 1924
rect 13136 1912 13142 1964
rect 11330 1884 11336 1896
rect 9548 1856 10833 1884
rect 11243 1856 11336 1884
rect 9548 1844 9554 1856
rect 7524 1788 8340 1816
rect 7524 1776 7530 1788
rect 8478 1776 8484 1828
rect 8536 1816 8542 1828
rect 9306 1816 9312 1828
rect 8536 1788 9312 1816
rect 8536 1776 8542 1788
rect 9306 1776 9312 1788
rect 9364 1776 9370 1828
rect 9401 1819 9459 1825
rect 9401 1785 9413 1819
rect 9447 1816 9459 1819
rect 10134 1816 10140 1828
rect 9447 1788 10140 1816
rect 9447 1785 9459 1788
rect 9401 1779 9459 1785
rect 10134 1776 10140 1788
rect 10192 1776 10198 1828
rect 10805 1816 10833 1856
rect 11330 1844 11336 1856
rect 11388 1884 11394 1896
rect 13188 1884 13216 1992
rect 15378 1980 15384 1992
rect 15436 1980 15442 2032
rect 17098 2023 17156 2029
rect 17098 2020 17110 2023
rect 16224 1992 17110 2020
rect 14001 1955 14059 1961
rect 14001 1921 14013 1955
rect 14047 1921 14059 1955
rect 14001 1915 14059 1921
rect 14185 1955 14243 1961
rect 14185 1921 14197 1955
rect 14231 1952 14243 1955
rect 14366 1952 14372 1964
rect 14231 1924 14372 1952
rect 14231 1921 14243 1924
rect 14185 1915 14243 1921
rect 13357 1887 13415 1893
rect 13357 1884 13369 1887
rect 11388 1856 13124 1884
rect 13188 1856 13369 1884
rect 11388 1844 11394 1856
rect 13096 1816 13124 1856
rect 13357 1853 13369 1856
rect 13403 1884 13415 1887
rect 13906 1884 13912 1896
rect 13403 1856 13912 1884
rect 13403 1853 13415 1856
rect 13357 1847 13415 1853
rect 13906 1844 13912 1856
rect 13964 1844 13970 1896
rect 14016 1816 14044 1915
rect 14366 1912 14372 1924
rect 14424 1912 14430 1964
rect 14826 1952 14832 1964
rect 14787 1924 14832 1952
rect 14826 1912 14832 1924
rect 14884 1912 14890 1964
rect 14918 1912 14924 1964
rect 14976 1952 14982 1964
rect 16224 1961 16252 1992
rect 17098 1989 17110 1992
rect 17144 2020 17156 2023
rect 17402 2020 17408 2032
rect 17144 1992 17408 2020
rect 17144 1989 17156 1992
rect 17098 1983 17156 1989
rect 17402 1980 17408 1992
rect 17460 1980 17466 2032
rect 16209 1955 16267 1961
rect 16209 1952 16221 1955
rect 14976 1924 16221 1952
rect 14976 1912 14982 1924
rect 16209 1921 16221 1924
rect 16255 1921 16267 1955
rect 16209 1915 16267 1921
rect 16301 1955 16359 1961
rect 16301 1921 16313 1955
rect 16347 1952 16359 1955
rect 16482 1952 16488 1964
rect 16347 1924 16488 1952
rect 16347 1921 16359 1924
rect 16301 1915 16359 1921
rect 16482 1912 16488 1924
rect 16540 1912 16546 1964
rect 14277 1887 14335 1893
rect 14277 1853 14289 1887
rect 14323 1884 14335 1887
rect 14458 1884 14464 1896
rect 14323 1856 14464 1884
rect 14323 1853 14335 1856
rect 14277 1847 14335 1853
rect 14458 1844 14464 1856
rect 14516 1844 14522 1896
rect 14936 1884 14964 1912
rect 14844 1856 14964 1884
rect 15013 1887 15071 1893
rect 14844 1816 14872 1856
rect 15013 1853 15025 1887
rect 15059 1884 15071 1887
rect 15470 1884 15476 1896
rect 15059 1856 15476 1884
rect 15059 1853 15071 1856
rect 15013 1847 15071 1853
rect 10805 1788 13032 1816
rect 13096 1788 14044 1816
rect 14108 1788 14872 1816
rect 842 1748 848 1760
rect 803 1720 848 1748
rect 842 1708 848 1720
rect 900 1708 906 1760
rect 5350 1708 5356 1760
rect 5408 1748 5414 1760
rect 7006 1748 7012 1760
rect 5408 1720 7012 1748
rect 5408 1708 5414 1720
rect 7006 1708 7012 1720
rect 7064 1708 7070 1760
rect 7282 1748 7288 1760
rect 7243 1720 7288 1748
rect 7282 1708 7288 1720
rect 7340 1708 7346 1760
rect 7834 1748 7840 1760
rect 7795 1720 7840 1748
rect 7834 1708 7840 1720
rect 7892 1708 7898 1760
rect 7926 1708 7932 1760
rect 7984 1748 7990 1760
rect 8754 1748 8760 1760
rect 7984 1720 8760 1748
rect 7984 1708 7990 1720
rect 8754 1708 8760 1720
rect 8812 1708 8818 1760
rect 9858 1708 9864 1760
rect 9916 1748 9922 1760
rect 10413 1751 10471 1757
rect 10413 1748 10425 1751
rect 9916 1720 10425 1748
rect 9916 1708 9922 1720
rect 10413 1717 10425 1720
rect 10459 1717 10471 1751
rect 10413 1711 10471 1717
rect 11054 1708 11060 1760
rect 11112 1748 11118 1760
rect 11330 1748 11336 1760
rect 11112 1720 11336 1748
rect 11112 1708 11118 1720
rect 11330 1708 11336 1720
rect 11388 1708 11394 1760
rect 12713 1751 12771 1757
rect 12713 1717 12725 1751
rect 12759 1748 12771 1751
rect 12802 1748 12808 1760
rect 12759 1720 12808 1748
rect 12759 1717 12771 1720
rect 12713 1711 12771 1717
rect 12802 1708 12808 1720
rect 12860 1708 12866 1760
rect 13004 1748 13032 1788
rect 14108 1748 14136 1788
rect 13004 1720 14136 1748
rect 14182 1708 14188 1760
rect 14240 1748 14246 1760
rect 14461 1751 14519 1757
rect 14461 1748 14473 1751
rect 14240 1720 14473 1748
rect 14240 1708 14246 1720
rect 14461 1717 14473 1720
rect 14507 1717 14519 1751
rect 14461 1711 14519 1717
rect 14734 1708 14740 1760
rect 14792 1748 14798 1760
rect 15028 1748 15056 1847
rect 15470 1844 15476 1856
rect 15528 1884 15534 1896
rect 16025 1887 16083 1893
rect 16025 1884 16037 1887
rect 15528 1856 16037 1884
rect 15528 1844 15534 1856
rect 16025 1853 16037 1856
rect 16071 1853 16083 1887
rect 16025 1847 16083 1853
rect 16114 1844 16120 1896
rect 16172 1884 16178 1896
rect 16853 1887 16911 1893
rect 16853 1884 16865 1887
rect 16172 1856 16865 1884
rect 16172 1844 16178 1856
rect 16853 1853 16865 1856
rect 16899 1853 16911 1887
rect 16853 1847 16911 1853
rect 16666 1748 16672 1760
rect 14792 1720 15056 1748
rect 16627 1720 16672 1748
rect 14792 1708 14798 1720
rect 16666 1708 16672 1720
rect 16724 1708 16730 1760
rect 0 1658 18860 1680
rect 0 1606 3110 1658
rect 3162 1606 3174 1658
rect 3226 1606 3238 1658
rect 3290 1606 3302 1658
rect 3354 1606 3366 1658
rect 3418 1606 6210 1658
rect 6262 1606 6274 1658
rect 6326 1606 6338 1658
rect 6390 1606 6402 1658
rect 6454 1606 6466 1658
rect 6518 1606 9310 1658
rect 9362 1606 9374 1658
rect 9426 1606 9438 1658
rect 9490 1606 9502 1658
rect 9554 1606 9566 1658
rect 9618 1606 12410 1658
rect 12462 1606 12474 1658
rect 12526 1606 12538 1658
rect 12590 1606 12602 1658
rect 12654 1606 12666 1658
rect 12718 1606 15510 1658
rect 15562 1606 15574 1658
rect 15626 1606 15638 1658
rect 15690 1606 15702 1658
rect 15754 1606 15766 1658
rect 15818 1606 18860 1658
rect 0 1584 18860 1606
rect 2774 1504 2780 1556
rect 2832 1544 2838 1556
rect 3053 1547 3111 1553
rect 3053 1544 3065 1547
rect 2832 1516 3065 1544
rect 2832 1504 2838 1516
rect 3053 1513 3065 1516
rect 3099 1513 3111 1547
rect 5902 1544 5908 1556
rect 5863 1516 5908 1544
rect 3053 1507 3111 1513
rect 845 1343 903 1349
rect 845 1309 857 1343
rect 891 1340 903 1343
rect 1302 1340 1308 1352
rect 891 1312 1308 1340
rect 891 1309 903 1312
rect 845 1303 903 1309
rect 1302 1300 1308 1312
rect 1360 1300 1366 1352
rect 3068 1340 3096 1507
rect 5902 1504 5908 1516
rect 5960 1504 5966 1556
rect 6638 1544 6644 1556
rect 6012 1516 6644 1544
rect 5629 1479 5687 1485
rect 5629 1445 5641 1479
rect 5675 1476 5687 1479
rect 6012 1476 6040 1516
rect 6638 1504 6644 1516
rect 6696 1504 6702 1556
rect 6914 1504 6920 1556
rect 6972 1544 6978 1556
rect 9674 1544 9680 1556
rect 6972 1516 9680 1544
rect 6972 1504 6978 1516
rect 9674 1504 9680 1516
rect 9732 1504 9738 1556
rect 10042 1544 10048 1556
rect 10003 1516 10048 1544
rect 10042 1504 10048 1516
rect 10100 1504 10106 1556
rect 11054 1544 11060 1556
rect 10428 1516 11060 1544
rect 7190 1476 7196 1488
rect 5675 1448 6040 1476
rect 6564 1448 7196 1476
rect 5675 1445 5687 1448
rect 5629 1439 5687 1445
rect 5258 1368 5264 1420
rect 5316 1408 5322 1420
rect 5353 1411 5411 1417
rect 5353 1408 5365 1411
rect 5316 1380 5365 1408
rect 5316 1368 5322 1380
rect 5353 1377 5365 1380
rect 5399 1377 5411 1411
rect 5994 1408 6000 1420
rect 5353 1371 5411 1377
rect 5644 1380 6000 1408
rect 3145 1343 3203 1349
rect 3145 1340 3157 1343
rect 3068 1312 3157 1340
rect 3145 1309 3157 1312
rect 3191 1309 3203 1343
rect 3145 1303 3203 1309
rect 3602 1300 3608 1352
rect 3660 1340 3666 1352
rect 4783 1343 4841 1349
rect 4783 1340 4795 1343
rect 3660 1312 4795 1340
rect 3660 1300 3666 1312
rect 4783 1309 4795 1312
rect 4829 1309 4841 1343
rect 4783 1303 4841 1309
rect 5077 1343 5135 1349
rect 5077 1309 5089 1343
rect 5123 1340 5135 1343
rect 5534 1340 5540 1352
rect 5123 1312 5540 1340
rect 5123 1309 5135 1312
rect 5077 1303 5135 1309
rect 5534 1300 5540 1312
rect 5592 1340 5598 1352
rect 5644 1340 5672 1380
rect 5994 1368 6000 1380
rect 6052 1368 6058 1420
rect 6564 1408 6592 1448
rect 7190 1436 7196 1448
rect 7248 1436 7254 1488
rect 7300 1448 7972 1476
rect 6380 1380 6592 1408
rect 5592 1312 5672 1340
rect 5721 1343 5779 1349
rect 5592 1300 5598 1312
rect 5721 1309 5733 1343
rect 5767 1309 5779 1343
rect 5721 1303 5779 1309
rect 5905 1343 5963 1349
rect 5905 1309 5917 1343
rect 5951 1340 5963 1343
rect 6380 1340 6408 1380
rect 6638 1368 6644 1420
rect 6696 1408 6702 1420
rect 6733 1411 6791 1417
rect 6733 1408 6745 1411
rect 6696 1380 6745 1408
rect 6696 1368 6702 1380
rect 6733 1377 6745 1380
rect 6779 1408 6791 1411
rect 7300 1408 7328 1448
rect 6779 1380 7328 1408
rect 6779 1377 6791 1380
rect 6733 1371 6791 1377
rect 7374 1368 7380 1420
rect 7432 1408 7438 1420
rect 7653 1411 7711 1417
rect 7432 1380 7477 1408
rect 7432 1368 7438 1380
rect 7653 1377 7665 1411
rect 7699 1408 7711 1411
rect 7834 1408 7840 1420
rect 7699 1380 7840 1408
rect 7699 1377 7711 1380
rect 7653 1371 7711 1377
rect 7834 1368 7840 1380
rect 7892 1368 7898 1420
rect 7944 1408 7972 1448
rect 8110 1436 8116 1488
rect 8168 1476 8174 1488
rect 10428 1476 10456 1516
rect 11054 1504 11060 1516
rect 11112 1504 11118 1556
rect 11146 1504 11152 1556
rect 11204 1544 11210 1556
rect 14642 1544 14648 1556
rect 11204 1516 12434 1544
rect 11204 1504 11210 1516
rect 10778 1476 10784 1488
rect 8168 1448 10456 1476
rect 10520 1448 10784 1476
rect 8168 1436 8174 1448
rect 9125 1411 9183 1417
rect 9125 1408 9137 1411
rect 7944 1380 9137 1408
rect 9125 1377 9137 1380
rect 9171 1408 9183 1411
rect 9766 1408 9772 1420
rect 9171 1380 9772 1408
rect 9171 1377 9183 1380
rect 9125 1371 9183 1377
rect 9766 1368 9772 1380
rect 9824 1368 9830 1420
rect 10520 1408 10548 1448
rect 10778 1436 10784 1448
rect 10836 1476 10842 1488
rect 11606 1476 11612 1488
rect 10836 1448 11612 1476
rect 10836 1436 10842 1448
rect 11606 1436 11612 1448
rect 11664 1476 11670 1488
rect 11790 1476 11796 1488
rect 11664 1448 11796 1476
rect 11664 1436 11670 1448
rect 11790 1436 11796 1448
rect 11848 1436 11854 1488
rect 9968 1380 10548 1408
rect 5951 1312 6408 1340
rect 6457 1343 6515 1349
rect 5951 1309 5963 1312
rect 5905 1303 5963 1309
rect 6457 1309 6469 1343
rect 6503 1340 6515 1343
rect 6546 1340 6552 1352
rect 6503 1312 6552 1340
rect 6503 1309 6515 1312
rect 6457 1303 6515 1309
rect 1578 1272 1584 1284
rect 1539 1244 1584 1272
rect 1578 1232 1584 1244
rect 1636 1232 1642 1284
rect 3418 1272 3424 1284
rect 382 1164 388 1216
rect 440 1204 446 1216
rect 569 1207 627 1213
rect 569 1204 581 1207
rect 440 1176 581 1204
rect 440 1164 446 1176
rect 569 1173 581 1176
rect 615 1173 627 1207
rect 569 1167 627 1173
rect 2590 1164 2596 1216
rect 2648 1204 2654 1216
rect 2792 1204 2820 1258
rect 3379 1244 3424 1272
rect 3418 1232 3424 1244
rect 3476 1232 3482 1284
rect 3970 1232 3976 1284
rect 4028 1272 4034 1284
rect 5261 1275 5319 1281
rect 5261 1272 5273 1275
rect 4028 1244 5273 1272
rect 4028 1232 4034 1244
rect 5261 1241 5273 1244
rect 5307 1272 5319 1275
rect 5629 1275 5687 1281
rect 5629 1272 5641 1275
rect 5307 1244 5641 1272
rect 5307 1241 5319 1244
rect 5261 1235 5319 1241
rect 5629 1241 5641 1244
rect 5675 1241 5687 1275
rect 5736 1272 5764 1303
rect 6546 1300 6552 1312
rect 6604 1300 6610 1352
rect 7098 1340 7104 1352
rect 6748 1312 7104 1340
rect 6362 1272 6368 1284
rect 5736 1244 6368 1272
rect 5629 1235 5687 1241
rect 6362 1232 6368 1244
rect 6420 1232 6426 1284
rect 3789 1207 3847 1213
rect 3789 1204 3801 1207
rect 2648 1176 3801 1204
rect 2648 1164 2654 1176
rect 3789 1173 3801 1176
rect 3835 1204 3847 1207
rect 3878 1204 3884 1216
rect 3835 1176 3884 1204
rect 3835 1173 3847 1176
rect 3789 1167 3847 1173
rect 3878 1164 3884 1176
rect 3936 1164 3942 1216
rect 6086 1204 6092 1216
rect 6047 1176 6092 1204
rect 6086 1164 6092 1176
rect 6144 1164 6150 1216
rect 6549 1207 6607 1213
rect 6549 1173 6561 1207
rect 6595 1204 6607 1207
rect 6748 1204 6776 1312
rect 7098 1300 7104 1312
rect 7156 1300 7162 1352
rect 7285 1343 7343 1349
rect 7285 1309 7297 1343
rect 7331 1340 7343 1343
rect 7466 1340 7472 1352
rect 7331 1312 7472 1340
rect 7331 1309 7343 1312
rect 7285 1303 7343 1309
rect 7466 1300 7472 1312
rect 7524 1300 7530 1352
rect 8021 1343 8079 1349
rect 8021 1309 8033 1343
rect 8067 1309 8079 1343
rect 8021 1303 8079 1309
rect 7190 1232 7196 1284
rect 7248 1272 7254 1284
rect 7374 1272 7380 1284
rect 7248 1244 7380 1272
rect 7248 1232 7254 1244
rect 7374 1232 7380 1244
rect 7432 1232 7438 1284
rect 8036 1272 8064 1303
rect 8110 1300 8116 1352
rect 8168 1340 8174 1352
rect 8297 1343 8355 1349
rect 8168 1312 8213 1340
rect 8168 1300 8174 1312
rect 8297 1309 8309 1343
rect 8343 1340 8355 1343
rect 8846 1340 8852 1352
rect 8343 1312 8852 1340
rect 8343 1309 8355 1312
rect 8297 1303 8355 1309
rect 8846 1300 8852 1312
rect 8904 1300 8910 1352
rect 9858 1340 9864 1352
rect 9819 1312 9864 1340
rect 9858 1300 9864 1312
rect 9916 1300 9922 1352
rect 8036 1244 8524 1272
rect 6914 1204 6920 1216
rect 6595 1176 6776 1204
rect 6875 1176 6920 1204
rect 6595 1173 6607 1176
rect 6549 1167 6607 1173
rect 6914 1164 6920 1176
rect 6972 1164 6978 1216
rect 7006 1164 7012 1216
rect 7064 1204 7070 1216
rect 8202 1204 8208 1216
rect 7064 1176 8208 1204
rect 7064 1164 7070 1176
rect 8202 1164 8208 1176
rect 8260 1164 8266 1216
rect 8496 1213 8524 1244
rect 9674 1232 9680 1284
rect 9732 1272 9738 1284
rect 9968 1272 9996 1380
rect 10134 1340 10140 1352
rect 10095 1312 10140 1340
rect 10134 1300 10140 1312
rect 10192 1300 10198 1352
rect 10318 1340 10324 1352
rect 10279 1312 10324 1340
rect 10318 1300 10324 1312
rect 10376 1300 10382 1352
rect 10520 1349 10548 1380
rect 11149 1411 11207 1417
rect 11149 1377 11161 1411
rect 11195 1408 11207 1411
rect 11330 1408 11336 1420
rect 11195 1380 11336 1408
rect 11195 1377 11207 1380
rect 11149 1371 11207 1377
rect 11330 1368 11336 1380
rect 11388 1368 11394 1420
rect 12406 1408 12434 1516
rect 12728 1516 14648 1544
rect 12728 1417 12756 1516
rect 14642 1504 14648 1516
rect 14700 1504 14706 1556
rect 14737 1547 14795 1553
rect 14737 1513 14749 1547
rect 14783 1544 14795 1547
rect 14826 1544 14832 1556
rect 14783 1516 14832 1544
rect 14783 1513 14795 1516
rect 14737 1507 14795 1513
rect 14826 1504 14832 1516
rect 14884 1504 14890 1556
rect 14182 1436 14188 1488
rect 14240 1436 14246 1488
rect 14274 1436 14280 1488
rect 14332 1476 14338 1488
rect 14332 1448 15424 1476
rect 14332 1436 14338 1448
rect 12713 1411 12771 1417
rect 12713 1408 12725 1411
rect 12406 1380 12725 1408
rect 12713 1377 12725 1380
rect 12759 1377 12771 1411
rect 12713 1371 12771 1377
rect 10505 1343 10563 1349
rect 10505 1309 10517 1343
rect 10551 1309 10563 1343
rect 11241 1343 11299 1349
rect 11241 1340 11253 1343
rect 10505 1303 10563 1309
rect 10888 1312 11253 1340
rect 9732 1244 9996 1272
rect 9732 1232 9738 1244
rect 8481 1207 8539 1213
rect 8481 1173 8493 1207
rect 8527 1173 8539 1207
rect 8481 1167 8539 1173
rect 8570 1164 8576 1216
rect 8628 1204 8634 1216
rect 8849 1207 8907 1213
rect 8849 1204 8861 1207
rect 8628 1176 8861 1204
rect 8628 1164 8634 1176
rect 8849 1173 8861 1176
rect 8895 1173 8907 1207
rect 8849 1167 8907 1173
rect 8941 1207 8999 1213
rect 8941 1173 8953 1207
rect 8987 1204 8999 1207
rect 9401 1207 9459 1213
rect 9401 1204 9413 1207
rect 8987 1176 9413 1204
rect 8987 1173 8999 1176
rect 8941 1167 8999 1173
rect 9401 1173 9413 1176
rect 9447 1173 9459 1207
rect 10336 1204 10364 1300
rect 10413 1275 10471 1281
rect 10413 1241 10425 1275
rect 10459 1272 10471 1275
rect 10888 1272 10916 1312
rect 11241 1309 11253 1312
rect 11287 1309 11299 1343
rect 11241 1303 11299 1309
rect 11425 1343 11483 1349
rect 11425 1309 11437 1343
rect 11471 1340 11483 1343
rect 11471 1312 12204 1340
rect 11471 1309 11483 1312
rect 11425 1303 11483 1309
rect 10459 1244 10916 1272
rect 10965 1275 11023 1281
rect 10459 1241 10471 1244
rect 10413 1235 10471 1241
rect 10965 1241 10977 1275
rect 11011 1241 11023 1275
rect 11256 1272 11284 1303
rect 12066 1272 12072 1284
rect 11256 1244 12072 1272
rect 10965 1235 11023 1241
rect 10980 1204 11008 1235
rect 12066 1232 12072 1244
rect 12124 1232 12130 1284
rect 11238 1204 11244 1216
rect 10336 1176 11008 1204
rect 11199 1176 11244 1204
rect 9401 1167 9459 1173
rect 11238 1164 11244 1176
rect 11296 1164 11302 1216
rect 12176 1213 12204 1312
rect 12250 1300 12256 1352
rect 12308 1340 12314 1352
rect 13265 1343 13323 1349
rect 13265 1340 13277 1343
rect 12308 1312 13277 1340
rect 12308 1300 12314 1312
rect 13265 1309 13277 1312
rect 13311 1309 13323 1343
rect 13265 1303 13323 1309
rect 13449 1343 13507 1349
rect 13449 1309 13461 1343
rect 13495 1309 13507 1343
rect 13449 1303 13507 1309
rect 12529 1275 12587 1281
rect 12529 1241 12541 1275
rect 12575 1272 12587 1275
rect 12802 1272 12808 1284
rect 12575 1244 12808 1272
rect 12575 1241 12587 1244
rect 12529 1235 12587 1241
rect 12802 1232 12808 1244
rect 12860 1232 12866 1284
rect 13170 1232 13176 1284
rect 13228 1272 13234 1284
rect 13464 1272 13492 1303
rect 13538 1300 13544 1352
rect 13596 1340 13602 1352
rect 14001 1343 14059 1349
rect 14001 1340 14013 1343
rect 13596 1312 14013 1340
rect 13596 1300 13602 1312
rect 14001 1309 14013 1312
rect 14047 1340 14059 1343
rect 14090 1340 14096 1352
rect 14047 1312 14096 1340
rect 14047 1309 14059 1312
rect 14001 1303 14059 1309
rect 14090 1300 14096 1312
rect 14148 1300 14154 1352
rect 14200 1349 14228 1436
rect 15102 1368 15108 1420
rect 15160 1408 15166 1420
rect 15396 1417 15424 1448
rect 15197 1411 15255 1417
rect 15197 1408 15209 1411
rect 15160 1380 15209 1408
rect 15160 1368 15166 1380
rect 15197 1377 15209 1380
rect 15243 1377 15255 1411
rect 15197 1371 15255 1377
rect 15381 1411 15439 1417
rect 15381 1377 15393 1411
rect 15427 1408 15439 1411
rect 15654 1408 15660 1420
rect 15427 1380 15660 1408
rect 15427 1377 15439 1380
rect 15381 1371 15439 1377
rect 15654 1368 15660 1380
rect 15712 1368 15718 1420
rect 14185 1343 14243 1349
rect 14185 1309 14197 1343
rect 14231 1309 14243 1343
rect 14185 1303 14243 1309
rect 14277 1343 14335 1349
rect 14277 1309 14289 1343
rect 14323 1309 14335 1343
rect 16114 1340 16120 1352
rect 16027 1312 16120 1340
rect 14277 1303 14335 1309
rect 13228 1244 13492 1272
rect 13228 1232 13234 1244
rect 13722 1232 13728 1284
rect 13780 1272 13786 1284
rect 14292 1272 14320 1303
rect 16114 1300 16120 1312
rect 16172 1300 16178 1352
rect 16132 1272 16160 1300
rect 16390 1272 16396 1284
rect 13780 1244 16160 1272
rect 16351 1244 16396 1272
rect 13780 1232 13786 1244
rect 16390 1232 16396 1244
rect 16448 1232 16454 1284
rect 12161 1207 12219 1213
rect 12161 1173 12173 1207
rect 12207 1173 12219 1207
rect 12618 1204 12624 1216
rect 12579 1176 12624 1204
rect 12161 1167 12219 1173
rect 12618 1164 12624 1176
rect 12676 1164 12682 1216
rect 12894 1164 12900 1216
rect 12952 1204 12958 1216
rect 13265 1207 13323 1213
rect 13265 1204 13277 1207
rect 12952 1176 13277 1204
rect 12952 1164 12958 1176
rect 13265 1173 13277 1176
rect 13311 1173 13323 1207
rect 13265 1167 13323 1173
rect 13814 1164 13820 1216
rect 13872 1204 13878 1216
rect 14001 1207 14059 1213
rect 14001 1204 14013 1207
rect 13872 1176 14013 1204
rect 13872 1164 13878 1176
rect 14001 1173 14013 1176
rect 14047 1173 14059 1207
rect 14001 1167 14059 1173
rect 14458 1164 14464 1216
rect 14516 1204 14522 1216
rect 14553 1207 14611 1213
rect 14553 1204 14565 1207
rect 14516 1176 14565 1204
rect 14516 1164 14522 1176
rect 14553 1173 14565 1176
rect 14599 1173 14611 1207
rect 14553 1167 14611 1173
rect 15010 1164 15016 1216
rect 15068 1204 15074 1216
rect 15105 1207 15163 1213
rect 15105 1204 15117 1207
rect 15068 1176 15117 1204
rect 15068 1164 15074 1176
rect 15105 1173 15117 1176
rect 15151 1173 15163 1207
rect 15105 1167 15163 1173
rect 15838 1164 15844 1216
rect 15896 1204 15902 1216
rect 16025 1207 16083 1213
rect 16025 1204 16037 1207
rect 15896 1176 16037 1204
rect 15896 1164 15902 1176
rect 16025 1173 16037 1176
rect 16071 1204 16083 1207
rect 16868 1204 16896 1258
rect 17862 1204 17868 1216
rect 16071 1176 16896 1204
rect 17823 1176 17868 1204
rect 16071 1173 16083 1176
rect 16025 1167 16083 1173
rect 17862 1164 17868 1176
rect 17920 1164 17926 1216
rect 0 1114 18860 1136
rect 0 1062 4660 1114
rect 4712 1062 4724 1114
rect 4776 1062 4788 1114
rect 4840 1062 4852 1114
rect 4904 1062 4916 1114
rect 4968 1062 7760 1114
rect 7812 1062 7824 1114
rect 7876 1062 7888 1114
rect 7940 1062 7952 1114
rect 8004 1062 8016 1114
rect 8068 1062 10860 1114
rect 10912 1062 10924 1114
rect 10976 1062 10988 1114
rect 11040 1062 11052 1114
rect 11104 1062 11116 1114
rect 11168 1062 13960 1114
rect 14012 1062 14024 1114
rect 14076 1062 14088 1114
rect 14140 1062 14152 1114
rect 14204 1062 14216 1114
rect 14268 1062 17060 1114
rect 17112 1062 17124 1114
rect 17176 1062 17188 1114
rect 17240 1062 17252 1114
rect 17304 1062 17316 1114
rect 17368 1062 18860 1114
rect 0 1040 18860 1062
rect 2774 960 2780 1012
rect 2832 1000 2838 1012
rect 2869 1003 2927 1009
rect 2869 1000 2881 1003
rect 2832 972 2881 1000
rect 2832 960 2838 972
rect 2869 969 2881 972
rect 2915 969 2927 1003
rect 2869 963 2927 969
rect 2961 1003 3019 1009
rect 2961 969 2973 1003
rect 3007 1000 3019 1003
rect 3329 1003 3387 1009
rect 3329 1000 3341 1003
rect 3007 972 3341 1000
rect 3007 969 3019 972
rect 2961 963 3019 969
rect 3329 969 3341 972
rect 3375 969 3387 1003
rect 3329 963 3387 969
rect 3418 960 3424 1012
rect 3476 1000 3482 1012
rect 3697 1003 3755 1009
rect 3697 1000 3709 1003
rect 3476 972 3709 1000
rect 3476 960 3482 972
rect 3697 969 3709 972
rect 3743 969 3755 1003
rect 3697 963 3755 969
rect 5810 960 5816 1012
rect 5868 1000 5874 1012
rect 6825 1003 6883 1009
rect 6825 1000 6837 1003
rect 5868 972 6837 1000
rect 5868 960 5874 972
rect 6825 969 6837 972
rect 6871 969 6883 1003
rect 9122 1000 9128 1012
rect 6825 963 6883 969
rect 6932 972 9128 1000
rect 2222 941 2228 944
rect 2179 935 2228 941
rect 382 864 388 876
rect 343 836 388 864
rect 382 824 388 836
rect 440 824 446 876
rect 753 867 811 873
rect 753 833 765 867
rect 799 864 811 867
rect 842 864 848 876
rect 799 836 848 864
rect 799 833 811 836
rect 753 827 811 833
rect 842 824 848 836
rect 900 824 906 876
rect 1780 864 1808 918
rect 2179 901 2191 935
rect 2225 901 2228 935
rect 2179 895 2228 901
rect 2222 892 2228 895
rect 2280 892 2286 944
rect 6932 932 6960 972
rect 8404 944 8432 972
rect 9122 960 9128 972
rect 9180 1000 9186 1012
rect 9306 1000 9312 1012
rect 9180 972 9312 1000
rect 9180 960 9186 972
rect 9306 960 9312 972
rect 9364 960 9370 1012
rect 13722 1000 13728 1012
rect 9876 972 13728 1000
rect 6302 918 6960 932
rect 6288 904 6960 918
rect 2590 864 2596 876
rect 1780 836 2596 864
rect 2590 824 2596 836
rect 2648 824 2654 876
rect 4893 867 4951 873
rect 4893 833 4905 867
rect 4939 864 4951 867
rect 5166 864 5172 876
rect 4939 836 5172 864
rect 4939 833 4951 836
rect 4893 827 4951 833
rect 5166 824 5172 836
rect 5224 824 5230 876
rect 3145 799 3203 805
rect 3145 765 3157 799
rect 3191 796 3203 799
rect 3602 796 3608 808
rect 3191 768 3608 796
rect 3191 765 3203 768
rect 3145 759 3203 765
rect 3602 756 3608 768
rect 3660 756 3666 808
rect 3786 796 3792 808
rect 3747 768 3792 796
rect 3786 756 3792 768
rect 3844 756 3850 808
rect 3970 796 3976 808
rect 3931 768 3976 796
rect 3970 756 3976 768
rect 4028 756 4034 808
rect 5258 796 5264 808
rect 5219 768 5264 796
rect 5258 756 5264 768
rect 5316 756 5322 808
rect 1302 620 1308 672
rect 1360 660 1366 672
rect 2501 663 2559 669
rect 2501 660 2513 663
rect 1360 632 2513 660
rect 1360 620 1366 632
rect 2501 629 2513 632
rect 2547 629 2559 663
rect 2501 623 2559 629
rect 3878 620 3884 672
rect 3936 660 3942 672
rect 4709 663 4767 669
rect 4709 660 4721 663
rect 3936 632 4721 660
rect 3936 620 3942 632
rect 4709 629 4721 632
rect 4755 660 4767 663
rect 6288 660 6316 904
rect 8386 892 8392 944
rect 8444 892 8450 944
rect 8846 932 8852 944
rect 8807 904 8852 932
rect 8846 892 8852 904
rect 8904 892 8910 944
rect 9876 932 9904 972
rect 13722 960 13728 972
rect 13780 960 13786 1012
rect 13909 1003 13967 1009
rect 13909 969 13921 1003
rect 13955 1000 13967 1003
rect 13955 972 14320 1000
rect 13955 969 13967 972
rect 13909 963 13967 969
rect 12158 932 12164 944
rect 9140 904 9904 932
rect 7006 864 7012 876
rect 6967 836 7012 864
rect 7006 824 7012 836
rect 7064 824 7070 876
rect 9140 873 9168 904
rect 9876 873 9904 904
rect 9968 904 10626 932
rect 12119 904 12164 932
rect 9125 867 9183 873
rect 9125 833 9137 867
rect 9171 833 9183 867
rect 9125 827 9183 833
rect 9217 867 9275 873
rect 9217 833 9229 867
rect 9263 833 9275 867
rect 9217 827 9275 833
rect 9861 867 9919 873
rect 9861 833 9873 867
rect 9907 833 9919 867
rect 9861 827 9919 833
rect 7374 796 7380 808
rect 7287 768 7380 796
rect 7374 756 7380 768
rect 7432 796 7438 808
rect 8754 796 8760 808
rect 7432 768 8760 796
rect 7432 756 7438 768
rect 8754 756 8760 768
rect 8812 796 8818 808
rect 9232 796 9260 827
rect 8812 768 9260 796
rect 8812 756 8818 768
rect 9306 756 9312 808
rect 9364 796 9370 808
rect 9769 799 9827 805
rect 9769 796 9781 799
rect 9364 768 9781 796
rect 9364 756 9370 768
rect 9769 765 9781 768
rect 9815 796 9827 799
rect 9968 796 9996 904
rect 12158 892 12164 904
rect 12216 892 12222 944
rect 12894 932 12900 944
rect 12855 904 12900 932
rect 12894 892 12900 904
rect 12952 892 12958 944
rect 13004 904 13584 932
rect 12342 874 12348 876
rect 12268 873 12348 874
rect 12069 867 12127 873
rect 12069 864 12081 867
rect 11624 836 12081 864
rect 9815 768 9996 796
rect 10137 799 10195 805
rect 9815 765 9827 768
rect 9769 759 9827 765
rect 10137 765 10149 799
rect 10183 796 10195 799
rect 10594 796 10600 808
rect 10183 768 10600 796
rect 10183 765 10195 768
rect 10137 759 10195 765
rect 10594 756 10600 768
rect 10652 756 10658 808
rect 6362 688 6368 740
rect 6420 728 6426 740
rect 6687 731 6745 737
rect 6687 728 6699 731
rect 6420 700 6699 728
rect 6420 688 6426 700
rect 6687 697 6699 700
rect 6733 728 6745 731
rect 7466 728 7472 740
rect 6733 700 7472 728
rect 6733 697 6745 700
rect 6687 691 6745 697
rect 7466 688 7472 700
rect 7524 688 7530 740
rect 11624 672 11652 836
rect 12069 833 12081 836
rect 12115 833 12127 867
rect 12069 827 12127 833
rect 12253 867 12348 873
rect 12253 833 12265 867
rect 12299 846 12348 867
rect 12299 833 12311 846
rect 12253 827 12311 833
rect 12084 796 12112 827
rect 12342 824 12348 846
rect 12400 824 12406 876
rect 12437 870 12495 873
rect 12437 867 12664 870
rect 12437 833 12449 867
rect 12483 842 12664 867
rect 12802 864 12808 876
rect 12483 833 12495 842
rect 12437 827 12495 833
rect 12636 796 12664 842
rect 12715 836 12808 864
rect 12802 824 12808 836
rect 12860 864 12866 876
rect 13004 864 13032 904
rect 13170 864 13176 876
rect 12860 836 13032 864
rect 13131 836 13176 864
rect 12860 824 12866 836
rect 13170 824 13176 836
rect 13228 824 13234 876
rect 13556 873 13584 904
rect 13814 892 13820 944
rect 13872 932 13878 944
rect 14292 932 14320 972
rect 14366 960 14372 1012
rect 14424 1000 14430 1012
rect 16390 1000 16396 1012
rect 14424 972 15976 1000
rect 16351 972 16396 1000
rect 14424 960 14430 972
rect 13872 904 14228 932
rect 14292 904 14596 932
rect 13872 892 13878 904
rect 14200 873 14228 904
rect 13265 867 13323 873
rect 13265 833 13277 867
rect 13311 833 13323 867
rect 13265 827 13323 833
rect 13357 867 13415 873
rect 13357 833 13369 867
rect 13403 833 13415 867
rect 13357 827 13415 833
rect 13541 867 13599 873
rect 13541 833 13553 867
rect 13587 864 13599 867
rect 13633 867 13691 873
rect 13633 864 13645 867
rect 13587 836 13645 864
rect 13587 833 13599 836
rect 13541 827 13599 833
rect 13633 833 13645 836
rect 13679 833 13691 867
rect 13633 827 13691 833
rect 14001 867 14059 873
rect 14001 833 14013 867
rect 14047 833 14059 867
rect 14001 827 14059 833
rect 14185 867 14243 873
rect 14185 833 14197 867
rect 14231 833 14243 867
rect 14458 864 14464 876
rect 14419 836 14464 864
rect 14185 827 14243 833
rect 12084 768 12664 796
rect 11790 688 11796 740
rect 11848 728 11854 740
rect 13280 728 13308 827
rect 11848 700 13308 728
rect 11848 688 11854 700
rect 4755 632 6316 660
rect 4755 629 4767 632
rect 4709 623 4767 629
rect 8846 620 8852 672
rect 8904 660 8910 672
rect 9217 663 9275 669
rect 9217 660 9229 663
rect 8904 632 9229 660
rect 8904 620 8910 632
rect 9217 629 9229 632
rect 9263 629 9275 663
rect 11606 660 11612 672
rect 11567 632 11612 660
rect 9217 623 9275 629
rect 11606 620 11612 632
rect 11664 620 11670 672
rect 11698 620 11704 672
rect 11756 660 11762 672
rect 13372 660 13400 827
rect 14016 796 14044 827
rect 14458 824 14464 836
rect 14516 824 14522 876
rect 14568 864 14596 904
rect 15838 892 15844 944
rect 15896 892 15902 944
rect 14568 836 14964 864
rect 13464 768 14044 796
rect 14093 799 14151 805
rect 13464 737 13492 768
rect 14093 765 14105 799
rect 14139 796 14151 799
rect 14829 799 14887 805
rect 14829 796 14841 799
rect 14139 768 14841 796
rect 14139 765 14151 768
rect 14093 759 14151 765
rect 14829 765 14841 768
rect 14875 765 14887 799
rect 14936 796 14964 836
rect 15194 796 15200 808
rect 14936 768 15200 796
rect 14829 759 14887 765
rect 15194 756 15200 768
rect 15252 796 15258 808
rect 15856 796 15884 892
rect 15948 864 15976 972
rect 16390 960 16396 972
rect 16448 960 16454 1012
rect 16482 960 16488 1012
rect 16540 1000 16546 1012
rect 16853 1003 16911 1009
rect 16853 1000 16865 1003
rect 16540 972 16865 1000
rect 16540 960 16546 972
rect 16853 969 16865 972
rect 16899 969 16911 1003
rect 16853 963 16911 969
rect 17313 1003 17371 1009
rect 17313 969 17325 1003
rect 17359 1000 17371 1003
rect 17402 1000 17408 1012
rect 17359 972 17408 1000
rect 17359 969 17371 972
rect 17313 963 17371 969
rect 17402 960 17408 972
rect 17460 960 17466 1012
rect 16574 864 16580 876
rect 15948 836 16580 864
rect 16574 824 16580 836
rect 16632 824 16638 876
rect 16669 867 16727 873
rect 16669 833 16681 867
rect 16715 864 16727 867
rect 17218 864 17224 876
rect 16715 836 17224 864
rect 16715 833 16727 836
rect 16669 827 16727 833
rect 17218 824 17224 836
rect 17276 824 17282 876
rect 18233 867 18291 873
rect 18233 833 18245 867
rect 18279 864 18291 867
rect 18322 864 18328 876
rect 18279 836 18328 864
rect 18279 833 18291 836
rect 18233 827 18291 833
rect 18322 824 18328 836
rect 18380 824 18386 876
rect 15252 768 15884 796
rect 16393 799 16451 805
rect 15252 756 15258 768
rect 16393 765 16405 799
rect 16439 796 16451 799
rect 16942 796 16948 808
rect 16439 768 16948 796
rect 16439 765 16451 768
rect 16393 759 16451 765
rect 16942 756 16948 768
rect 17000 756 17006 808
rect 17405 799 17463 805
rect 17405 765 17417 799
rect 17451 765 17463 799
rect 18506 796 18512 808
rect 18467 768 18512 796
rect 17405 759 17463 765
rect 13449 731 13507 737
rect 13449 697 13461 731
rect 13495 697 13507 731
rect 13449 691 13507 697
rect 15654 688 15660 740
rect 15712 728 15718 740
rect 17420 728 17448 759
rect 18506 756 18512 768
rect 18564 756 18570 808
rect 15712 700 17448 728
rect 15712 688 15718 700
rect 11756 632 13400 660
rect 13633 663 13691 669
rect 11756 620 11762 632
rect 13633 629 13645 663
rect 13679 660 13691 663
rect 14734 660 14740 672
rect 13679 632 14740 660
rect 13679 629 13691 632
rect 13633 623 13691 629
rect 14734 620 14740 632
rect 14792 660 14798 672
rect 16255 663 16313 669
rect 16255 660 16267 663
rect 14792 632 16267 660
rect 14792 620 14798 632
rect 16255 629 16267 632
rect 16301 629 16313 663
rect 16255 623 16313 629
rect 0 570 18860 592
rect 0 518 3110 570
rect 3162 518 3174 570
rect 3226 518 3238 570
rect 3290 518 3302 570
rect 3354 518 3366 570
rect 3418 518 6210 570
rect 6262 518 6274 570
rect 6326 518 6338 570
rect 6390 518 6402 570
rect 6454 518 6466 570
rect 6518 518 9310 570
rect 9362 518 9374 570
rect 9426 518 9438 570
rect 9490 518 9502 570
rect 9554 518 9566 570
rect 9618 518 12410 570
rect 12462 518 12474 570
rect 12526 518 12538 570
rect 12590 518 12602 570
rect 12654 518 12666 570
rect 12718 518 15510 570
rect 15562 518 15574 570
rect 15626 518 15638 570
rect 15690 518 15702 570
rect 15754 518 15766 570
rect 15818 518 18860 570
rect 0 496 18860 518
rect 1489 459 1547 465
rect 1489 425 1501 459
rect 1535 456 1547 459
rect 1578 456 1584 468
rect 1535 428 1584 456
rect 1535 425 1547 428
rect 1489 419 1547 425
rect 1578 416 1584 428
rect 1636 416 1642 468
rect 2590 456 2596 468
rect 2551 428 2596 456
rect 2590 416 2596 428
rect 2648 416 2654 468
rect 3421 459 3479 465
rect 3421 425 3433 459
rect 3467 456 3479 459
rect 3786 456 3792 468
rect 3467 428 3792 456
rect 3467 425 3479 428
rect 3421 419 3479 425
rect 3786 416 3792 428
rect 3844 416 3850 468
rect 4893 459 4951 465
rect 4893 425 4905 459
rect 4939 456 4951 459
rect 5258 456 5264 468
rect 4939 428 5264 456
rect 4939 425 4951 428
rect 4893 419 4951 425
rect 5258 416 5264 428
rect 5316 416 5322 468
rect 6365 459 6423 465
rect 6365 425 6377 459
rect 6411 456 6423 459
rect 6546 456 6552 468
rect 6411 428 6552 456
rect 6411 425 6423 428
rect 6365 419 6423 425
rect 6546 416 6552 428
rect 6604 416 6610 468
rect 7098 456 7104 468
rect 6840 428 7104 456
rect 5534 388 5540 400
rect 5092 360 5540 388
rect 3237 323 3295 329
rect 3237 289 3249 323
rect 3283 320 3295 323
rect 3510 320 3516 332
rect 3283 292 3516 320
rect 3283 289 3295 292
rect 3237 283 3295 289
rect 3510 280 3516 292
rect 3568 280 3574 332
rect 5092 329 5120 360
rect 5534 348 5540 360
rect 5592 348 5598 400
rect 5077 323 5135 329
rect 5077 289 5089 323
rect 5123 289 5135 323
rect 5077 283 5135 289
rect 5169 323 5227 329
rect 5169 289 5181 323
rect 5215 320 5227 323
rect 6086 320 6092 332
rect 5215 292 6092 320
rect 5215 289 5227 292
rect 5169 283 5227 289
rect 6086 280 6092 292
rect 6144 280 6150 332
rect 6840 329 6868 428
rect 7098 416 7104 428
rect 7156 456 7162 468
rect 7285 459 7343 465
rect 7285 456 7297 459
rect 7156 428 7297 456
rect 7156 416 7162 428
rect 7285 425 7297 428
rect 7331 425 7343 459
rect 7285 419 7343 425
rect 7561 459 7619 465
rect 7561 425 7573 459
rect 7607 456 7619 459
rect 8386 456 8392 468
rect 7607 428 8392 456
rect 7607 425 7619 428
rect 7561 419 7619 425
rect 8386 416 8392 428
rect 8444 416 8450 468
rect 8481 459 8539 465
rect 8481 425 8493 459
rect 8527 456 8539 459
rect 8570 456 8576 468
rect 8527 428 8576 456
rect 8527 425 8539 428
rect 8481 419 8539 425
rect 8570 416 8576 428
rect 8628 416 8634 468
rect 10594 456 10600 468
rect 10555 428 10600 456
rect 10594 416 10600 428
rect 10652 416 10658 468
rect 12713 459 12771 465
rect 12713 425 12725 459
rect 12759 456 12771 459
rect 13078 456 13084 468
rect 12759 428 13084 456
rect 12759 425 12771 428
rect 12713 419 12771 425
rect 13078 416 13084 428
rect 13136 416 13142 468
rect 15010 456 15016 468
rect 14971 428 15016 456
rect 15010 416 15016 428
rect 15068 416 15074 468
rect 16942 456 16948 468
rect 16903 428 16948 456
rect 16942 416 16948 428
rect 17000 416 17006 468
rect 17218 456 17224 468
rect 17179 428 17224 456
rect 17218 416 17224 428
rect 17276 416 17282 468
rect 18506 456 18512 468
rect 18467 428 18512 456
rect 18506 416 18512 428
rect 18564 416 18570 468
rect 12989 391 13047 397
rect 12989 388 13001 391
rect 12452 360 13001 388
rect 6825 323 6883 329
rect 6825 289 6837 323
rect 6871 289 6883 323
rect 6825 283 6883 289
rect 7009 323 7067 329
rect 7009 289 7021 323
rect 7055 320 7067 323
rect 9030 320 9036 332
rect 7055 292 9036 320
rect 7055 289 7067 292
rect 7009 283 7067 289
rect 9030 280 9036 292
rect 9088 280 9094 332
rect 11238 320 11244 332
rect 10520 292 11244 320
rect 1302 252 1308 264
rect 1263 224 1308 252
rect 1302 212 1308 224
rect 1360 212 1366 264
rect 2958 212 2964 264
rect 3016 252 3022 264
rect 3145 255 3203 261
rect 3145 252 3157 255
rect 3016 224 3157 252
rect 3016 212 3022 224
rect 3145 221 3157 224
rect 3191 221 3203 255
rect 3145 215 3203 221
rect 5537 255 5595 261
rect 5537 221 5549 255
rect 5583 252 5595 255
rect 7282 252 7288 264
rect 5583 224 7288 252
rect 5583 221 5595 224
rect 5537 215 5595 221
rect 7282 212 7288 224
rect 7340 212 7346 264
rect 8846 252 8852 264
rect 8807 224 8852 252
rect 8846 212 8852 224
rect 8904 212 8910 264
rect 8941 255 8999 261
rect 8941 221 8953 255
rect 8987 252 8999 255
rect 9858 252 9864 264
rect 8987 224 9864 252
rect 8987 221 8999 224
rect 8941 215 8999 221
rect 9858 212 9864 224
rect 9916 212 9922 264
rect 10520 261 10548 292
rect 11238 280 11244 292
rect 11296 280 11302 332
rect 12452 329 12480 360
rect 12989 357 13001 360
rect 13035 357 13047 391
rect 12989 351 13047 357
rect 14844 360 17356 388
rect 12437 323 12495 329
rect 12437 289 12449 323
rect 12483 289 12495 323
rect 13170 320 13176 332
rect 12437 283 12495 289
rect 13004 292 13176 320
rect 10505 255 10563 261
rect 10505 221 10517 255
rect 10551 221 10563 255
rect 10505 215 10563 221
rect 10689 255 10747 261
rect 10689 221 10701 255
rect 10735 221 10747 255
rect 10689 215 10747 221
rect 6733 187 6791 193
rect 6733 153 6745 187
rect 6779 184 6791 187
rect 6914 184 6920 196
rect 6779 156 6920 184
rect 6779 153 6791 156
rect 6733 147 6791 153
rect 6914 144 6920 156
rect 6972 144 6978 196
rect 10704 184 10732 215
rect 10778 212 10784 264
rect 10836 252 10842 264
rect 10873 255 10931 261
rect 10873 252 10885 255
rect 10836 224 10885 252
rect 10836 212 10842 224
rect 10873 221 10885 224
rect 10919 221 10931 255
rect 10873 215 10931 221
rect 11149 255 11207 261
rect 11149 221 11161 255
rect 11195 252 11207 255
rect 11606 252 11612 264
rect 11195 224 11612 252
rect 11195 221 11207 224
rect 11149 215 11207 221
rect 11606 212 11612 224
rect 11664 252 11670 264
rect 12345 255 12403 261
rect 12345 252 12357 255
rect 11664 224 12357 252
rect 11664 212 11670 224
rect 12345 221 12357 224
rect 12391 221 12403 255
rect 12802 252 12808 264
rect 12763 224 12808 252
rect 12345 215 12403 221
rect 12802 212 12808 224
rect 12860 212 12866 264
rect 13004 261 13032 292
rect 13170 280 13176 292
rect 13228 320 13234 332
rect 14844 329 14872 360
rect 14829 323 14887 329
rect 14829 320 14841 323
rect 13228 292 14841 320
rect 13228 280 13234 292
rect 14829 289 14841 292
rect 14875 289 14887 323
rect 14829 283 14887 289
rect 16666 280 16672 332
rect 16724 320 16730 332
rect 16724 292 17080 320
rect 16724 280 16730 292
rect 12989 255 13047 261
rect 12989 221 13001 255
rect 13035 221 13047 255
rect 14734 252 14740 264
rect 14695 224 14740 252
rect 12989 215 13047 221
rect 14734 212 14740 224
rect 14792 212 14798 264
rect 16574 212 16580 264
rect 16632 252 16638 264
rect 17052 261 17080 292
rect 17328 261 17356 360
rect 16853 255 16911 261
rect 16853 252 16865 255
rect 16632 224 16865 252
rect 16632 212 16638 224
rect 16853 221 16865 224
rect 16899 221 16911 255
rect 16853 215 16911 221
rect 17037 255 17095 261
rect 17037 221 17049 255
rect 17083 221 17095 255
rect 17037 215 17095 221
rect 17313 255 17371 261
rect 17313 221 17325 255
rect 17359 252 17371 255
rect 17862 252 17868 264
rect 17359 224 17868 252
rect 17359 221 17371 224
rect 17313 215 17371 221
rect 17862 212 17868 224
rect 17920 212 17926 264
rect 10965 187 11023 193
rect 10704 156 10916 184
rect 10888 125 10916 156
rect 10965 153 10977 187
rect 11011 184 11023 187
rect 11330 184 11336 196
rect 11011 156 11336 184
rect 11011 153 11023 156
rect 10965 147 11023 153
rect 11330 144 11336 156
rect 11388 144 11394 196
rect 10873 119 10931 125
rect 10873 85 10885 119
rect 10919 85 10931 119
rect 10873 79 10931 85
rect 0 26 18860 48
rect 0 -26 4660 26
rect 4712 -26 4724 26
rect 4776 -26 4788 26
rect 4840 -26 4852 26
rect 4904 -26 4916 26
rect 4968 -26 7760 26
rect 7812 -26 7824 26
rect 7876 -26 7888 26
rect 7940 -26 7952 26
rect 8004 -26 8016 26
rect 8068 -26 10860 26
rect 10912 -26 10924 26
rect 10976 -26 10988 26
rect 11040 -26 11052 26
rect 11104 -26 11116 26
rect 11168 -26 13960 26
rect 14012 -26 14024 26
rect 14076 -26 14088 26
rect 14140 -26 14152 26
rect 14204 -26 14216 26
rect 14268 -26 17060 26
rect 17112 -26 17124 26
rect 17176 -26 17188 26
rect 17240 -26 17252 26
rect 17304 -26 17316 26
rect 17368 -26 18860 26
rect 0 -48 18860 -26
<< via1 >>
rect 4660 10854 4712 10906
rect 4724 10854 4776 10906
rect 4788 10854 4840 10906
rect 4852 10854 4904 10906
rect 4916 10854 4968 10906
rect 7760 10854 7812 10906
rect 7824 10854 7876 10906
rect 7888 10854 7940 10906
rect 7952 10854 8004 10906
rect 8016 10854 8068 10906
rect 10860 10854 10912 10906
rect 10924 10854 10976 10906
rect 10988 10854 11040 10906
rect 11052 10854 11104 10906
rect 11116 10854 11168 10906
rect 13960 10854 14012 10906
rect 14024 10854 14076 10906
rect 14088 10854 14140 10906
rect 14152 10854 14204 10906
rect 14216 10854 14268 10906
rect 17060 10854 17112 10906
rect 17124 10854 17176 10906
rect 17188 10854 17240 10906
rect 17252 10854 17304 10906
rect 17316 10854 17368 10906
rect 7104 10752 7156 10804
rect 8852 10752 8904 10804
rect 9956 10752 10008 10804
rect 12808 10752 12860 10804
rect 10876 10727 10928 10736
rect 10876 10693 10885 10727
rect 10885 10693 10919 10727
rect 10919 10693 10928 10727
rect 10876 10684 10928 10693
rect 13084 10684 13136 10736
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 3516 10616 3568 10668
rect 6092 10616 6144 10668
rect 2044 10548 2096 10600
rect 3792 10591 3844 10600
rect 3792 10557 3801 10591
rect 3801 10557 3835 10591
rect 3835 10557 3844 10591
rect 3792 10548 3844 10557
rect 8944 10591 8996 10600
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 11888 10616 11940 10668
rect 12900 10616 12952 10668
rect 11244 10548 11296 10600
rect 1952 10412 2004 10464
rect 5264 10412 5316 10464
rect 6000 10412 6052 10464
rect 7656 10412 7708 10464
rect 12808 10548 12860 10600
rect 15108 10616 15160 10668
rect 18052 10659 18104 10668
rect 18052 10625 18061 10659
rect 18061 10625 18095 10659
rect 18095 10625 18104 10659
rect 18052 10616 18104 10625
rect 18788 10616 18840 10668
rect 13268 10412 13320 10464
rect 14464 10455 14516 10464
rect 14464 10421 14473 10455
rect 14473 10421 14507 10455
rect 14507 10421 14516 10455
rect 14464 10412 14516 10421
rect 14740 10412 14792 10464
rect 15200 10412 15252 10464
rect 16948 10455 17000 10464
rect 16948 10421 16957 10455
rect 16957 10421 16991 10455
rect 16991 10421 17000 10455
rect 16948 10412 17000 10421
rect 3110 10310 3162 10362
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 3302 10310 3354 10362
rect 3366 10310 3418 10362
rect 6210 10310 6262 10362
rect 6274 10310 6326 10362
rect 6338 10310 6390 10362
rect 6402 10310 6454 10362
rect 6466 10310 6518 10362
rect 9310 10310 9362 10362
rect 9374 10310 9426 10362
rect 9438 10310 9490 10362
rect 9502 10310 9554 10362
rect 9566 10310 9618 10362
rect 12410 10310 12462 10362
rect 12474 10310 12526 10362
rect 12538 10310 12590 10362
rect 12602 10310 12654 10362
rect 12666 10310 12718 10362
rect 15510 10310 15562 10362
rect 15574 10310 15626 10362
rect 15638 10310 15690 10362
rect 15702 10310 15754 10362
rect 15766 10310 15818 10362
rect 3516 10208 3568 10260
rect 3792 10208 3844 10260
rect 6920 10208 6972 10260
rect 8852 10183 8904 10192
rect 296 10004 348 10056
rect 1952 10115 2004 10124
rect 1952 10081 1961 10115
rect 1961 10081 1995 10115
rect 1995 10081 2004 10115
rect 1952 10072 2004 10081
rect 6000 10072 6052 10124
rect 940 10047 992 10056
rect 940 10013 949 10047
rect 949 10013 983 10047
rect 983 10013 992 10047
rect 940 10004 992 10013
rect 388 9979 440 9988
rect 388 9945 397 9979
rect 397 9945 431 9979
rect 431 9945 440 9979
rect 388 9936 440 9945
rect 1216 10004 1268 10056
rect 3700 10047 3752 10056
rect 3700 10013 3709 10047
rect 3709 10013 3743 10047
rect 3743 10013 3752 10047
rect 3700 10004 3752 10013
rect 3884 10047 3936 10056
rect 3884 10013 3893 10047
rect 3893 10013 3927 10047
rect 3927 10013 3936 10047
rect 3884 10004 3936 10013
rect 6460 10047 6512 10056
rect 6460 10013 6469 10047
rect 6469 10013 6503 10047
rect 6503 10013 6512 10047
rect 6460 10004 6512 10013
rect 8852 10149 8861 10183
rect 8861 10149 8895 10183
rect 8895 10149 8904 10183
rect 8852 10140 8904 10149
rect 12808 10208 12860 10260
rect 13820 10208 13872 10260
rect 15108 10208 15160 10260
rect 18052 10208 18104 10260
rect 9220 10072 9272 10124
rect 11520 10072 11572 10124
rect 13268 10115 13320 10124
rect 13268 10081 13277 10115
rect 13277 10081 13311 10115
rect 13311 10081 13320 10115
rect 13268 10072 13320 10081
rect 14464 10072 14516 10124
rect 16948 10072 17000 10124
rect 16488 10004 16540 10056
rect 18604 10004 18656 10056
rect 664 9868 716 9920
rect 1584 9979 1636 9988
rect 1584 9945 1593 9979
rect 1593 9945 1627 9979
rect 1627 9945 1636 9979
rect 1584 9936 1636 9945
rect 2596 9868 2648 9920
rect 7472 9936 7524 9988
rect 3608 9868 3660 9920
rect 10232 9868 10284 9920
rect 10692 9911 10744 9920
rect 10692 9877 10701 9911
rect 10701 9877 10735 9911
rect 10735 9877 10744 9911
rect 10692 9868 10744 9877
rect 10876 9936 10928 9988
rect 12440 9868 12492 9920
rect 16120 9868 16172 9920
rect 18328 9911 18380 9920
rect 18328 9877 18337 9911
rect 18337 9877 18371 9911
rect 18371 9877 18380 9911
rect 18328 9868 18380 9877
rect 4660 9766 4712 9818
rect 4724 9766 4776 9818
rect 4788 9766 4840 9818
rect 4852 9766 4904 9818
rect 4916 9766 4968 9818
rect 7760 9766 7812 9818
rect 7824 9766 7876 9818
rect 7888 9766 7940 9818
rect 7952 9766 8004 9818
rect 8016 9766 8068 9818
rect 10860 9766 10912 9818
rect 10924 9766 10976 9818
rect 10988 9766 11040 9818
rect 11052 9766 11104 9818
rect 11116 9766 11168 9818
rect 13960 9766 14012 9818
rect 14024 9766 14076 9818
rect 14088 9766 14140 9818
rect 14152 9766 14204 9818
rect 14216 9766 14268 9818
rect 17060 9766 17112 9818
rect 17124 9766 17176 9818
rect 17188 9766 17240 9818
rect 17252 9766 17304 9818
rect 17316 9766 17368 9818
rect 2136 9664 2188 9716
rect 2964 9664 3016 9716
rect 5264 9707 5316 9716
rect 5264 9673 5273 9707
rect 5273 9673 5307 9707
rect 5307 9673 5316 9707
rect 5264 9664 5316 9673
rect 6460 9707 6512 9716
rect 2228 9596 2280 9648
rect 388 9528 440 9580
rect 664 9571 716 9580
rect 664 9537 673 9571
rect 673 9537 707 9571
rect 707 9537 716 9571
rect 664 9528 716 9537
rect 1584 9528 1636 9580
rect 2688 9596 2740 9648
rect 1216 9460 1268 9512
rect 2596 9571 2648 9580
rect 2596 9537 2605 9571
rect 2605 9537 2639 9571
rect 2639 9537 2648 9571
rect 2596 9528 2648 9537
rect 2872 9571 2924 9580
rect 2872 9537 2881 9571
rect 2881 9537 2915 9571
rect 2915 9537 2924 9571
rect 3700 9596 3752 9648
rect 2872 9528 2924 9537
rect 3516 9528 3568 9580
rect 5632 9596 5684 9648
rect 6460 9673 6469 9707
rect 6469 9673 6503 9707
rect 6503 9673 6512 9707
rect 6460 9664 6512 9673
rect 11244 9707 11296 9716
rect 6644 9596 6696 9648
rect 8852 9596 8904 9648
rect 11244 9673 11253 9707
rect 11253 9673 11287 9707
rect 11287 9673 11296 9707
rect 11244 9664 11296 9673
rect 12440 9664 12492 9716
rect 16580 9664 16632 9716
rect 9864 9596 9916 9648
rect 16120 9596 16172 9648
rect 2228 9367 2280 9376
rect 2228 9333 2237 9367
rect 2237 9333 2271 9367
rect 2271 9333 2280 9367
rect 2228 9324 2280 9333
rect 2872 9392 2924 9444
rect 3884 9392 3936 9444
rect 5448 9503 5500 9512
rect 5448 9469 5457 9503
rect 5457 9469 5491 9503
rect 5491 9469 5500 9503
rect 5448 9460 5500 9469
rect 3976 9324 4028 9376
rect 5172 9392 5224 9444
rect 6000 9528 6052 9580
rect 6920 9528 6972 9580
rect 7472 9571 7524 9580
rect 7472 9537 7481 9571
rect 7481 9537 7515 9571
rect 7515 9537 7524 9571
rect 7472 9528 7524 9537
rect 9772 9528 9824 9580
rect 14740 9571 14792 9580
rect 14740 9537 14749 9571
rect 14749 9537 14783 9571
rect 14783 9537 14792 9571
rect 14740 9528 14792 9537
rect 15200 9528 15252 9580
rect 6092 9460 6144 9512
rect 8484 9460 8536 9512
rect 9036 9460 9088 9512
rect 8852 9392 8904 9444
rect 9864 9392 9916 9444
rect 12256 9460 12308 9512
rect 18328 9460 18380 9512
rect 4896 9367 4948 9376
rect 4896 9333 4905 9367
rect 4905 9333 4939 9367
rect 4939 9333 4948 9367
rect 4896 9324 4948 9333
rect 5540 9324 5592 9376
rect 7472 9324 7524 9376
rect 9036 9324 9088 9376
rect 9772 9367 9824 9376
rect 9772 9333 9781 9367
rect 9781 9333 9815 9367
rect 9815 9333 9824 9367
rect 9772 9324 9824 9333
rect 9956 9324 10008 9376
rect 11336 9324 11388 9376
rect 12164 9367 12216 9376
rect 12164 9333 12173 9367
rect 12173 9333 12207 9367
rect 12207 9333 12216 9367
rect 12164 9324 12216 9333
rect 14740 9392 14792 9444
rect 12992 9324 13044 9376
rect 15292 9324 15344 9376
rect 16120 9324 16172 9376
rect 3110 9222 3162 9274
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 3302 9222 3354 9274
rect 3366 9222 3418 9274
rect 6210 9222 6262 9274
rect 6274 9222 6326 9274
rect 6338 9222 6390 9274
rect 6402 9222 6454 9274
rect 6466 9222 6518 9274
rect 9310 9222 9362 9274
rect 9374 9222 9426 9274
rect 9438 9222 9490 9274
rect 9502 9222 9554 9274
rect 9566 9222 9618 9274
rect 12410 9222 12462 9274
rect 12474 9222 12526 9274
rect 12538 9222 12590 9274
rect 12602 9222 12654 9274
rect 12666 9222 12718 9274
rect 15510 9222 15562 9274
rect 15574 9222 15626 9274
rect 15638 9222 15690 9274
rect 15702 9222 15754 9274
rect 15766 9222 15818 9274
rect 940 9120 992 9172
rect 1400 9163 1452 9172
rect 1400 9129 1409 9163
rect 1409 9129 1443 9163
rect 1443 9129 1452 9163
rect 1400 9120 1452 9129
rect 6000 9120 6052 9172
rect 8484 9163 8536 9172
rect 8484 9129 8493 9163
rect 8493 9129 8527 9163
rect 8527 9129 8536 9163
rect 8484 9120 8536 9129
rect 11888 9163 11940 9172
rect 2596 9052 2648 9104
rect 6644 9052 6696 9104
rect 7196 9052 7248 9104
rect 10508 9095 10560 9104
rect 2136 8984 2188 9036
rect 3700 8984 3752 9036
rect 1400 8916 1452 8968
rect 2228 8916 2280 8968
rect 3608 8916 3660 8968
rect 4896 8916 4948 8968
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 8852 8984 8904 9036
rect 10508 9061 10517 9095
rect 10517 9061 10551 9095
rect 10551 9061 10560 9095
rect 10508 9052 10560 9061
rect 10324 9027 10376 9036
rect 5632 8916 5684 8925
rect 7288 8916 7340 8968
rect 7472 8916 7524 8968
rect 2320 8848 2372 8900
rect 2136 8780 2188 8832
rect 2780 8848 2832 8900
rect 2596 8780 2648 8832
rect 4068 8848 4120 8900
rect 5448 8848 5500 8900
rect 6092 8848 6144 8900
rect 6552 8848 6604 8900
rect 7104 8891 7156 8900
rect 7104 8857 7113 8891
rect 7113 8857 7147 8891
rect 7147 8857 7156 8891
rect 7104 8848 7156 8857
rect 8116 8916 8168 8968
rect 10324 8993 10333 9027
rect 10333 8993 10367 9027
rect 10367 8993 10376 9027
rect 10324 8984 10376 8993
rect 8484 8848 8536 8900
rect 9036 8848 9088 8900
rect 9404 8916 9456 8968
rect 5724 8780 5776 8832
rect 7564 8780 7616 8832
rect 9864 8848 9916 8900
rect 10784 8916 10836 8968
rect 11888 9129 11897 9163
rect 11897 9129 11931 9163
rect 11931 9129 11940 9163
rect 11888 9120 11940 9129
rect 12072 9120 12124 9172
rect 11428 9027 11480 9036
rect 11428 8993 11437 9027
rect 11437 8993 11471 9027
rect 11471 8993 11480 9027
rect 11428 8984 11480 8993
rect 11336 8916 11388 8968
rect 12440 9052 12492 9104
rect 12900 9052 12952 9104
rect 12808 8984 12860 9036
rect 14464 8984 14516 9036
rect 11980 8848 12032 8900
rect 12716 8959 12768 8968
rect 12716 8925 12725 8959
rect 12725 8925 12759 8959
rect 12759 8925 12768 8959
rect 12716 8916 12768 8925
rect 9956 8780 10008 8832
rect 10140 8823 10192 8832
rect 10140 8789 10149 8823
rect 10149 8789 10183 8823
rect 10183 8789 10192 8823
rect 10140 8780 10192 8789
rect 12072 8780 12124 8832
rect 12256 8780 12308 8832
rect 12624 8780 12676 8832
rect 17408 9120 17460 9172
rect 14740 8984 14792 9036
rect 13176 8848 13228 8900
rect 13636 8780 13688 8832
rect 15200 8848 15252 8900
rect 14924 8780 14976 8832
rect 15936 8916 15988 8968
rect 17868 8959 17920 8968
rect 17868 8925 17877 8959
rect 17877 8925 17911 8959
rect 17911 8925 17920 8959
rect 17868 8916 17920 8925
rect 16212 8780 16264 8832
rect 4660 8678 4712 8730
rect 4724 8678 4776 8730
rect 4788 8678 4840 8730
rect 4852 8678 4904 8730
rect 4916 8678 4968 8730
rect 7760 8678 7812 8730
rect 7824 8678 7876 8730
rect 7888 8678 7940 8730
rect 7952 8678 8004 8730
rect 8016 8678 8068 8730
rect 10860 8678 10912 8730
rect 10924 8678 10976 8730
rect 10988 8678 11040 8730
rect 11052 8678 11104 8730
rect 11116 8678 11168 8730
rect 13960 8678 14012 8730
rect 14024 8678 14076 8730
rect 14088 8678 14140 8730
rect 14152 8678 14204 8730
rect 14216 8678 14268 8730
rect 17060 8678 17112 8730
rect 17124 8678 17176 8730
rect 17188 8678 17240 8730
rect 17252 8678 17304 8730
rect 17316 8678 17368 8730
rect 2044 8576 2096 8628
rect 2320 8576 2372 8628
rect 6644 8576 6696 8628
rect 2228 8508 2280 8560
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 2596 8508 2648 8560
rect 2780 8508 2832 8560
rect 2688 8483 2740 8492
rect 2688 8449 2697 8483
rect 2697 8449 2731 8483
rect 2731 8449 2740 8483
rect 2688 8440 2740 8449
rect 296 8415 348 8424
rect 296 8381 305 8415
rect 305 8381 339 8415
rect 339 8381 348 8415
rect 296 8372 348 8381
rect 572 8415 624 8424
rect 572 8381 581 8415
rect 581 8381 615 8415
rect 615 8381 624 8415
rect 572 8372 624 8381
rect 2872 8372 2924 8424
rect 5172 8483 5224 8492
rect 5172 8449 5181 8483
rect 5181 8449 5215 8483
rect 5215 8449 5224 8483
rect 5172 8440 5224 8449
rect 5540 8508 5592 8560
rect 6552 8508 6604 8560
rect 8760 8576 8812 8628
rect 8944 8576 8996 8628
rect 9588 8576 9640 8628
rect 10232 8576 10284 8628
rect 10692 8576 10744 8628
rect 12164 8576 12216 8628
rect 12716 8576 12768 8628
rect 13176 8619 13228 8628
rect 13176 8585 13185 8619
rect 13185 8585 13219 8619
rect 13219 8585 13228 8619
rect 13176 8576 13228 8585
rect 13636 8619 13688 8628
rect 13636 8585 13645 8619
rect 13645 8585 13679 8619
rect 13679 8585 13688 8619
rect 13636 8576 13688 8585
rect 14464 8576 14516 8628
rect 5724 8483 5776 8492
rect 5724 8449 5733 8483
rect 5733 8449 5767 8483
rect 5767 8449 5776 8483
rect 7656 8508 7708 8560
rect 5724 8440 5776 8449
rect 3700 8415 3752 8424
rect 3700 8381 3709 8415
rect 3709 8381 3743 8415
rect 3743 8381 3752 8415
rect 3700 8372 3752 8381
rect 3884 8304 3936 8356
rect 4068 8304 4120 8356
rect 5816 8372 5868 8424
rect 2044 8279 2096 8288
rect 2044 8245 2053 8279
rect 2053 8245 2087 8279
rect 2087 8245 2096 8279
rect 2044 8236 2096 8245
rect 2964 8236 3016 8288
rect 5172 8236 5224 8288
rect 5908 8279 5960 8288
rect 5908 8245 5917 8279
rect 5917 8245 5951 8279
rect 5951 8245 5960 8279
rect 10508 8508 10560 8560
rect 8208 8440 8260 8492
rect 7196 8372 7248 8424
rect 7472 8415 7524 8424
rect 7472 8381 7481 8415
rect 7481 8381 7515 8415
rect 7515 8381 7524 8415
rect 7472 8372 7524 8381
rect 8760 8372 8812 8424
rect 9404 8372 9456 8424
rect 9588 8440 9640 8492
rect 9864 8440 9916 8492
rect 11796 8440 11848 8492
rect 10600 8372 10652 8424
rect 11520 8372 11572 8424
rect 11980 8440 12032 8492
rect 12348 8508 12400 8560
rect 12900 8483 12952 8492
rect 12900 8449 12909 8483
rect 12909 8449 12943 8483
rect 12943 8449 12952 8483
rect 16212 8508 16264 8560
rect 16948 8508 17000 8560
rect 12900 8440 12952 8449
rect 14924 8440 14976 8492
rect 13820 8415 13872 8424
rect 13820 8381 13829 8415
rect 13829 8381 13863 8415
rect 13863 8381 13872 8415
rect 13820 8372 13872 8381
rect 11152 8304 11204 8356
rect 12348 8304 12400 8356
rect 12624 8304 12676 8356
rect 5908 8236 5960 8245
rect 10140 8236 10192 8288
rect 11428 8236 11480 8288
rect 11888 8236 11940 8288
rect 12900 8304 12952 8356
rect 14004 8304 14056 8356
rect 14648 8304 14700 8356
rect 16580 8372 16632 8424
rect 18604 8440 18656 8492
rect 17408 8415 17460 8424
rect 17408 8381 17417 8415
rect 17417 8381 17451 8415
rect 17451 8381 17460 8415
rect 17408 8372 17460 8381
rect 14832 8236 14884 8288
rect 16764 8236 16816 8288
rect 3110 8134 3162 8186
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 3302 8134 3354 8186
rect 3366 8134 3418 8186
rect 6210 8134 6262 8186
rect 6274 8134 6326 8186
rect 6338 8134 6390 8186
rect 6402 8134 6454 8186
rect 6466 8134 6518 8186
rect 9310 8134 9362 8186
rect 9374 8134 9426 8186
rect 9438 8134 9490 8186
rect 9502 8134 9554 8186
rect 9566 8134 9618 8186
rect 12410 8134 12462 8186
rect 12474 8134 12526 8186
rect 12538 8134 12590 8186
rect 12602 8134 12654 8186
rect 12666 8134 12718 8186
rect 15510 8134 15562 8186
rect 15574 8134 15626 8186
rect 15638 8134 15690 8186
rect 15702 8134 15754 8186
rect 15766 8134 15818 8186
rect 572 8032 624 8084
rect 2136 8032 2188 8084
rect 2320 8032 2372 8084
rect 2504 8075 2556 8084
rect 2504 8041 2513 8075
rect 2513 8041 2547 8075
rect 2547 8041 2556 8075
rect 2504 8032 2556 8041
rect 4252 8032 4304 8084
rect 9772 8032 9824 8084
rect 11796 8075 11848 8084
rect 11796 8041 11805 8075
rect 11805 8041 11839 8075
rect 11839 8041 11848 8075
rect 11796 8032 11848 8041
rect 1308 7939 1360 7948
rect 1308 7905 1317 7939
rect 1317 7905 1351 7939
rect 1351 7905 1360 7939
rect 1308 7896 1360 7905
rect 3700 7964 3752 8016
rect 5540 7964 5592 8016
rect 2964 7896 3016 7948
rect 7564 7896 7616 7948
rect 8852 7939 8904 7948
rect 8852 7905 8861 7939
rect 8861 7905 8895 7939
rect 8895 7905 8904 7939
rect 8852 7896 8904 7905
rect 11428 7939 11480 7948
rect 11428 7905 11437 7939
rect 11437 7905 11471 7939
rect 11471 7905 11480 7939
rect 11428 7896 11480 7905
rect 1952 7828 2004 7880
rect 3700 7828 3752 7880
rect 6092 7828 6144 7880
rect 11152 7828 11204 7880
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 11704 7828 11756 7837
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 2504 7760 2556 7812
rect 7380 7760 7432 7812
rect 18512 8032 18564 8084
rect 12072 7964 12124 8016
rect 13636 7964 13688 8016
rect 15936 7964 15988 8016
rect 14372 7939 14424 7948
rect 3792 7692 3844 7744
rect 6920 7692 6972 7744
rect 7104 7692 7156 7744
rect 8208 7692 8260 7744
rect 9128 7692 9180 7744
rect 11244 7692 11296 7744
rect 14372 7905 14381 7939
rect 14381 7905 14415 7939
rect 14415 7905 14424 7939
rect 14372 7896 14424 7905
rect 12164 7760 12216 7812
rect 14004 7828 14056 7880
rect 14648 7871 14700 7880
rect 14648 7837 14657 7871
rect 14657 7837 14691 7871
rect 14691 7837 14700 7871
rect 14648 7828 14700 7837
rect 14832 7828 14884 7880
rect 16580 7896 16632 7948
rect 16764 7896 16816 7948
rect 17868 7871 17920 7880
rect 14740 7760 14792 7812
rect 12256 7692 12308 7744
rect 17868 7837 17877 7871
rect 17877 7837 17911 7871
rect 17911 7837 17920 7871
rect 17868 7828 17920 7837
rect 16304 7760 16356 7812
rect 4660 7590 4712 7642
rect 4724 7590 4776 7642
rect 4788 7590 4840 7642
rect 4852 7590 4904 7642
rect 4916 7590 4968 7642
rect 7760 7590 7812 7642
rect 7824 7590 7876 7642
rect 7888 7590 7940 7642
rect 7952 7590 8004 7642
rect 8016 7590 8068 7642
rect 10860 7590 10912 7642
rect 10924 7590 10976 7642
rect 10988 7590 11040 7642
rect 11052 7590 11104 7642
rect 11116 7590 11168 7642
rect 13960 7590 14012 7642
rect 14024 7590 14076 7642
rect 14088 7590 14140 7642
rect 14152 7590 14204 7642
rect 14216 7590 14268 7642
rect 17060 7590 17112 7642
rect 17124 7590 17176 7642
rect 17188 7590 17240 7642
rect 17252 7590 17304 7642
rect 17316 7590 17368 7642
rect 1308 7488 1360 7540
rect 1952 7463 2004 7472
rect 1952 7429 1961 7463
rect 1961 7429 1995 7463
rect 1995 7429 2004 7463
rect 1952 7420 2004 7429
rect 3792 7420 3844 7472
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 2320 7395 2372 7404
rect 2320 7361 2329 7395
rect 2329 7361 2363 7395
rect 2363 7361 2372 7395
rect 2320 7352 2372 7361
rect 2504 7352 2556 7404
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 2596 7327 2648 7336
rect 2596 7293 2605 7327
rect 2605 7293 2639 7327
rect 2639 7293 2648 7327
rect 2596 7284 2648 7293
rect 3884 7284 3936 7336
rect 4344 7352 4396 7404
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 5632 7488 5684 7540
rect 7288 7488 7340 7540
rect 8484 7531 8536 7540
rect 8484 7497 8493 7531
rect 8493 7497 8527 7531
rect 8527 7497 8536 7531
rect 8484 7488 8536 7497
rect 8852 7488 8904 7540
rect 8944 7488 8996 7540
rect 11244 7488 11296 7540
rect 12072 7488 12124 7540
rect 4804 7284 4856 7336
rect 5172 7398 5224 7404
rect 5172 7364 5181 7398
rect 5181 7364 5215 7398
rect 5215 7364 5224 7398
rect 5172 7352 5224 7364
rect 5356 7352 5408 7404
rect 5724 7352 5776 7404
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 5540 7284 5592 7336
rect 6000 7284 6052 7336
rect 6552 7284 6604 7336
rect 7656 7420 7708 7472
rect 8116 7420 8168 7472
rect 7012 7284 7064 7336
rect 7380 7284 7432 7336
rect 8208 7284 8260 7336
rect 9128 7352 9180 7404
rect 11060 7395 11112 7404
rect 11060 7361 11069 7395
rect 11069 7361 11103 7395
rect 11103 7361 11112 7395
rect 11060 7352 11112 7361
rect 11704 7352 11756 7404
rect 8944 7327 8996 7336
rect 8944 7293 8953 7327
rect 8953 7293 8987 7327
rect 8987 7293 8996 7327
rect 8944 7284 8996 7293
rect 9036 7327 9088 7336
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 10324 7284 10376 7336
rect 2964 7148 3016 7200
rect 4252 7191 4304 7200
rect 4252 7157 4261 7191
rect 4261 7157 4295 7191
rect 4295 7157 4304 7191
rect 4252 7148 4304 7157
rect 7380 7148 7432 7200
rect 7564 7148 7616 7200
rect 11428 7284 11480 7336
rect 10784 7216 10836 7268
rect 12164 7352 12216 7404
rect 12256 7284 12308 7336
rect 12900 7352 12952 7404
rect 14188 7463 14240 7472
rect 14188 7429 14197 7463
rect 14197 7429 14231 7463
rect 14231 7429 14240 7463
rect 14188 7420 14240 7429
rect 14004 7395 14056 7404
rect 14372 7420 14424 7472
rect 12808 7284 12860 7336
rect 14004 7361 14032 7395
rect 14032 7361 14056 7395
rect 14004 7352 14056 7361
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 16948 7395 17000 7404
rect 16948 7361 16957 7395
rect 16957 7361 16991 7395
rect 16991 7361 17000 7395
rect 16948 7352 17000 7361
rect 14096 7216 14148 7268
rect 9036 7148 9088 7200
rect 11428 7191 11480 7200
rect 11428 7157 11437 7191
rect 11437 7157 11471 7191
rect 11471 7157 11480 7191
rect 11428 7148 11480 7157
rect 12164 7191 12216 7200
rect 12164 7157 12173 7191
rect 12173 7157 12207 7191
rect 12207 7157 12216 7191
rect 12164 7148 12216 7157
rect 12256 7191 12308 7200
rect 12256 7157 12265 7191
rect 12265 7157 12299 7191
rect 12299 7157 12308 7191
rect 12256 7148 12308 7157
rect 16304 7148 16356 7200
rect 3110 7046 3162 7098
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 3302 7046 3354 7098
rect 3366 7046 3418 7098
rect 6210 7046 6262 7098
rect 6274 7046 6326 7098
rect 6338 7046 6390 7098
rect 6402 7046 6454 7098
rect 6466 7046 6518 7098
rect 9310 7046 9362 7098
rect 9374 7046 9426 7098
rect 9438 7046 9490 7098
rect 9502 7046 9554 7098
rect 9566 7046 9618 7098
rect 12410 7046 12462 7098
rect 12474 7046 12526 7098
rect 12538 7046 12590 7098
rect 12602 7046 12654 7098
rect 12666 7046 12718 7098
rect 15510 7046 15562 7098
rect 15574 7046 15626 7098
rect 15638 7046 15690 7098
rect 15702 7046 15754 7098
rect 15766 7046 15818 7098
rect 3884 6944 3936 6996
rect 6552 6944 6604 6996
rect 7380 6944 7432 6996
rect 8208 6944 8260 6996
rect 10784 6944 10836 6996
rect 12256 6944 12308 6996
rect 14096 6987 14148 6996
rect 14096 6953 14105 6987
rect 14105 6953 14139 6987
rect 14139 6953 14148 6987
rect 14096 6944 14148 6953
rect 4436 6876 4488 6928
rect 2504 6808 2556 6860
rect 3700 6808 3752 6860
rect 3976 6808 4028 6860
rect 2412 6783 2464 6792
rect 572 6604 624 6656
rect 2412 6749 2421 6783
rect 2421 6749 2455 6783
rect 2455 6749 2464 6783
rect 2412 6740 2464 6749
rect 2872 6740 2924 6792
rect 4896 6808 4948 6860
rect 5172 6876 5224 6928
rect 7012 6876 7064 6928
rect 4344 6672 4396 6724
rect 4528 6672 4580 6724
rect 5356 6740 5408 6792
rect 6000 6740 6052 6792
rect 7288 6808 7340 6860
rect 10324 6740 10376 6792
rect 11428 6740 11480 6792
rect 12808 6808 12860 6860
rect 4804 6672 4856 6724
rect 5724 6672 5776 6724
rect 2964 6604 3016 6656
rect 7012 6672 7064 6724
rect 8852 6715 8904 6724
rect 8852 6681 8861 6715
rect 8861 6681 8895 6715
rect 8895 6681 8904 6715
rect 8852 6672 8904 6681
rect 10692 6672 10744 6724
rect 8760 6604 8812 6656
rect 10968 6672 11020 6724
rect 12900 6740 12952 6792
rect 13544 6740 13596 6792
rect 14280 6876 14332 6928
rect 14372 6808 14424 6860
rect 16948 6808 17000 6860
rect 17868 6851 17920 6860
rect 17868 6817 17877 6851
rect 17877 6817 17911 6851
rect 17911 6817 17920 6851
rect 17868 6808 17920 6817
rect 14004 6672 14056 6724
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 15844 6715 15896 6724
rect 15844 6681 15853 6715
rect 15853 6681 15887 6715
rect 15887 6681 15896 6715
rect 15844 6672 15896 6681
rect 16304 6672 16356 6724
rect 17500 6672 17552 6724
rect 12808 6604 12860 6656
rect 14556 6604 14608 6656
rect 15108 6647 15160 6656
rect 15108 6613 15117 6647
rect 15117 6613 15151 6647
rect 15151 6613 15160 6647
rect 15108 6604 15160 6613
rect 15936 6604 15988 6656
rect 18328 6647 18380 6656
rect 18328 6613 18337 6647
rect 18337 6613 18371 6647
rect 18371 6613 18380 6647
rect 18328 6604 18380 6613
rect 4660 6502 4712 6554
rect 4724 6502 4776 6554
rect 4788 6502 4840 6554
rect 4852 6502 4904 6554
rect 4916 6502 4968 6554
rect 7760 6502 7812 6554
rect 7824 6502 7876 6554
rect 7888 6502 7940 6554
rect 7952 6502 8004 6554
rect 8016 6502 8068 6554
rect 10860 6502 10912 6554
rect 10924 6502 10976 6554
rect 10988 6502 11040 6554
rect 11052 6502 11104 6554
rect 11116 6502 11168 6554
rect 13960 6502 14012 6554
rect 14024 6502 14076 6554
rect 14088 6502 14140 6554
rect 14152 6502 14204 6554
rect 14216 6502 14268 6554
rect 17060 6502 17112 6554
rect 17124 6502 17176 6554
rect 17188 6502 17240 6554
rect 17252 6502 17304 6554
rect 17316 6502 17368 6554
rect 2412 6400 2464 6452
rect 2596 6443 2648 6452
rect 2596 6409 2605 6443
rect 2605 6409 2639 6443
rect 2639 6409 2648 6443
rect 2596 6400 2648 6409
rect 4252 6400 4304 6452
rect 8852 6400 8904 6452
rect 13544 6400 13596 6452
rect 15108 6400 15160 6452
rect 572 6375 624 6384
rect 572 6341 581 6375
rect 581 6341 615 6375
rect 615 6341 624 6375
rect 572 6332 624 6341
rect 2228 6332 2280 6384
rect 4344 6332 4396 6384
rect 2688 6307 2740 6316
rect 296 6239 348 6248
rect 296 6205 305 6239
rect 305 6205 339 6239
rect 339 6205 348 6239
rect 296 6196 348 6205
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 2688 6264 2740 6273
rect 2780 6264 2832 6316
rect 4068 6264 4120 6316
rect 2872 6196 2924 6248
rect 3700 6239 3752 6248
rect 3700 6205 3709 6239
rect 3709 6205 3743 6239
rect 3743 6205 3752 6239
rect 3700 6196 3752 6205
rect 4528 6196 4580 6248
rect 2504 6128 2556 6180
rect 5448 6128 5500 6180
rect 5632 6128 5684 6180
rect 6000 6264 6052 6316
rect 7656 6307 7708 6316
rect 7656 6273 7665 6307
rect 7665 6273 7699 6307
rect 7699 6273 7708 6307
rect 7656 6264 7708 6273
rect 12164 6332 12216 6384
rect 16212 6400 16264 6452
rect 16948 6443 17000 6452
rect 16948 6409 16957 6443
rect 16957 6409 16991 6443
rect 16991 6409 17000 6443
rect 16948 6400 17000 6409
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 13820 6307 13872 6316
rect 6552 6239 6604 6248
rect 6552 6205 6561 6239
rect 6561 6205 6595 6239
rect 6595 6205 6604 6239
rect 6552 6196 6604 6205
rect 7564 6196 7616 6248
rect 8392 6196 8444 6248
rect 8944 6128 8996 6180
rect 13820 6273 13829 6307
rect 13829 6273 13863 6307
rect 13863 6273 13872 6307
rect 13820 6264 13872 6273
rect 14648 6264 14700 6316
rect 16304 6264 16356 6316
rect 16488 6264 16540 6316
rect 12808 6239 12860 6248
rect 12808 6205 12817 6239
rect 12817 6205 12851 6239
rect 12851 6205 12860 6239
rect 12808 6196 12860 6205
rect 14372 6196 14424 6248
rect 14464 6196 14516 6248
rect 16580 6196 16632 6248
rect 17408 6196 17460 6248
rect 16212 6128 16264 6180
rect 2228 6103 2280 6112
rect 2228 6069 2237 6103
rect 2237 6069 2271 6103
rect 2271 6069 2280 6103
rect 2228 6060 2280 6069
rect 2964 6060 3016 6112
rect 4436 6060 4488 6112
rect 5540 6060 5592 6112
rect 8300 6103 8352 6112
rect 8300 6069 8309 6103
rect 8309 6069 8343 6103
rect 8343 6069 8352 6103
rect 8300 6060 8352 6069
rect 8576 6060 8628 6112
rect 8668 6103 8720 6112
rect 8668 6069 8677 6103
rect 8677 6069 8711 6103
rect 8711 6069 8720 6103
rect 9036 6103 9088 6112
rect 8668 6060 8720 6069
rect 9036 6069 9045 6103
rect 9045 6069 9079 6103
rect 9079 6069 9088 6103
rect 9036 6060 9088 6069
rect 10692 6060 10744 6112
rect 11704 6103 11756 6112
rect 11704 6069 11713 6103
rect 11713 6069 11747 6103
rect 11747 6069 11756 6103
rect 11704 6060 11756 6069
rect 14280 6060 14332 6112
rect 14740 6060 14792 6112
rect 15844 6060 15896 6112
rect 3110 5958 3162 6010
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 3302 5958 3354 6010
rect 3366 5958 3418 6010
rect 6210 5958 6262 6010
rect 6274 5958 6326 6010
rect 6338 5958 6390 6010
rect 6402 5958 6454 6010
rect 6466 5958 6518 6010
rect 9310 5958 9362 6010
rect 9374 5958 9426 6010
rect 9438 5958 9490 6010
rect 9502 5958 9554 6010
rect 9566 5958 9618 6010
rect 12410 5958 12462 6010
rect 12474 5958 12526 6010
rect 12538 5958 12590 6010
rect 12602 5958 12654 6010
rect 12666 5958 12718 6010
rect 15510 5958 15562 6010
rect 15574 5958 15626 6010
rect 15638 5958 15690 6010
rect 15702 5958 15754 6010
rect 15766 5958 15818 6010
rect 2872 5856 2924 5908
rect 4436 5856 4488 5908
rect 6552 5899 6604 5908
rect 296 5720 348 5772
rect 6092 5720 6144 5772
rect 6552 5865 6561 5899
rect 6561 5865 6595 5899
rect 6595 5865 6604 5899
rect 6552 5856 6604 5865
rect 8300 5899 8352 5908
rect 8300 5865 8309 5899
rect 8309 5865 8343 5899
rect 8343 5865 8352 5899
rect 8300 5856 8352 5865
rect 6276 5788 6328 5840
rect 1216 5584 1268 5636
rect 5724 5652 5776 5704
rect 4436 5627 4488 5636
rect 2228 5516 2280 5568
rect 4436 5593 4445 5627
rect 4445 5593 4479 5627
rect 4479 5593 4488 5627
rect 4436 5584 4488 5593
rect 8024 5652 8076 5704
rect 8668 5652 8720 5704
rect 15384 5856 15436 5908
rect 16948 5856 17000 5908
rect 11428 5720 11480 5772
rect 14464 5788 14516 5840
rect 14280 5763 14332 5772
rect 14280 5729 14289 5763
rect 14289 5729 14323 5763
rect 14323 5729 14332 5763
rect 14280 5720 14332 5729
rect 16488 5788 16540 5840
rect 15844 5720 15896 5772
rect 17500 5720 17552 5772
rect 18328 5720 18380 5772
rect 14556 5695 14608 5704
rect 3516 5516 3568 5568
rect 8208 5584 8260 5636
rect 11704 5584 11756 5636
rect 5908 5559 5960 5568
rect 5908 5525 5917 5559
rect 5917 5525 5951 5559
rect 5951 5525 5960 5559
rect 5908 5516 5960 5525
rect 9312 5516 9364 5568
rect 10692 5516 10744 5568
rect 12348 5516 12400 5568
rect 12808 5516 12860 5568
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 14648 5584 14700 5636
rect 13820 5559 13872 5568
rect 13820 5525 13829 5559
rect 13829 5525 13863 5559
rect 13863 5525 13872 5559
rect 13820 5516 13872 5525
rect 14372 5516 14424 5568
rect 16212 5652 16264 5704
rect 17868 5695 17920 5704
rect 17868 5661 17877 5695
rect 17877 5661 17911 5695
rect 17911 5661 17920 5695
rect 17868 5652 17920 5661
rect 18512 5695 18564 5704
rect 18512 5661 18521 5695
rect 18521 5661 18555 5695
rect 18555 5661 18564 5695
rect 18512 5652 18564 5661
rect 16120 5584 16172 5636
rect 15016 5559 15068 5568
rect 15016 5525 15025 5559
rect 15025 5525 15059 5559
rect 15059 5525 15068 5559
rect 15016 5516 15068 5525
rect 18052 5516 18104 5568
rect 4660 5414 4712 5466
rect 4724 5414 4776 5466
rect 4788 5414 4840 5466
rect 4852 5414 4904 5466
rect 4916 5414 4968 5466
rect 7760 5414 7812 5466
rect 7824 5414 7876 5466
rect 7888 5414 7940 5466
rect 7952 5414 8004 5466
rect 8016 5414 8068 5466
rect 10860 5414 10912 5466
rect 10924 5414 10976 5466
rect 10988 5414 11040 5466
rect 11052 5414 11104 5466
rect 11116 5414 11168 5466
rect 13960 5414 14012 5466
rect 14024 5414 14076 5466
rect 14088 5414 14140 5466
rect 14152 5414 14204 5466
rect 14216 5414 14268 5466
rect 17060 5414 17112 5466
rect 17124 5414 17176 5466
rect 17188 5414 17240 5466
rect 17252 5414 17304 5466
rect 17316 5414 17368 5466
rect 1216 5355 1268 5364
rect 1216 5321 1225 5355
rect 1225 5321 1259 5355
rect 1259 5321 1268 5355
rect 1216 5312 1268 5321
rect 2780 5312 2832 5364
rect 2964 5355 3016 5364
rect 2964 5321 2973 5355
rect 2973 5321 3007 5355
rect 3007 5321 3016 5355
rect 2964 5312 3016 5321
rect 4436 5312 4488 5364
rect 2504 5244 2556 5296
rect 2872 5219 2924 5228
rect 2872 5185 2881 5219
rect 2881 5185 2915 5219
rect 2915 5185 2924 5219
rect 2872 5176 2924 5185
rect 2688 5108 2740 5160
rect 3608 5176 3660 5228
rect 5540 5312 5592 5364
rect 6092 5312 6144 5364
rect 7472 5312 7524 5364
rect 8484 5312 8536 5364
rect 9220 5312 9272 5364
rect 11336 5355 11388 5364
rect 11336 5321 11345 5355
rect 11345 5321 11379 5355
rect 11379 5321 11388 5355
rect 11336 5312 11388 5321
rect 11520 5312 11572 5364
rect 12532 5312 12584 5364
rect 6000 5244 6052 5296
rect 9312 5244 9364 5296
rect 13452 5312 13504 5364
rect 13268 5244 13320 5296
rect 5908 5219 5960 5228
rect 3884 5108 3936 5160
rect 5908 5185 5917 5219
rect 5917 5185 5951 5219
rect 5951 5185 5960 5219
rect 5908 5176 5960 5185
rect 8852 5176 8904 5228
rect 9036 5176 9088 5228
rect 5448 5151 5500 5160
rect 5448 5117 5457 5151
rect 5457 5117 5491 5151
rect 5491 5117 5500 5151
rect 5448 5108 5500 5117
rect 8208 5108 8260 5160
rect 8576 5108 8628 5160
rect 9220 5040 9272 5092
rect 10784 5219 10836 5228
rect 10784 5185 10802 5219
rect 10802 5185 10836 5219
rect 10784 5176 10836 5185
rect 11428 5176 11480 5228
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 14464 5219 14516 5228
rect 14464 5185 14473 5219
rect 14473 5185 14507 5219
rect 14507 5185 14516 5219
rect 14464 5176 14516 5185
rect 17960 5312 18012 5364
rect 16120 5244 16172 5296
rect 16212 5244 16264 5296
rect 15016 5108 15068 5160
rect 15384 5108 15436 5160
rect 17408 5176 17460 5228
rect 16948 5108 17000 5160
rect 4068 4972 4120 5024
rect 8392 4972 8444 5024
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 14372 4972 14424 5024
rect 15200 4972 15252 5024
rect 15292 4972 15344 5024
rect 16580 5040 16632 5092
rect 3110 4870 3162 4922
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 3302 4870 3354 4922
rect 3366 4870 3418 4922
rect 6210 4870 6262 4922
rect 6274 4870 6326 4922
rect 6338 4870 6390 4922
rect 6402 4870 6454 4922
rect 6466 4870 6518 4922
rect 9310 4870 9362 4922
rect 9374 4870 9426 4922
rect 9438 4870 9490 4922
rect 9502 4870 9554 4922
rect 9566 4870 9618 4922
rect 12410 4870 12462 4922
rect 12474 4870 12526 4922
rect 12538 4870 12590 4922
rect 12602 4870 12654 4922
rect 12666 4870 12718 4922
rect 15510 4870 15562 4922
rect 15574 4870 15626 4922
rect 15638 4870 15690 4922
rect 15702 4870 15754 4922
rect 15766 4870 15818 4922
rect 5540 4768 5592 4820
rect 8208 4811 8260 4820
rect 3976 4632 4028 4684
rect 1124 4564 1176 4616
rect 1308 4607 1360 4616
rect 1308 4573 1317 4607
rect 1317 4573 1351 4607
rect 1351 4573 1360 4607
rect 1308 4564 1360 4573
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4068 4564 4120 4573
rect 5816 4700 5868 4752
rect 5632 4675 5684 4684
rect 5632 4641 5641 4675
rect 5641 4641 5675 4675
rect 5675 4641 5684 4675
rect 5632 4632 5684 4641
rect 6092 4675 6144 4684
rect 6092 4641 6101 4675
rect 6101 4641 6135 4675
rect 6135 4641 6144 4675
rect 6092 4632 6144 4641
rect 8208 4777 8217 4811
rect 8217 4777 8251 4811
rect 8251 4777 8260 4811
rect 8208 4768 8260 4777
rect 8852 4768 8904 4820
rect 9128 4632 9180 4684
rect 9220 4675 9272 4684
rect 9220 4641 9229 4675
rect 9229 4641 9263 4675
rect 9263 4641 9272 4675
rect 9220 4632 9272 4641
rect 1860 4496 1912 4548
rect 3516 4496 3568 4548
rect 4988 4496 5040 4548
rect 8208 4607 8260 4616
rect 5448 4496 5500 4548
rect 3056 4471 3108 4480
rect 3056 4437 3065 4471
rect 3065 4437 3099 4471
rect 3099 4437 3108 4471
rect 3056 4428 3108 4437
rect 3700 4471 3752 4480
rect 3700 4437 3709 4471
rect 3709 4437 3743 4471
rect 3743 4437 3752 4471
rect 3700 4428 3752 4437
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 11336 4675 11388 4684
rect 11336 4641 11345 4675
rect 11345 4641 11379 4675
rect 11379 4641 11388 4675
rect 11336 4632 11388 4641
rect 11520 4675 11572 4684
rect 11520 4641 11529 4675
rect 11529 4641 11563 4675
rect 11563 4641 11572 4675
rect 11520 4632 11572 4641
rect 13084 4632 13136 4684
rect 16580 4632 16632 4684
rect 17500 4675 17552 4684
rect 17500 4641 17509 4675
rect 17509 4641 17543 4675
rect 17543 4641 17552 4675
rect 17500 4632 17552 4641
rect 13268 4564 13320 4616
rect 15016 4564 15068 4616
rect 15844 4564 15896 4616
rect 7012 4496 7064 4548
rect 8944 4496 8996 4548
rect 7380 4428 7432 4480
rect 9128 4428 9180 4480
rect 13728 4539 13780 4548
rect 10784 4428 10836 4480
rect 13728 4505 13737 4539
rect 13737 4505 13771 4539
rect 13771 4505 13780 4539
rect 13728 4496 13780 4505
rect 12440 4428 12492 4480
rect 13452 4428 13504 4480
rect 15384 4496 15436 4548
rect 15200 4428 15252 4480
rect 16120 4428 16172 4480
rect 17776 4428 17828 4480
rect 4660 4326 4712 4378
rect 4724 4326 4776 4378
rect 4788 4326 4840 4378
rect 4852 4326 4904 4378
rect 4916 4326 4968 4378
rect 7760 4326 7812 4378
rect 7824 4326 7876 4378
rect 7888 4326 7940 4378
rect 7952 4326 8004 4378
rect 8016 4326 8068 4378
rect 10860 4326 10912 4378
rect 10924 4326 10976 4378
rect 10988 4326 11040 4378
rect 11052 4326 11104 4378
rect 11116 4326 11168 4378
rect 13960 4326 14012 4378
rect 14024 4326 14076 4378
rect 14088 4326 14140 4378
rect 14152 4326 14204 4378
rect 14216 4326 14268 4378
rect 17060 4326 17112 4378
rect 17124 4326 17176 4378
rect 17188 4326 17240 4378
rect 17252 4326 17304 4378
rect 17316 4326 17368 4378
rect 3700 4224 3752 4276
rect 5632 4267 5684 4276
rect 5632 4233 5641 4267
rect 5641 4233 5675 4267
rect 5675 4233 5684 4267
rect 5632 4224 5684 4233
rect 7012 4224 7064 4276
rect 8208 4224 8260 4276
rect 13728 4224 13780 4276
rect 17960 4267 18012 4276
rect 17960 4233 17969 4267
rect 17969 4233 18003 4267
rect 18003 4233 18012 4267
rect 17960 4224 18012 4233
rect 1860 4156 1912 4208
rect 3056 4199 3108 4208
rect 3056 4165 3065 4199
rect 3065 4165 3099 4199
rect 3099 4165 3108 4199
rect 3056 4156 3108 4165
rect 3608 4156 3660 4208
rect 4988 4156 5040 4208
rect 848 4063 900 4072
rect 848 4029 857 4063
rect 857 4029 891 4063
rect 891 4029 900 4063
rect 848 4020 900 4029
rect 3792 4131 3844 4140
rect 1308 4020 1360 4072
rect 3792 4097 3801 4131
rect 3801 4097 3835 4131
rect 3835 4097 3844 4131
rect 3792 4088 3844 4097
rect 3884 4131 3936 4140
rect 3884 4097 3893 4131
rect 3893 4097 3927 4131
rect 3927 4097 3936 4131
rect 3884 4088 3936 4097
rect 5540 4088 5592 4140
rect 7380 4088 7432 4140
rect 8208 4088 8260 4140
rect 11796 4156 11848 4208
rect 12256 4156 12308 4208
rect 13452 4156 13504 4208
rect 13820 4156 13872 4208
rect 8852 4131 8904 4140
rect 8852 4097 8861 4131
rect 8861 4097 8895 4131
rect 8895 4097 8904 4131
rect 8852 4088 8904 4097
rect 10784 4088 10836 4140
rect 11244 4131 11296 4140
rect 11244 4097 11253 4131
rect 11253 4097 11287 4131
rect 11287 4097 11296 4131
rect 11244 4088 11296 4097
rect 12440 4088 12492 4140
rect 16120 4156 16172 4208
rect 1124 3884 1176 3936
rect 4896 4020 4948 4072
rect 5356 4020 5408 4072
rect 8944 4063 8996 4072
rect 8944 4029 8953 4063
rect 8953 4029 8987 4063
rect 8987 4029 8996 4063
rect 8944 4020 8996 4029
rect 11336 4063 11388 4072
rect 11336 4029 11345 4063
rect 11345 4029 11379 4063
rect 11379 4029 11388 4063
rect 11336 4020 11388 4029
rect 13176 4020 13228 4072
rect 13820 4020 13872 4072
rect 14556 4088 14608 4140
rect 15292 4088 15344 4140
rect 2688 3884 2740 3936
rect 3884 3884 3936 3936
rect 4068 3884 4120 3936
rect 6828 3884 6880 3936
rect 11704 3884 11756 3936
rect 12900 3952 12952 4004
rect 15016 4020 15068 4072
rect 15200 4063 15252 4072
rect 15200 4029 15209 4063
rect 15209 4029 15243 4063
rect 15243 4029 15252 4063
rect 15200 4020 15252 4029
rect 15936 4020 15988 4072
rect 16580 4088 16632 4140
rect 18328 4088 18380 4140
rect 16396 4020 16448 4072
rect 14740 3884 14792 3936
rect 18052 3952 18104 4004
rect 3110 3782 3162 3834
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 3302 3782 3354 3834
rect 3366 3782 3418 3834
rect 6210 3782 6262 3834
rect 6274 3782 6326 3834
rect 6338 3782 6390 3834
rect 6402 3782 6454 3834
rect 6466 3782 6518 3834
rect 9310 3782 9362 3834
rect 9374 3782 9426 3834
rect 9438 3782 9490 3834
rect 9502 3782 9554 3834
rect 9566 3782 9618 3834
rect 12410 3782 12462 3834
rect 12474 3782 12526 3834
rect 12538 3782 12590 3834
rect 12602 3782 12654 3834
rect 12666 3782 12718 3834
rect 15510 3782 15562 3834
rect 15574 3782 15626 3834
rect 15638 3782 15690 3834
rect 15702 3782 15754 3834
rect 15766 3782 15818 3834
rect 848 3680 900 3732
rect 3792 3680 3844 3732
rect 11152 3680 11204 3732
rect 11244 3680 11296 3732
rect 12256 3680 12308 3732
rect 4528 3612 4580 3664
rect 2872 3544 2924 3596
rect 2688 3476 2740 3528
rect 3976 3544 4028 3596
rect 8208 3612 8260 3664
rect 15200 3680 15252 3732
rect 4068 3519 4120 3528
rect 2596 3340 2648 3392
rect 2688 3340 2740 3392
rect 4068 3485 4077 3519
rect 4077 3485 4111 3519
rect 4111 3485 4120 3519
rect 4068 3476 4120 3485
rect 6644 3544 6696 3596
rect 7012 3544 7064 3596
rect 11796 3544 11848 3596
rect 13268 3587 13320 3596
rect 4896 3519 4948 3528
rect 4896 3485 4905 3519
rect 4905 3485 4939 3519
rect 4939 3485 4948 3519
rect 4896 3476 4948 3485
rect 5264 3519 5316 3528
rect 5264 3485 5273 3519
rect 5273 3485 5307 3519
rect 5307 3485 5316 3519
rect 5264 3476 5316 3485
rect 5816 3476 5868 3528
rect 6828 3519 6880 3528
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 8392 3476 8444 3528
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 10048 3476 10100 3528
rect 13268 3553 13277 3587
rect 13277 3553 13311 3587
rect 13311 3553 13320 3587
rect 13268 3544 13320 3553
rect 14740 3587 14792 3596
rect 14740 3553 14749 3587
rect 14749 3553 14783 3587
rect 14783 3553 14792 3587
rect 14740 3544 14792 3553
rect 12900 3519 12952 3528
rect 12900 3485 12909 3519
rect 12909 3485 12943 3519
rect 12943 3485 12952 3519
rect 12900 3476 12952 3485
rect 4436 3408 4488 3460
rect 7012 3408 7064 3460
rect 7564 3408 7616 3460
rect 6552 3340 6604 3392
rect 6736 3383 6788 3392
rect 6736 3349 6745 3383
rect 6745 3349 6779 3383
rect 6779 3349 6788 3383
rect 6736 3340 6788 3349
rect 8116 3408 8168 3460
rect 9220 3408 9272 3460
rect 11704 3340 11756 3392
rect 12072 3340 12124 3392
rect 13820 3340 13872 3392
rect 14924 3476 14976 3528
rect 15844 3519 15896 3528
rect 15844 3485 15853 3519
rect 15853 3485 15887 3519
rect 15887 3485 15896 3519
rect 15844 3476 15896 3485
rect 18512 3519 18564 3528
rect 18512 3485 18521 3519
rect 18521 3485 18555 3519
rect 18555 3485 18564 3519
rect 18512 3476 18564 3485
rect 16120 3451 16172 3460
rect 14648 3383 14700 3392
rect 14648 3349 14657 3383
rect 14657 3349 14691 3383
rect 14691 3349 14700 3383
rect 14648 3340 14700 3349
rect 14740 3340 14792 3392
rect 15844 3340 15896 3392
rect 16120 3417 16129 3451
rect 16129 3417 16163 3451
rect 16163 3417 16172 3451
rect 16120 3408 16172 3417
rect 16396 3408 16448 3460
rect 17408 3408 17460 3460
rect 16856 3340 16908 3392
rect 4660 3238 4712 3290
rect 4724 3238 4776 3290
rect 4788 3238 4840 3290
rect 4852 3238 4904 3290
rect 4916 3238 4968 3290
rect 7760 3238 7812 3290
rect 7824 3238 7876 3290
rect 7888 3238 7940 3290
rect 7952 3238 8004 3290
rect 8016 3238 8068 3290
rect 10860 3238 10912 3290
rect 10924 3238 10976 3290
rect 10988 3238 11040 3290
rect 11052 3238 11104 3290
rect 11116 3238 11168 3290
rect 13960 3238 14012 3290
rect 14024 3238 14076 3290
rect 14088 3238 14140 3290
rect 14152 3238 14204 3290
rect 14216 3238 14268 3290
rect 17060 3238 17112 3290
rect 17124 3238 17176 3290
rect 17188 3238 17240 3290
rect 17252 3238 17304 3290
rect 17316 3238 17368 3290
rect 1308 3136 1360 3188
rect 1860 3068 1912 3120
rect 2688 3068 2740 3120
rect 572 2975 624 2984
rect 572 2941 581 2975
rect 581 2941 615 2975
rect 615 2941 624 2975
rect 572 2932 624 2941
rect 2044 2975 2096 2984
rect 2044 2941 2053 2975
rect 2053 2941 2087 2975
rect 2087 2941 2096 2975
rect 6092 3136 6144 3188
rect 8116 3136 8168 3188
rect 8392 3136 8444 3188
rect 7012 3068 7064 3120
rect 3700 3043 3752 3052
rect 3700 3009 3709 3043
rect 3709 3009 3743 3043
rect 3743 3009 3752 3043
rect 3700 3000 3752 3009
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 4344 3043 4396 3052
rect 4344 3009 4353 3043
rect 4353 3009 4387 3043
rect 4387 3009 4396 3043
rect 4344 3000 4396 3009
rect 4528 3000 4580 3052
rect 5172 3043 5224 3052
rect 2044 2932 2096 2941
rect 940 2796 992 2848
rect 3608 2932 3660 2984
rect 3976 2975 4028 2984
rect 3976 2941 3985 2975
rect 3985 2941 4019 2975
rect 4019 2941 4028 2975
rect 3976 2932 4028 2941
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 7564 3043 7616 3052
rect 2596 2796 2648 2848
rect 4528 2839 4580 2848
rect 4528 2805 4537 2839
rect 4537 2805 4571 2839
rect 4571 2805 4580 2839
rect 4528 2796 4580 2805
rect 5080 2839 5132 2848
rect 5080 2805 5089 2839
rect 5089 2805 5123 2839
rect 5123 2805 5132 2839
rect 5080 2796 5132 2805
rect 6092 2932 6144 2984
rect 6920 2975 6972 2984
rect 6920 2941 6929 2975
rect 6929 2941 6963 2975
rect 6963 2941 6972 2975
rect 7564 3009 7573 3043
rect 7573 3009 7607 3043
rect 7607 3009 7616 3043
rect 7564 3000 7616 3009
rect 8024 3043 8076 3052
rect 8024 3009 8033 3043
rect 8033 3009 8067 3043
rect 8067 3009 8076 3043
rect 8024 3000 8076 3009
rect 8668 3000 8720 3052
rect 6920 2932 6972 2941
rect 8944 3043 8996 3052
rect 8944 3009 8953 3043
rect 8953 3009 8987 3043
rect 8987 3009 8996 3043
rect 8944 3000 8996 3009
rect 10048 3000 10100 3052
rect 12072 3043 12124 3052
rect 12072 3009 12081 3043
rect 12081 3009 12115 3043
rect 12115 3009 12124 3043
rect 12072 3000 12124 3009
rect 13452 3068 13504 3120
rect 12532 3000 12584 3052
rect 12808 2932 12860 2984
rect 12992 2932 13044 2984
rect 13820 3000 13872 3052
rect 14648 3043 14700 3052
rect 14648 3009 14657 3043
rect 14657 3009 14691 3043
rect 14691 3009 14700 3043
rect 14648 3000 14700 3009
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 15016 3136 15068 3188
rect 16120 3136 16172 3188
rect 15844 3068 15896 3120
rect 16856 3000 16908 3052
rect 17776 3043 17828 3052
rect 17776 3009 17785 3043
rect 17785 3009 17819 3043
rect 17819 3009 17828 3043
rect 17776 3000 17828 3009
rect 14740 2932 14792 2984
rect 17684 2932 17736 2984
rect 6828 2864 6880 2916
rect 8668 2864 8720 2916
rect 8944 2864 8996 2916
rect 16396 2864 16448 2916
rect 18144 2864 18196 2916
rect 7196 2796 7248 2848
rect 11796 2796 11848 2848
rect 11980 2796 12032 2848
rect 14372 2796 14424 2848
rect 17132 2839 17184 2848
rect 17132 2805 17141 2839
rect 17141 2805 17175 2839
rect 17175 2805 17184 2839
rect 17132 2796 17184 2805
rect 17868 2796 17920 2848
rect 3110 2694 3162 2746
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 3302 2694 3354 2746
rect 3366 2694 3418 2746
rect 6210 2694 6262 2746
rect 6274 2694 6326 2746
rect 6338 2694 6390 2746
rect 6402 2694 6454 2746
rect 6466 2694 6518 2746
rect 9310 2694 9362 2746
rect 9374 2694 9426 2746
rect 9438 2694 9490 2746
rect 9502 2694 9554 2746
rect 9566 2694 9618 2746
rect 12410 2694 12462 2746
rect 12474 2694 12526 2746
rect 12538 2694 12590 2746
rect 12602 2694 12654 2746
rect 12666 2694 12718 2746
rect 15510 2694 15562 2746
rect 15574 2694 15626 2746
rect 15638 2694 15690 2746
rect 15702 2694 15754 2746
rect 15766 2694 15818 2746
rect 572 2592 624 2644
rect 3700 2592 3752 2644
rect 3884 2592 3936 2644
rect 4528 2592 4580 2644
rect 4712 2592 4764 2644
rect 5356 2592 5408 2644
rect 6092 2635 6144 2644
rect 6092 2601 6101 2635
rect 6101 2601 6135 2635
rect 6135 2601 6144 2635
rect 6092 2592 6144 2601
rect 6736 2592 6788 2644
rect 3516 2524 3568 2576
rect 8852 2592 8904 2644
rect 10048 2592 10100 2644
rect 11336 2592 11388 2644
rect 12808 2592 12860 2644
rect 12992 2592 13044 2644
rect 15108 2592 15160 2644
rect 17132 2592 17184 2644
rect 17684 2635 17736 2644
rect 2228 2456 2280 2508
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 2780 2456 2832 2465
rect 4344 2456 4396 2508
rect 7656 2524 7708 2576
rect 8024 2524 8076 2576
rect 940 2431 992 2440
rect 940 2397 949 2431
rect 949 2397 983 2431
rect 983 2397 992 2431
rect 940 2388 992 2397
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 2872 2388 2924 2440
rect 3516 2431 3568 2440
rect 3516 2397 3525 2431
rect 3525 2397 3559 2431
rect 3559 2397 3568 2431
rect 3516 2388 3568 2397
rect 4528 2431 4580 2440
rect 2964 2320 3016 2372
rect 4528 2397 4537 2431
rect 4537 2397 4571 2431
rect 4571 2397 4580 2431
rect 4528 2388 4580 2397
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 6552 2456 6604 2508
rect 6828 2456 6880 2508
rect 4620 2320 4672 2372
rect 6000 2388 6052 2440
rect 7196 2388 7248 2440
rect 9036 2456 9088 2508
rect 9220 2456 9272 2508
rect 13176 2524 13228 2576
rect 17684 2601 17693 2635
rect 17693 2601 17727 2635
rect 17727 2601 17736 2635
rect 17684 2592 17736 2601
rect 8116 2388 8168 2440
rect 8668 2431 8720 2440
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 9496 2388 9548 2440
rect 3424 2252 3476 2304
rect 4344 2252 4396 2304
rect 4436 2252 4488 2304
rect 9312 2320 9364 2372
rect 11244 2388 11296 2440
rect 13268 2456 13320 2508
rect 13728 2456 13780 2508
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 15108 2388 15160 2440
rect 17776 2524 17828 2576
rect 17132 2431 17184 2440
rect 17132 2397 17141 2431
rect 17141 2397 17175 2431
rect 17175 2397 17184 2431
rect 17132 2388 17184 2397
rect 17868 2431 17920 2440
rect 17868 2397 17877 2431
rect 17877 2397 17911 2431
rect 17911 2397 17920 2431
rect 17868 2388 17920 2397
rect 18144 2431 18196 2440
rect 18144 2397 18153 2431
rect 18153 2397 18187 2431
rect 18187 2397 18196 2431
rect 18144 2388 18196 2397
rect 5264 2252 5316 2304
rect 5448 2295 5500 2304
rect 5448 2261 5457 2295
rect 5457 2261 5491 2295
rect 5491 2261 5500 2295
rect 5448 2252 5500 2261
rect 7012 2252 7064 2304
rect 9220 2252 9272 2304
rect 11336 2363 11388 2372
rect 11336 2329 11345 2363
rect 11345 2329 11379 2363
rect 11379 2329 11388 2363
rect 11336 2320 11388 2329
rect 11612 2320 11664 2372
rect 11704 2363 11756 2372
rect 11704 2329 11713 2363
rect 11713 2329 11747 2363
rect 11747 2329 11756 2363
rect 11704 2320 11756 2329
rect 13820 2320 13872 2372
rect 15476 2363 15528 2372
rect 15476 2329 15485 2363
rect 15485 2329 15519 2363
rect 15519 2329 15528 2363
rect 15476 2320 15528 2329
rect 18236 2320 18288 2372
rect 11428 2252 11480 2304
rect 14464 2252 14516 2304
rect 4660 2150 4712 2202
rect 4724 2150 4776 2202
rect 4788 2150 4840 2202
rect 4852 2150 4904 2202
rect 4916 2150 4968 2202
rect 7760 2150 7812 2202
rect 7824 2150 7876 2202
rect 7888 2150 7940 2202
rect 7952 2150 8004 2202
rect 8016 2150 8068 2202
rect 10860 2150 10912 2202
rect 10924 2150 10976 2202
rect 10988 2150 11040 2202
rect 11052 2150 11104 2202
rect 11116 2150 11168 2202
rect 13960 2150 14012 2202
rect 14024 2150 14076 2202
rect 14088 2150 14140 2202
rect 14152 2150 14204 2202
rect 14216 2150 14268 2202
rect 17060 2150 17112 2202
rect 17124 2150 17176 2202
rect 17188 2150 17240 2202
rect 17252 2150 17304 2202
rect 17316 2150 17368 2202
rect 2228 2091 2280 2100
rect 2228 2057 2237 2091
rect 2237 2057 2271 2091
rect 2271 2057 2280 2091
rect 2228 2048 2280 2057
rect 2872 2091 2924 2100
rect 2872 2057 2881 2091
rect 2881 2057 2915 2091
rect 2915 2057 2924 2091
rect 2872 2048 2924 2057
rect 3424 2048 3476 2100
rect 7104 2048 7156 2100
rect 8208 2048 8260 2100
rect 8668 2048 8720 2100
rect 9312 2048 9364 2100
rect 11244 2048 11296 2100
rect 11612 2091 11664 2100
rect 11612 2057 11621 2091
rect 11621 2057 11655 2091
rect 11655 2057 11664 2091
rect 11612 2048 11664 2057
rect 13176 2091 13228 2100
rect 13176 2057 13185 2091
rect 13185 2057 13219 2091
rect 13219 2057 13228 2091
rect 13820 2091 13872 2100
rect 13176 2048 13228 2057
rect 4528 1980 4580 2032
rect 2780 1912 2832 1964
rect 4160 1955 4212 1964
rect 4160 1921 4169 1955
rect 4169 1921 4203 1955
rect 4203 1921 4212 1955
rect 4160 1912 4212 1921
rect 4344 1955 4396 1964
rect 4344 1921 4353 1955
rect 4353 1921 4387 1955
rect 4387 1921 4396 1955
rect 4344 1912 4396 1921
rect 4436 1912 4488 1964
rect 5080 1955 5132 1964
rect 5080 1921 5089 1955
rect 5089 1921 5123 1955
rect 5123 1921 5132 1955
rect 5080 1912 5132 1921
rect 5448 1955 5500 1964
rect 5448 1921 5457 1955
rect 5457 1921 5491 1955
rect 5491 1921 5500 1955
rect 5448 1912 5500 1921
rect 6920 1980 6972 2032
rect 7288 1955 7340 1964
rect 7288 1921 7297 1955
rect 7297 1921 7331 1955
rect 7331 1921 7340 1955
rect 7288 1912 7340 1921
rect 2228 1844 2280 1896
rect 2872 1844 2924 1896
rect 3608 1844 3660 1896
rect 3976 1887 4028 1896
rect 3976 1853 3985 1887
rect 3985 1853 4019 1887
rect 4019 1853 4028 1887
rect 3976 1844 4028 1853
rect 5816 1887 5868 1896
rect 5816 1853 5825 1887
rect 5825 1853 5859 1887
rect 5859 1853 5868 1887
rect 5816 1844 5868 1853
rect 5908 1844 5960 1896
rect 7012 1887 7064 1896
rect 7012 1853 7021 1887
rect 7021 1853 7055 1887
rect 7055 1853 7064 1887
rect 7012 1844 7064 1853
rect 3516 1776 3568 1828
rect 6920 1776 6972 1828
rect 7656 1912 7708 1964
rect 7932 1955 7984 1964
rect 7932 1921 7941 1955
rect 7941 1921 7975 1955
rect 7975 1921 7984 1955
rect 7932 1912 7984 1921
rect 8024 1844 8076 1896
rect 7472 1776 7524 1828
rect 8760 1912 8812 1964
rect 9220 1955 9272 1964
rect 9220 1921 9229 1955
rect 9229 1921 9263 1955
rect 9263 1921 9272 1955
rect 9220 1912 9272 1921
rect 9404 1980 9456 2032
rect 10324 1980 10376 2032
rect 9772 1912 9824 1964
rect 10692 1912 10744 1964
rect 11336 1980 11388 2032
rect 12992 1980 13044 2032
rect 13820 2057 13829 2091
rect 13829 2057 13863 2091
rect 13863 2057 13872 2091
rect 13820 2048 13872 2057
rect 14740 2048 14792 2100
rect 15108 2048 15160 2100
rect 17500 2048 17552 2100
rect 18236 2091 18288 2100
rect 18236 2057 18245 2091
rect 18245 2057 18279 2091
rect 18279 2057 18288 2091
rect 18236 2048 18288 2057
rect 9496 1887 9548 1896
rect 9496 1853 9505 1887
rect 9505 1853 9539 1887
rect 9539 1853 9548 1887
rect 11152 1955 11204 1964
rect 11152 1921 11161 1955
rect 11161 1921 11195 1955
rect 11195 1921 11204 1955
rect 11428 1955 11480 1964
rect 11152 1912 11204 1921
rect 11428 1921 11437 1955
rect 11437 1921 11471 1955
rect 11471 1921 11480 1955
rect 11428 1912 11480 1921
rect 11612 1912 11664 1964
rect 12900 1912 12952 1964
rect 13084 1955 13136 1964
rect 13084 1921 13093 1955
rect 13093 1921 13127 1955
rect 13127 1921 13136 1955
rect 13084 1912 13136 1921
rect 11336 1887 11388 1896
rect 9496 1844 9548 1853
rect 8484 1776 8536 1828
rect 9312 1776 9364 1828
rect 10140 1776 10192 1828
rect 11336 1853 11345 1887
rect 11345 1853 11379 1887
rect 11379 1853 11388 1887
rect 15384 1980 15436 2032
rect 11336 1844 11388 1853
rect 13912 1844 13964 1896
rect 14372 1912 14424 1964
rect 14832 1955 14884 1964
rect 14832 1921 14841 1955
rect 14841 1921 14875 1955
rect 14875 1921 14884 1955
rect 14832 1912 14884 1921
rect 14924 1912 14976 1964
rect 17408 1980 17460 2032
rect 16488 1912 16540 1964
rect 14464 1844 14516 1896
rect 848 1751 900 1760
rect 848 1717 857 1751
rect 857 1717 891 1751
rect 891 1717 900 1751
rect 848 1708 900 1717
rect 5356 1708 5408 1760
rect 7012 1708 7064 1760
rect 7288 1751 7340 1760
rect 7288 1717 7297 1751
rect 7297 1717 7331 1751
rect 7331 1717 7340 1751
rect 7288 1708 7340 1717
rect 7840 1751 7892 1760
rect 7840 1717 7849 1751
rect 7849 1717 7883 1751
rect 7883 1717 7892 1751
rect 7840 1708 7892 1717
rect 7932 1708 7984 1760
rect 8760 1708 8812 1760
rect 9864 1708 9916 1760
rect 11060 1708 11112 1760
rect 11336 1708 11388 1760
rect 12808 1708 12860 1760
rect 14188 1708 14240 1760
rect 14740 1708 14792 1760
rect 15476 1844 15528 1896
rect 16120 1844 16172 1896
rect 16672 1751 16724 1760
rect 16672 1717 16681 1751
rect 16681 1717 16715 1751
rect 16715 1717 16724 1751
rect 16672 1708 16724 1717
rect 3110 1606 3162 1658
rect 3174 1606 3226 1658
rect 3238 1606 3290 1658
rect 3302 1606 3354 1658
rect 3366 1606 3418 1658
rect 6210 1606 6262 1658
rect 6274 1606 6326 1658
rect 6338 1606 6390 1658
rect 6402 1606 6454 1658
rect 6466 1606 6518 1658
rect 9310 1606 9362 1658
rect 9374 1606 9426 1658
rect 9438 1606 9490 1658
rect 9502 1606 9554 1658
rect 9566 1606 9618 1658
rect 12410 1606 12462 1658
rect 12474 1606 12526 1658
rect 12538 1606 12590 1658
rect 12602 1606 12654 1658
rect 12666 1606 12718 1658
rect 15510 1606 15562 1658
rect 15574 1606 15626 1658
rect 15638 1606 15690 1658
rect 15702 1606 15754 1658
rect 15766 1606 15818 1658
rect 2780 1504 2832 1556
rect 5908 1547 5960 1556
rect 1308 1343 1360 1352
rect 1308 1309 1317 1343
rect 1317 1309 1351 1343
rect 1351 1309 1360 1343
rect 1308 1300 1360 1309
rect 5908 1513 5917 1547
rect 5917 1513 5951 1547
rect 5951 1513 5960 1547
rect 5908 1504 5960 1513
rect 6644 1504 6696 1556
rect 6920 1504 6972 1556
rect 9680 1504 9732 1556
rect 10048 1547 10100 1556
rect 10048 1513 10057 1547
rect 10057 1513 10091 1547
rect 10091 1513 10100 1547
rect 10048 1504 10100 1513
rect 5264 1368 5316 1420
rect 3608 1300 3660 1352
rect 5540 1300 5592 1352
rect 6000 1368 6052 1420
rect 7196 1436 7248 1488
rect 6644 1368 6696 1420
rect 7380 1411 7432 1420
rect 7380 1377 7389 1411
rect 7389 1377 7423 1411
rect 7423 1377 7432 1411
rect 7380 1368 7432 1377
rect 7840 1368 7892 1420
rect 8116 1436 8168 1488
rect 11060 1504 11112 1556
rect 11152 1504 11204 1556
rect 9772 1368 9824 1420
rect 10784 1436 10836 1488
rect 11612 1436 11664 1488
rect 11796 1436 11848 1488
rect 1584 1275 1636 1284
rect 1584 1241 1593 1275
rect 1593 1241 1627 1275
rect 1627 1241 1636 1275
rect 1584 1232 1636 1241
rect 3424 1275 3476 1284
rect 388 1164 440 1216
rect 2596 1164 2648 1216
rect 3424 1241 3433 1275
rect 3433 1241 3467 1275
rect 3467 1241 3476 1275
rect 3424 1232 3476 1241
rect 3976 1232 4028 1284
rect 6552 1300 6604 1352
rect 6368 1232 6420 1284
rect 3884 1164 3936 1216
rect 6092 1207 6144 1216
rect 6092 1173 6101 1207
rect 6101 1173 6135 1207
rect 6135 1173 6144 1207
rect 6092 1164 6144 1173
rect 7104 1300 7156 1352
rect 7472 1300 7524 1352
rect 7196 1232 7248 1284
rect 7380 1232 7432 1284
rect 8116 1343 8168 1352
rect 8116 1309 8125 1343
rect 8125 1309 8159 1343
rect 8159 1309 8168 1343
rect 8116 1300 8168 1309
rect 8852 1300 8904 1352
rect 9864 1343 9916 1352
rect 9864 1309 9873 1343
rect 9873 1309 9907 1343
rect 9907 1309 9916 1343
rect 9864 1300 9916 1309
rect 6920 1207 6972 1216
rect 6920 1173 6929 1207
rect 6929 1173 6963 1207
rect 6963 1173 6972 1207
rect 6920 1164 6972 1173
rect 7012 1164 7064 1216
rect 8208 1164 8260 1216
rect 9680 1232 9732 1284
rect 10140 1343 10192 1352
rect 10140 1309 10149 1343
rect 10149 1309 10183 1343
rect 10183 1309 10192 1343
rect 10140 1300 10192 1309
rect 10324 1343 10376 1352
rect 10324 1309 10333 1343
rect 10333 1309 10367 1343
rect 10367 1309 10376 1343
rect 10324 1300 10376 1309
rect 11336 1368 11388 1420
rect 14648 1504 14700 1556
rect 14832 1504 14884 1556
rect 14188 1436 14240 1488
rect 14280 1436 14332 1488
rect 8576 1164 8628 1216
rect 12072 1232 12124 1284
rect 11244 1207 11296 1216
rect 11244 1173 11253 1207
rect 11253 1173 11287 1207
rect 11287 1173 11296 1207
rect 11244 1164 11296 1173
rect 12256 1300 12308 1352
rect 12808 1232 12860 1284
rect 13176 1232 13228 1284
rect 13544 1300 13596 1352
rect 14096 1300 14148 1352
rect 15108 1368 15160 1420
rect 15660 1368 15712 1420
rect 16120 1343 16172 1352
rect 13728 1232 13780 1284
rect 16120 1309 16129 1343
rect 16129 1309 16163 1343
rect 16163 1309 16172 1343
rect 16120 1300 16172 1309
rect 16396 1275 16448 1284
rect 16396 1241 16405 1275
rect 16405 1241 16439 1275
rect 16439 1241 16448 1275
rect 16396 1232 16448 1241
rect 12624 1207 12676 1216
rect 12624 1173 12633 1207
rect 12633 1173 12667 1207
rect 12667 1173 12676 1207
rect 12624 1164 12676 1173
rect 12900 1164 12952 1216
rect 13820 1164 13872 1216
rect 14464 1164 14516 1216
rect 15016 1164 15068 1216
rect 15844 1164 15896 1216
rect 17868 1207 17920 1216
rect 17868 1173 17877 1207
rect 17877 1173 17911 1207
rect 17911 1173 17920 1207
rect 17868 1164 17920 1173
rect 4660 1062 4712 1114
rect 4724 1062 4776 1114
rect 4788 1062 4840 1114
rect 4852 1062 4904 1114
rect 4916 1062 4968 1114
rect 7760 1062 7812 1114
rect 7824 1062 7876 1114
rect 7888 1062 7940 1114
rect 7952 1062 8004 1114
rect 8016 1062 8068 1114
rect 10860 1062 10912 1114
rect 10924 1062 10976 1114
rect 10988 1062 11040 1114
rect 11052 1062 11104 1114
rect 11116 1062 11168 1114
rect 13960 1062 14012 1114
rect 14024 1062 14076 1114
rect 14088 1062 14140 1114
rect 14152 1062 14204 1114
rect 14216 1062 14268 1114
rect 17060 1062 17112 1114
rect 17124 1062 17176 1114
rect 17188 1062 17240 1114
rect 17252 1062 17304 1114
rect 17316 1062 17368 1114
rect 2780 960 2832 1012
rect 3424 960 3476 1012
rect 5816 960 5868 1012
rect 388 867 440 876
rect 388 833 397 867
rect 397 833 431 867
rect 431 833 440 867
rect 388 824 440 833
rect 848 824 900 876
rect 2228 892 2280 944
rect 9128 960 9180 1012
rect 9312 960 9364 1012
rect 2596 824 2648 876
rect 5172 824 5224 876
rect 3608 756 3660 808
rect 3792 799 3844 808
rect 3792 765 3801 799
rect 3801 765 3835 799
rect 3835 765 3844 799
rect 3792 756 3844 765
rect 3976 799 4028 808
rect 3976 765 3985 799
rect 3985 765 4019 799
rect 4019 765 4028 799
rect 3976 756 4028 765
rect 5264 799 5316 808
rect 5264 765 5273 799
rect 5273 765 5307 799
rect 5307 765 5316 799
rect 5264 756 5316 765
rect 1308 620 1360 672
rect 3884 620 3936 672
rect 8392 892 8444 944
rect 8852 935 8904 944
rect 8852 901 8861 935
rect 8861 901 8895 935
rect 8895 901 8904 935
rect 8852 892 8904 901
rect 13728 960 13780 1012
rect 12164 935 12216 944
rect 7012 867 7064 876
rect 7012 833 7021 867
rect 7021 833 7055 867
rect 7055 833 7064 867
rect 7012 824 7064 833
rect 7380 799 7432 808
rect 7380 765 7389 799
rect 7389 765 7423 799
rect 7423 765 7432 799
rect 7380 756 7432 765
rect 8760 756 8812 808
rect 9312 756 9364 808
rect 12164 901 12173 935
rect 12173 901 12207 935
rect 12207 901 12216 935
rect 12164 892 12216 901
rect 12900 935 12952 944
rect 12900 901 12909 935
rect 12909 901 12943 935
rect 12943 901 12952 935
rect 12900 892 12952 901
rect 10600 756 10652 808
rect 6368 688 6420 740
rect 7472 688 7524 740
rect 12348 824 12400 876
rect 12808 867 12860 876
rect 12808 833 12817 867
rect 12817 833 12851 867
rect 12851 833 12860 867
rect 13176 867 13228 876
rect 12808 824 12860 833
rect 13176 833 13185 867
rect 13185 833 13219 867
rect 13219 833 13228 867
rect 13176 824 13228 833
rect 13820 892 13872 944
rect 14372 960 14424 1012
rect 16396 1003 16448 1012
rect 14464 867 14516 876
rect 11796 688 11848 740
rect 8852 620 8904 672
rect 11612 663 11664 672
rect 11612 629 11621 663
rect 11621 629 11655 663
rect 11655 629 11664 663
rect 11612 620 11664 629
rect 11704 620 11756 672
rect 14464 833 14473 867
rect 14473 833 14507 867
rect 14507 833 14516 867
rect 14464 824 14516 833
rect 15844 892 15896 944
rect 15200 756 15252 808
rect 16396 969 16405 1003
rect 16405 969 16439 1003
rect 16439 969 16448 1003
rect 16396 960 16448 969
rect 16488 960 16540 1012
rect 17408 960 17460 1012
rect 16580 867 16632 876
rect 16580 833 16589 867
rect 16589 833 16623 867
rect 16623 833 16632 867
rect 16580 824 16632 833
rect 17224 867 17276 876
rect 17224 833 17233 867
rect 17233 833 17267 867
rect 17267 833 17276 867
rect 17224 824 17276 833
rect 18328 824 18380 876
rect 16948 756 17000 808
rect 18512 799 18564 808
rect 15660 688 15712 740
rect 18512 765 18521 799
rect 18521 765 18555 799
rect 18555 765 18564 799
rect 18512 756 18564 765
rect 14740 620 14792 672
rect 3110 518 3162 570
rect 3174 518 3226 570
rect 3238 518 3290 570
rect 3302 518 3354 570
rect 3366 518 3418 570
rect 6210 518 6262 570
rect 6274 518 6326 570
rect 6338 518 6390 570
rect 6402 518 6454 570
rect 6466 518 6518 570
rect 9310 518 9362 570
rect 9374 518 9426 570
rect 9438 518 9490 570
rect 9502 518 9554 570
rect 9566 518 9618 570
rect 12410 518 12462 570
rect 12474 518 12526 570
rect 12538 518 12590 570
rect 12602 518 12654 570
rect 12666 518 12718 570
rect 15510 518 15562 570
rect 15574 518 15626 570
rect 15638 518 15690 570
rect 15702 518 15754 570
rect 15766 518 15818 570
rect 1584 416 1636 468
rect 2596 459 2648 468
rect 2596 425 2605 459
rect 2605 425 2639 459
rect 2639 425 2648 459
rect 2596 416 2648 425
rect 3792 416 3844 468
rect 5264 416 5316 468
rect 6552 416 6604 468
rect 3516 280 3568 332
rect 5540 348 5592 400
rect 6092 280 6144 332
rect 7104 416 7156 468
rect 8392 416 8444 468
rect 8576 416 8628 468
rect 10600 459 10652 468
rect 10600 425 10609 459
rect 10609 425 10643 459
rect 10643 425 10652 459
rect 10600 416 10652 425
rect 13084 416 13136 468
rect 15016 459 15068 468
rect 15016 425 15025 459
rect 15025 425 15059 459
rect 15059 425 15068 459
rect 15016 416 15068 425
rect 16948 459 17000 468
rect 16948 425 16957 459
rect 16957 425 16991 459
rect 16991 425 17000 459
rect 16948 416 17000 425
rect 17224 459 17276 468
rect 17224 425 17233 459
rect 17233 425 17267 459
rect 17267 425 17276 459
rect 17224 416 17276 425
rect 18512 459 18564 468
rect 18512 425 18521 459
rect 18521 425 18555 459
rect 18555 425 18564 459
rect 18512 416 18564 425
rect 9036 323 9088 332
rect 9036 289 9045 323
rect 9045 289 9079 323
rect 9079 289 9088 323
rect 9036 280 9088 289
rect 1308 255 1360 264
rect 1308 221 1317 255
rect 1317 221 1351 255
rect 1351 221 1360 255
rect 1308 212 1360 221
rect 2964 212 3016 264
rect 7288 212 7340 264
rect 8852 255 8904 264
rect 8852 221 8861 255
rect 8861 221 8895 255
rect 8895 221 8904 255
rect 8852 212 8904 221
rect 9864 212 9916 264
rect 11244 280 11296 332
rect 6920 144 6972 196
rect 10784 212 10836 264
rect 11612 212 11664 264
rect 12808 255 12860 264
rect 12808 221 12817 255
rect 12817 221 12851 255
rect 12851 221 12860 255
rect 12808 212 12860 221
rect 13176 280 13228 332
rect 16672 280 16724 332
rect 14740 255 14792 264
rect 14740 221 14749 255
rect 14749 221 14783 255
rect 14783 221 14792 255
rect 14740 212 14792 221
rect 16580 212 16632 264
rect 17868 212 17920 264
rect 11336 144 11388 196
rect 4660 -26 4712 26
rect 4724 -26 4776 26
rect 4788 -26 4840 26
rect 4852 -26 4904 26
rect 4916 -26 4968 26
rect 7760 -26 7812 26
rect 7824 -26 7876 26
rect 7888 -26 7940 26
rect 7952 -26 8004 26
rect 8016 -26 8068 26
rect 10860 -26 10912 26
rect 10924 -26 10976 26
rect 10988 -26 11040 26
rect 11052 -26 11104 26
rect 11116 -26 11168 26
rect 13960 -26 14012 26
rect 14024 -26 14076 26
rect 14088 -26 14140 26
rect 14152 -26 14204 26
rect 14216 -26 14268 26
rect 17060 -26 17112 26
rect 17124 -26 17176 26
rect 17188 -26 17240 26
rect 17252 -26 17304 26
rect 17316 -26 17368 26
<< metal2 >>
rect 1398 11200 1454 12000
rect 4250 11200 4306 12000
rect 7102 11200 7158 12000
rect 9954 11200 10010 12000
rect 12806 11200 12862 12000
rect 15396 11206 15608 11234
rect 296 10056 348 10062
rect 296 9998 348 10004
rect 940 10056 992 10062
rect 940 9998 992 10004
rect 1216 10056 1268 10062
rect 1216 9998 1268 10004
rect 308 8430 336 9998
rect 388 9988 440 9994
rect 388 9930 440 9936
rect 400 9586 428 9930
rect 664 9920 716 9926
rect 664 9862 716 9868
rect 676 9586 704 9862
rect 388 9580 440 9586
rect 388 9522 440 9528
rect 664 9580 716 9586
rect 664 9522 716 9528
rect 952 9178 980 9998
rect 1228 9518 1256 9998
rect 1216 9512 1268 9518
rect 1216 9454 1268 9460
rect 1412 9178 1440 11200
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 2044 10600 2096 10606
rect 2044 10542 2096 10548
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1964 10130 1992 10406
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 1584 9988 1636 9994
rect 1584 9930 1636 9936
rect 1596 9586 1624 9930
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 940 9172 992 9178
rect 940 9114 992 9120
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1412 8974 1440 9114
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 2056 8634 2084 10542
rect 2148 9722 2176 10610
rect 3110 10364 3418 10384
rect 3110 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3276 10364
rect 3332 10362 3356 10364
rect 3412 10362 3418 10364
rect 3172 10310 3174 10362
rect 3354 10310 3356 10362
rect 3110 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3276 10310
rect 3332 10308 3356 10310
rect 3412 10308 3418 10310
rect 3110 10288 3418 10308
rect 3528 10266 3556 10610
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3804 10266 3832 10542
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2240 9382 2268 9590
rect 2608 9586 2636 9862
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2688 9648 2740 9654
rect 2688 9590 2740 9596
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2148 8838 2176 8978
rect 2240 8974 2268 9318
rect 2608 9110 2636 9522
rect 2596 9104 2648 9110
rect 2596 9046 2648 9052
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2136 8832 2188 8838
rect 2136 8774 2188 8780
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2148 8498 2176 8774
rect 2240 8566 2268 8910
rect 2320 8900 2372 8906
rect 2320 8842 2372 8848
rect 2332 8634 2360 8842
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2608 8566 2636 8774
rect 2228 8560 2280 8566
rect 2228 8502 2280 8508
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 296 8424 348 8430
rect 296 8366 348 8372
rect 572 8424 624 8430
rect 572 8366 624 8372
rect 308 6254 336 8366
rect 584 8090 612 8366
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 572 8084 624 8090
rect 572 8026 624 8032
rect 1308 7948 1360 7954
rect 1308 7890 1360 7896
rect 1320 7546 1348 7890
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 1308 7540 1360 7546
rect 1308 7482 1360 7488
rect 1964 7478 1992 7822
rect 1952 7472 2004 7478
rect 1952 7414 2004 7420
rect 2056 7410 2084 8230
rect 2148 8090 2176 8434
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2148 7410 2176 8026
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 572 6656 624 6662
rect 572 6598 624 6604
rect 584 6390 612 6598
rect 2240 6390 2268 8502
rect 2700 8498 2728 9590
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2884 9450 2912 9522
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2780 8900 2832 8906
rect 2780 8842 2832 8848
rect 2792 8566 2820 8842
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2884 8430 2912 9386
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2976 8294 3004 9658
rect 3528 9586 3556 10202
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3110 9276 3418 9296
rect 3110 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3276 9276
rect 3332 9274 3356 9276
rect 3412 9274 3418 9276
rect 3172 9222 3174 9274
rect 3354 9222 3356 9274
rect 3110 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3276 9222
rect 3332 9220 3356 9222
rect 3412 9220 3418 9222
rect 3110 9200 3418 9220
rect 3620 8974 3648 9862
rect 3712 9654 3740 9998
rect 3700 9648 3752 9654
rect 3700 9590 3752 9596
rect 3896 9450 3924 9998
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3700 9036 3752 9042
rect 3700 8978 3752 8984
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3712 8430 3740 8978
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2332 7410 2360 8026
rect 2516 7818 2544 8026
rect 2976 7954 3004 8230
rect 3110 8188 3418 8208
rect 3110 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3276 8188
rect 3332 8186 3356 8188
rect 3412 8186 3418 8188
rect 3172 8134 3174 8186
rect 3354 8134 3356 8186
rect 3110 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3276 8134
rect 3332 8132 3356 8134
rect 3412 8132 3418 8134
rect 3110 8112 3418 8132
rect 3712 8022 3740 8366
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 3700 8016 3752 8022
rect 3700 7958 3752 7964
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 3712 7886 3740 7958
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 2504 7812 2556 7818
rect 2504 7754 2556 7760
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2516 7154 2544 7346
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2424 7126 2544 7154
rect 2424 6798 2452 7126
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2424 6458 2452 6734
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 572 6384 624 6390
rect 572 6326 624 6332
rect 2228 6384 2280 6390
rect 2228 6326 2280 6332
rect 296 6248 348 6254
rect 296 6190 348 6196
rect 308 5778 336 6190
rect 2240 6118 2268 6326
rect 2516 6186 2544 6802
rect 2608 6458 2636 7278
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 296 5772 348 5778
rect 296 5714 348 5720
rect 1216 5636 1268 5642
rect 1216 5578 1268 5584
rect 1228 5370 1256 5578
rect 2240 5574 2268 6054
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 1216 5364 1268 5370
rect 1216 5306 1268 5312
rect 2516 5302 2544 6122
rect 2504 5296 2556 5302
rect 2504 5238 2556 5244
rect 2700 5166 2728 6258
rect 2792 5370 2820 6258
rect 2884 6254 2912 6734
rect 2976 6662 3004 7142
rect 3110 7100 3418 7120
rect 3110 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3276 7100
rect 3332 7098 3356 7100
rect 3412 7098 3418 7100
rect 3172 7046 3174 7098
rect 3354 7046 3356 7098
rect 3110 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3276 7046
rect 3332 7044 3356 7046
rect 3412 7044 3418 7046
rect 3110 7024 3418 7044
rect 3712 6866 3740 7822
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3804 7478 3832 7686
rect 3792 7472 3844 7478
rect 3790 7440 3792 7449
rect 3844 7440 3846 7449
rect 3790 7375 3846 7384
rect 3896 7342 3924 8298
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3896 7002 3924 7278
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3988 6866 4016 9318
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 4080 8362 4108 8842
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4264 8090 4292 11200
rect 4660 10908 4968 10928
rect 4660 10906 4666 10908
rect 4722 10906 4746 10908
rect 4802 10906 4826 10908
rect 4882 10906 4906 10908
rect 4962 10906 4968 10908
rect 4722 10854 4724 10906
rect 4904 10854 4906 10906
rect 4660 10852 4666 10854
rect 4722 10852 4746 10854
rect 4802 10852 4826 10854
rect 4882 10852 4906 10854
rect 4962 10852 4968 10854
rect 4660 10832 4968 10852
rect 7116 10810 7144 11200
rect 7760 10908 8068 10928
rect 7760 10906 7766 10908
rect 7822 10906 7846 10908
rect 7902 10906 7926 10908
rect 7982 10906 8006 10908
rect 8062 10906 8068 10908
rect 7822 10854 7824 10906
rect 8004 10854 8006 10906
rect 7760 10852 7766 10854
rect 7822 10852 7846 10854
rect 7902 10852 7926 10854
rect 7982 10852 8006 10854
rect 8062 10852 8068 10854
rect 7760 10832 8068 10852
rect 9968 10810 9996 11200
rect 10860 10908 11168 10928
rect 10860 10906 10866 10908
rect 10922 10906 10946 10908
rect 11002 10906 11026 10908
rect 11082 10906 11106 10908
rect 11162 10906 11168 10908
rect 10922 10854 10924 10906
rect 11104 10854 11106 10906
rect 10860 10852 10866 10854
rect 10922 10852 10946 10854
rect 11002 10852 11026 10854
rect 11082 10852 11106 10854
rect 11162 10852 11168 10854
rect 10860 10832 11168 10852
rect 12820 10810 12848 11200
rect 13960 10908 14268 10928
rect 13960 10906 13966 10908
rect 14022 10906 14046 10908
rect 14102 10906 14126 10908
rect 14182 10906 14206 10908
rect 14262 10906 14268 10908
rect 14022 10854 14024 10906
rect 14204 10854 14206 10906
rect 13960 10852 13966 10854
rect 14022 10852 14046 10854
rect 14102 10852 14126 10854
rect 14182 10852 14206 10854
rect 14262 10852 14268 10854
rect 13960 10832 14268 10852
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 6092 10668 6144 10674
rect 6092 10610 6144 10616
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 4660 9820 4968 9840
rect 4660 9818 4666 9820
rect 4722 9818 4746 9820
rect 4802 9818 4826 9820
rect 4882 9818 4906 9820
rect 4962 9818 4968 9820
rect 4722 9766 4724 9818
rect 4904 9766 4906 9818
rect 4660 9764 4666 9766
rect 4722 9764 4746 9766
rect 4802 9764 4826 9766
rect 4882 9764 4906 9766
rect 4962 9764 4968 9766
rect 4660 9744 4968 9764
rect 5276 9722 5304 10406
rect 6012 10130 6040 10406
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5632 9648 5684 9654
rect 5684 9608 5764 9636
rect 5632 9590 5684 9596
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4908 8974 4936 9318
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4660 8732 4968 8752
rect 4660 8730 4666 8732
rect 4722 8730 4746 8732
rect 4802 8730 4826 8732
rect 4882 8730 4906 8732
rect 4962 8730 4968 8732
rect 4722 8678 4724 8730
rect 4904 8678 4906 8730
rect 4660 8676 4666 8678
rect 4722 8676 4746 8678
rect 4802 8676 4826 8678
rect 4882 8676 4906 8678
rect 4962 8676 4968 8678
rect 4660 8656 4968 8676
rect 5184 8498 5212 9386
rect 5460 8906 5488 9454
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5552 8974 5580 9318
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4660 7644 4968 7664
rect 4660 7642 4666 7644
rect 4722 7642 4746 7644
rect 4802 7642 4826 7644
rect 4882 7642 4906 7644
rect 4962 7642 4968 7644
rect 4722 7590 4724 7642
rect 4904 7590 4906 7642
rect 4660 7588 4666 7590
rect 4722 7588 4746 7590
rect 4802 7588 4826 7590
rect 4882 7588 4906 7590
rect 4962 7588 4968 7590
rect 4660 7568 4968 7588
rect 4802 7440 4858 7449
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4344 7404 4396 7410
rect 5184 7410 5212 8230
rect 5552 8022 5580 8502
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 4802 7375 4858 7384
rect 4896 7404 4948 7410
rect 4344 7346 4396 7352
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 3712 6254 3740 6802
rect 4080 6322 4108 7346
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4264 6458 4292 7142
rect 4356 6730 4384 7346
rect 4816 7342 4844 7375
rect 4896 7346 4948 7352
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4436 6928 4488 6934
rect 4436 6870 4488 6876
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4356 6390 4384 6666
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 2884 5914 2912 6190
rect 4448 6118 4476 6870
rect 4816 6730 4844 7278
rect 4908 6866 4936 7346
rect 5184 6934 5212 7346
rect 5172 6928 5224 6934
rect 5172 6870 5224 6876
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 5368 6798 5396 7346
rect 5552 7342 5580 7958
rect 5644 7546 5672 8910
rect 5736 8838 5764 9608
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6012 9178 6040 9522
rect 6104 9518 6132 10610
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 6210 10364 6518 10384
rect 6210 10362 6216 10364
rect 6272 10362 6296 10364
rect 6352 10362 6376 10364
rect 6432 10362 6456 10364
rect 6512 10362 6518 10364
rect 6272 10310 6274 10362
rect 6454 10310 6456 10362
rect 6210 10308 6216 10310
rect 6272 10308 6296 10310
rect 6352 10308 6376 10310
rect 6432 10308 6456 10310
rect 6512 10308 6518 10310
rect 6210 10288 6518 10308
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6472 9722 6500 9998
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 6104 8906 6132 9454
rect 6210 9276 6518 9296
rect 6210 9274 6216 9276
rect 6272 9274 6296 9276
rect 6352 9274 6376 9276
rect 6432 9274 6456 9276
rect 6512 9274 6518 9276
rect 6272 9222 6274 9274
rect 6454 9222 6456 9274
rect 6210 9220 6216 9222
rect 6272 9220 6296 9222
rect 6352 9220 6376 9222
rect 6432 9220 6456 9222
rect 6512 9220 6518 9222
rect 6210 9200 6518 9220
rect 6656 9110 6684 9590
rect 6932 9586 6960 10202
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7484 9586 7512 9930
rect 6920 9580 6972 9586
rect 7472 9580 7524 9586
rect 6920 9522 6972 9528
rect 7392 9540 7472 9568
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 6092 8900 6144 8906
rect 6092 8842 6144 8848
rect 6552 8900 6604 8906
rect 6552 8842 6604 8848
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5736 8498 5764 8774
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 4528 6724 4580 6730
rect 4528 6666 4580 6672
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4540 6254 4568 6666
rect 4660 6556 4968 6576
rect 4660 6554 4666 6556
rect 4722 6554 4746 6556
rect 4802 6554 4826 6556
rect 4882 6554 4906 6556
rect 4962 6554 4968 6556
rect 4722 6502 4724 6554
rect 4904 6502 4906 6554
rect 4660 6500 4666 6502
rect 4722 6500 4746 6502
rect 4802 6500 4826 6502
rect 4882 6500 4906 6502
rect 4962 6500 4968 6502
rect 4660 6480 4968 6500
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 5644 6186 5672 7482
rect 5736 7410 5764 8434
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5724 6724 5776 6730
rect 5828 6712 5856 8366
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5920 7410 5948 8230
rect 6104 7886 6132 8842
rect 6564 8566 6592 8842
rect 6656 8634 6684 9046
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6210 8188 6518 8208
rect 6210 8186 6216 8188
rect 6272 8186 6296 8188
rect 6352 8186 6376 8188
rect 6432 8186 6456 8188
rect 6512 8186 6518 8188
rect 6272 8134 6274 8186
rect 6454 8134 6456 8186
rect 6210 8132 6216 8134
rect 6272 8132 6296 8134
rect 6352 8132 6376 8134
rect 6432 8132 6456 8134
rect 6512 8132 6518 8134
rect 6210 8112 6518 8132
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 6012 6798 6040 7278
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5776 6684 5856 6712
rect 5724 6666 5776 6672
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2884 5234 2912 5850
rect 2976 5370 3004 6054
rect 3110 6012 3418 6032
rect 3110 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3276 6012
rect 3332 6010 3356 6012
rect 3412 6010 3418 6012
rect 3172 5958 3174 6010
rect 3354 5958 3356 6010
rect 3110 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3276 5958
rect 3332 5956 3356 5958
rect 3412 5956 3418 5958
rect 3110 5936 3418 5956
rect 4448 5914 4476 6054
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 3110 4924 3418 4944
rect 3110 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3276 4924
rect 3332 4922 3356 4924
rect 3412 4922 3418 4924
rect 3172 4870 3174 4922
rect 3354 4870 3356 4922
rect 3110 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3276 4870
rect 3332 4868 3356 4870
rect 3412 4868 3418 4870
rect 3110 4848 3418 4868
rect 1124 4616 1176 4622
rect 1124 4558 1176 4564
rect 1308 4616 1360 4622
rect 1308 4558 1360 4564
rect 848 4072 900 4078
rect 848 4014 900 4020
rect 860 3738 888 4014
rect 1136 3942 1164 4558
rect 1320 4078 1348 4558
rect 3528 4554 3556 5510
rect 4448 5370 4476 5578
rect 4660 5468 4968 5488
rect 4660 5466 4666 5468
rect 4722 5466 4746 5468
rect 4802 5466 4826 5468
rect 4882 5466 4906 5468
rect 4962 5466 4968 5468
rect 4722 5414 4724 5466
rect 4904 5414 4906 5466
rect 4660 5412 4666 5414
rect 4722 5412 4746 5414
rect 4802 5412 4826 5414
rect 4882 5412 4906 5414
rect 4962 5412 4968 5414
rect 4660 5392 4968 5412
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 1860 4548 1912 4554
rect 1860 4490 1912 4496
rect 3516 4548 3568 4554
rect 3516 4490 3568 4496
rect 1872 4214 1900 4490
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 3068 4214 3096 4422
rect 3620 4214 3648 5170
rect 5460 5166 5488 6122
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5552 5370 5580 6054
rect 5736 5710 5764 6666
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5920 5234 5948 5510
rect 6012 5302 6040 6258
rect 6104 5794 6132 7822
rect 7116 7750 7144 8842
rect 7208 8430 7236 9046
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 6920 7744 6972 7750
rect 7104 7744 7156 7750
rect 6972 7704 7052 7732
rect 6920 7686 6972 7692
rect 7024 7342 7052 7704
rect 7104 7686 7156 7692
rect 7300 7546 7328 8910
rect 7392 7818 7420 9540
rect 7472 9522 7524 9528
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7484 8974 7512 9318
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 6210 7100 6518 7120
rect 6210 7098 6216 7100
rect 6272 7098 6296 7100
rect 6352 7098 6376 7100
rect 6432 7098 6456 7100
rect 6512 7098 6518 7100
rect 6272 7046 6274 7098
rect 6454 7046 6456 7098
rect 6210 7044 6216 7046
rect 6272 7044 6296 7046
rect 6352 7044 6376 7046
rect 6432 7044 6456 7046
rect 6512 7044 6518 7046
rect 6210 7024 6518 7044
rect 6564 7002 6592 7278
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 7024 6934 7052 7278
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 7024 6730 7052 6870
rect 7300 6866 7328 7482
rect 7392 7342 7420 7754
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7392 7002 7420 7142
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6210 6012 6518 6032
rect 6210 6010 6216 6012
rect 6272 6010 6296 6012
rect 6352 6010 6376 6012
rect 6432 6010 6456 6012
rect 6512 6010 6518 6012
rect 6272 5958 6274 6010
rect 6454 5958 6456 6010
rect 6210 5956 6216 5958
rect 6272 5956 6296 5958
rect 6352 5956 6376 5958
rect 6432 5956 6456 5958
rect 6512 5956 6518 5958
rect 6210 5936 6518 5956
rect 6564 5914 6592 6190
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6276 5840 6328 5846
rect 6104 5788 6276 5794
rect 6104 5782 6328 5788
rect 6104 5778 6316 5782
rect 6092 5772 6316 5778
rect 6144 5766 6316 5772
rect 6092 5714 6144 5720
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 3700 4480 3752 4486
rect 3700 4422 3752 4428
rect 3712 4282 3740 4422
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 1860 4208 1912 4214
rect 1860 4150 1912 4156
rect 3056 4208 3108 4214
rect 3056 4150 3108 4156
rect 3608 4208 3660 4214
rect 3608 4150 3660 4156
rect 1308 4072 1360 4078
rect 1308 4014 1360 4020
rect 1124 3936 1176 3942
rect 1124 3878 1176 3884
rect 848 3732 900 3738
rect 848 3674 900 3680
rect 1320 3194 1348 4014
rect 1308 3188 1360 3194
rect 1308 3130 1360 3136
rect 572 2984 624 2990
rect 572 2926 624 2932
rect 584 2650 612 2926
rect 940 2848 992 2854
rect 940 2790 992 2796
rect 572 2644 624 2650
rect 572 2586 624 2592
rect 952 2446 980 2790
rect 940 2440 992 2446
rect 940 2382 992 2388
rect 848 1760 900 1766
rect 848 1702 900 1708
rect 388 1216 440 1222
rect 388 1158 440 1164
rect 400 882 428 1158
rect 860 882 888 1702
rect 1320 1358 1348 3130
rect 1872 3126 1900 4150
rect 3896 4146 3924 5102
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2700 3534 2728 3878
rect 3110 3836 3418 3856
rect 3110 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3276 3836
rect 3332 3834 3356 3836
rect 3412 3834 3418 3836
rect 3172 3782 3174 3834
rect 3354 3782 3356 3834
rect 3110 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3276 3782
rect 3332 3780 3356 3782
rect 3412 3780 3418 3782
rect 3110 3760 3418 3780
rect 3804 3738 3832 4082
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 1860 3120 1912 3126
rect 1860 3062 1912 3068
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 2056 2446 2084 2926
rect 2608 2854 2636 3334
rect 2700 3126 2728 3334
rect 2688 3120 2740 3126
rect 2688 3062 2740 3068
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2240 2106 2268 2450
rect 2228 2100 2280 2106
rect 2228 2042 2280 2048
rect 2228 1896 2280 1902
rect 2228 1838 2280 1844
rect 1308 1352 1360 1358
rect 1308 1294 1360 1300
rect 1584 1284 1636 1290
rect 1584 1226 1636 1232
rect 388 876 440 882
rect 388 818 440 824
rect 848 876 900 882
rect 848 818 900 824
rect 1308 672 1360 678
rect 1308 614 1360 620
rect 1320 270 1348 614
rect 1596 474 1624 1226
rect 2240 950 2268 1838
rect 2608 1222 2636 2790
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2792 1970 2820 2450
rect 2884 2446 2912 3538
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 3110 2748 3418 2768
rect 3110 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3276 2748
rect 3332 2746 3356 2748
rect 3412 2746 3418 2748
rect 3172 2694 3174 2746
rect 3354 2694 3356 2746
rect 3110 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3276 2694
rect 3332 2692 3356 2694
rect 3412 2692 3418 2694
rect 3110 2672 3418 2692
rect 3516 2576 3568 2582
rect 3516 2518 3568 2524
rect 3528 2446 3556 2518
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 2884 2106 2912 2382
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 2780 1964 2832 1970
rect 2780 1906 2832 1912
rect 2792 1562 2820 1906
rect 2884 1902 2912 2042
rect 2872 1896 2924 1902
rect 2872 1838 2924 1844
rect 2780 1556 2832 1562
rect 2780 1498 2832 1504
rect 2596 1216 2648 1222
rect 2596 1158 2648 1164
rect 2228 944 2280 950
rect 2228 886 2280 892
rect 2608 882 2636 1158
rect 2792 1018 2820 1498
rect 2780 1012 2832 1018
rect 2780 954 2832 960
rect 2596 876 2648 882
rect 2596 818 2648 824
rect 2608 474 2636 818
rect 1584 468 1636 474
rect 1584 410 1636 416
rect 2596 468 2648 474
rect 2596 410 2648 416
rect 2976 270 3004 2314
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3436 2106 3464 2246
rect 3424 2100 3476 2106
rect 3424 2042 3476 2048
rect 3528 1834 3556 2382
rect 3620 1902 3648 2926
rect 3712 2650 3740 2994
rect 3896 2650 3924 3878
rect 3988 3602 4016 4626
rect 4080 4622 4108 4966
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 4068 4616 4120 4622
rect 5552 4570 5580 4762
rect 5816 4752 5868 4758
rect 5816 4694 5868 4700
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 4068 4558 4120 4564
rect 5460 4554 5580 4570
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 5448 4548 5580 4554
rect 5500 4542 5580 4548
rect 5448 4490 5500 4496
rect 4660 4380 4968 4400
rect 4660 4378 4666 4380
rect 4722 4378 4746 4380
rect 4802 4378 4826 4380
rect 4882 4378 4906 4380
rect 4962 4378 4968 4380
rect 4722 4326 4724 4378
rect 4904 4326 4906 4378
rect 4660 4324 4666 4326
rect 4722 4324 4746 4326
rect 4802 4324 4826 4326
rect 4882 4324 4906 4326
rect 4962 4324 4968 4326
rect 4660 4304 4968 4324
rect 5000 4214 5028 4490
rect 4988 4208 5040 4214
rect 4988 4150 5040 4156
rect 5552 4146 5580 4542
rect 5644 4282 5672 4626
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 4080 3534 4108 3878
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3988 1902 4016 2926
rect 4172 1970 4200 2994
rect 4356 2514 4384 2994
rect 4448 2530 4476 3402
rect 4540 3058 4568 3606
rect 4908 3534 4936 4014
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 4660 3292 4968 3312
rect 4660 3290 4666 3292
rect 4722 3290 4746 3292
rect 4802 3290 4826 3292
rect 4882 3290 4906 3292
rect 4962 3290 4968 3292
rect 4722 3238 4724 3290
rect 4904 3238 4906 3290
rect 4660 3236 4666 3238
rect 4722 3236 4746 3238
rect 4802 3236 4826 3238
rect 4882 3236 4906 3238
rect 4962 3236 4968 3238
rect 4660 3216 4968 3236
rect 4528 3052 4580 3058
rect 5172 3052 5224 3058
rect 4580 3012 4660 3040
rect 4528 2994 4580 3000
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 4540 2650 4568 2790
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 4344 2508 4396 2514
rect 4448 2502 4568 2530
rect 4344 2450 4396 2456
rect 4540 2446 4568 2502
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4344 2304 4396 2310
rect 4344 2246 4396 2252
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4356 1970 4384 2246
rect 4448 1970 4476 2246
rect 4540 2038 4568 2382
rect 4632 2378 4660 3012
rect 5172 2994 5224 3000
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4724 2446 4752 2586
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4620 2372 4672 2378
rect 4620 2314 4672 2320
rect 4660 2204 4968 2224
rect 4660 2202 4666 2204
rect 4722 2202 4746 2204
rect 4802 2202 4826 2204
rect 4882 2202 4906 2204
rect 4962 2202 4968 2204
rect 4722 2150 4724 2202
rect 4904 2150 4906 2202
rect 4660 2148 4666 2150
rect 4722 2148 4746 2150
rect 4802 2148 4826 2150
rect 4882 2148 4906 2150
rect 4962 2148 4968 2150
rect 4660 2128 4968 2148
rect 4528 2032 4580 2038
rect 4528 1974 4580 1980
rect 5092 1970 5120 2790
rect 4160 1964 4212 1970
rect 4160 1906 4212 1912
rect 4344 1964 4396 1970
rect 4344 1906 4396 1912
rect 4436 1964 4488 1970
rect 4436 1906 4488 1912
rect 5080 1964 5132 1970
rect 5080 1906 5132 1912
rect 3608 1896 3660 1902
rect 3608 1838 3660 1844
rect 3976 1896 4028 1902
rect 3976 1838 4028 1844
rect 3516 1828 3568 1834
rect 3516 1770 3568 1776
rect 3110 1660 3418 1680
rect 3110 1658 3116 1660
rect 3172 1658 3196 1660
rect 3252 1658 3276 1660
rect 3332 1658 3356 1660
rect 3412 1658 3418 1660
rect 3172 1606 3174 1658
rect 3354 1606 3356 1658
rect 3110 1604 3116 1606
rect 3172 1604 3196 1606
rect 3252 1604 3276 1606
rect 3332 1604 3356 1606
rect 3412 1604 3418 1606
rect 3110 1584 3418 1604
rect 3424 1284 3476 1290
rect 3424 1226 3476 1232
rect 3436 1018 3464 1226
rect 3424 1012 3476 1018
rect 3424 954 3476 960
rect 3110 572 3418 592
rect 3110 570 3116 572
rect 3172 570 3196 572
rect 3252 570 3276 572
rect 3332 570 3356 572
rect 3412 570 3418 572
rect 3172 518 3174 570
rect 3354 518 3356 570
rect 3110 516 3116 518
rect 3172 516 3196 518
rect 3252 516 3276 518
rect 3332 516 3356 518
rect 3412 516 3418 518
rect 3110 496 3418 516
rect 3528 338 3556 1770
rect 3620 1358 3648 1838
rect 3608 1352 3660 1358
rect 3608 1294 3660 1300
rect 3620 814 3648 1294
rect 3988 1290 4016 1838
rect 3976 1284 4028 1290
rect 3976 1226 4028 1232
rect 3884 1216 3936 1222
rect 3884 1158 3936 1164
rect 3608 808 3660 814
rect 3608 750 3660 756
rect 3792 808 3844 814
rect 3792 750 3844 756
rect 3804 474 3832 750
rect 3896 678 3924 1158
rect 3988 814 4016 1226
rect 4660 1116 4968 1136
rect 4660 1114 4666 1116
rect 4722 1114 4746 1116
rect 4802 1114 4826 1116
rect 4882 1114 4906 1116
rect 4962 1114 4968 1116
rect 4722 1062 4724 1114
rect 4904 1062 4906 1114
rect 4660 1060 4666 1062
rect 4722 1060 4746 1062
rect 4802 1060 4826 1062
rect 4882 1060 4906 1062
rect 4962 1060 4968 1062
rect 4660 1040 4968 1060
rect 5184 882 5212 2994
rect 5276 2310 5304 3470
rect 5368 2650 5396 4014
rect 5828 3534 5856 4694
rect 6104 4690 6132 5306
rect 6210 4924 6518 4944
rect 6210 4922 6216 4924
rect 6272 4922 6296 4924
rect 6352 4922 6376 4924
rect 6432 4922 6456 4924
rect 6512 4922 6518 4924
rect 6272 4870 6274 4922
rect 6454 4870 6456 4922
rect 6210 4868 6216 4870
rect 6272 4868 6296 4870
rect 6352 4868 6376 4870
rect 6432 4868 6456 4870
rect 6512 4868 6518 4870
rect 6210 4848 6518 4868
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 6104 3194 6132 4626
rect 7024 4554 7052 6666
rect 7484 5370 7512 8366
rect 7576 7954 7604 8774
rect 7668 8566 7696 10406
rect 8864 10198 8892 10746
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8852 10192 8904 10198
rect 8852 10134 8904 10140
rect 7760 9820 8068 9840
rect 7760 9818 7766 9820
rect 7822 9818 7846 9820
rect 7902 9818 7926 9820
rect 7982 9818 8006 9820
rect 8062 9818 8068 9820
rect 7822 9766 7824 9818
rect 8004 9766 8006 9818
rect 7760 9764 7766 9766
rect 7822 9764 7846 9766
rect 7902 9764 7926 9766
rect 7982 9764 8006 9766
rect 8062 9764 8068 9766
rect 7760 9744 8068 9764
rect 8864 9654 8892 10134
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8496 9178 8524 9454
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8864 9330 8892 9386
rect 8772 9302 8892 9330
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 7760 8732 8068 8752
rect 7760 8730 7766 8732
rect 7822 8730 7846 8732
rect 7902 8730 7926 8732
rect 7982 8730 8006 8732
rect 8062 8730 8068 8732
rect 7822 8678 7824 8730
rect 8004 8678 8006 8730
rect 7760 8676 7766 8678
rect 7822 8676 7846 8678
rect 7902 8676 7926 8678
rect 7982 8676 8006 8678
rect 8062 8676 8068 8678
rect 7760 8656 8068 8676
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7760 7644 8068 7664
rect 7760 7642 7766 7644
rect 7822 7642 7846 7644
rect 7902 7642 7926 7644
rect 7982 7642 8006 7644
rect 8062 7642 8068 7644
rect 7822 7590 7824 7642
rect 8004 7590 8006 7642
rect 7760 7588 7766 7590
rect 7822 7588 7846 7590
rect 7902 7588 7926 7590
rect 7982 7588 8006 7590
rect 8062 7588 8068 7590
rect 7760 7568 8068 7588
rect 8128 7478 8156 8910
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8220 7750 8248 8434
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8496 7546 8524 8842
rect 8772 8634 8800 9302
rect 8852 9036 8904 9042
rect 8852 8978 8904 8984
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 7656 7472 7708 7478
rect 7656 7414 7708 7420
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 6254 7604 7142
rect 7668 6322 7696 7414
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8220 7002 8248 7278
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 7760 6556 8068 6576
rect 7760 6554 7766 6556
rect 7822 6554 7846 6556
rect 7902 6554 7926 6556
rect 7982 6554 8006 6556
rect 8062 6554 8068 6556
rect 7822 6502 7824 6554
rect 8004 6502 8006 6554
rect 7760 6500 7766 6502
rect 7822 6500 7846 6502
rect 7902 6500 7926 6502
rect 7982 6500 8006 6502
rect 8062 6500 8068 6502
rect 7760 6480 8068 6500
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 8036 5710 8064 6258
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8220 5642 8248 6938
rect 8772 6662 8800 8366
rect 8864 7954 8892 8978
rect 8956 8634 8984 10542
rect 9310 10364 9618 10384
rect 9310 10362 9316 10364
rect 9372 10362 9396 10364
rect 9452 10362 9476 10364
rect 9532 10362 9556 10364
rect 9612 10362 9618 10364
rect 9372 10310 9374 10362
rect 9554 10310 9556 10362
rect 9310 10308 9316 10310
rect 9372 10308 9396 10310
rect 9452 10308 9476 10310
rect 9532 10308 9556 10310
rect 9612 10308 9618 10310
rect 9310 10288 9618 10308
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9048 9382 9076 9454
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9048 8906 9076 9318
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8864 7546 8892 7890
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8956 7342 8984 7482
rect 9140 7410 9168 7686
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 8852 6724 8904 6730
rect 8852 6666 8904 6672
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8864 6458 8892 6666
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8312 5914 8340 6054
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8208 5636 8260 5642
rect 8208 5578 8260 5584
rect 7760 5468 8068 5488
rect 7760 5466 7766 5468
rect 7822 5466 7846 5468
rect 7902 5466 7926 5468
rect 7982 5466 8006 5468
rect 8062 5466 8068 5468
rect 7822 5414 7824 5466
rect 8004 5414 8006 5466
rect 7760 5412 7766 5414
rect 7822 5412 7846 5414
rect 7902 5412 7926 5414
rect 7982 5412 8006 5414
rect 8062 5412 8068 5414
rect 7760 5392 8068 5412
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8220 4826 8248 5102
rect 8404 5030 8432 6190
rect 8956 6186 8984 7278
rect 9048 7206 9076 7278
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 7012 4548 7064 4554
rect 7012 4490 7064 4496
rect 7024 4282 7052 4490
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6210 3836 6518 3856
rect 6210 3834 6216 3836
rect 6272 3834 6296 3836
rect 6352 3834 6376 3836
rect 6432 3834 6456 3836
rect 6512 3834 6518 3836
rect 6272 3782 6274 3834
rect 6454 3782 6456 3834
rect 6210 3780 6216 3782
rect 6272 3780 6296 3782
rect 6352 3780 6376 3782
rect 6432 3780 6456 3782
rect 6512 3780 6518 3782
rect 6210 3760 6518 3780
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 6104 2650 6132 2926
rect 6210 2748 6518 2768
rect 6210 2746 6216 2748
rect 6272 2746 6296 2748
rect 6352 2746 6376 2748
rect 6432 2746 6456 2748
rect 6512 2746 6518 2748
rect 6272 2694 6274 2746
rect 6454 2694 6456 2746
rect 6210 2692 6216 2694
rect 6272 2692 6296 2694
rect 6352 2692 6376 2694
rect 6432 2692 6456 2694
rect 6512 2692 6518 2694
rect 6210 2672 6518 2692
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 5276 1426 5304 2246
rect 5368 1766 5396 2586
rect 6564 2514 6592 3334
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5460 1970 5488 2246
rect 5448 1964 5500 1970
rect 5448 1906 5500 1912
rect 5816 1896 5868 1902
rect 5816 1838 5868 1844
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 5356 1760 5408 1766
rect 5356 1702 5408 1708
rect 5264 1420 5316 1426
rect 5264 1362 5316 1368
rect 5540 1352 5592 1358
rect 5540 1294 5592 1300
rect 5172 876 5224 882
rect 5172 818 5224 824
rect 3976 808 4028 814
rect 3976 750 4028 756
rect 5264 808 5316 814
rect 5264 750 5316 756
rect 3884 672 3936 678
rect 3884 614 3936 620
rect 5276 474 5304 750
rect 3792 468 3844 474
rect 3792 410 3844 416
rect 5264 468 5316 474
rect 5264 410 5316 416
rect 5552 406 5580 1294
rect 5828 1018 5856 1838
rect 5920 1562 5948 1838
rect 5908 1556 5960 1562
rect 5908 1498 5960 1504
rect 6012 1426 6040 2382
rect 6210 1660 6518 1680
rect 6210 1658 6216 1660
rect 6272 1658 6296 1660
rect 6352 1658 6376 1660
rect 6432 1658 6456 1660
rect 6512 1658 6518 1660
rect 6272 1606 6274 1658
rect 6454 1606 6456 1658
rect 6210 1604 6216 1606
rect 6272 1604 6296 1606
rect 6352 1604 6376 1606
rect 6432 1604 6456 1606
rect 6512 1604 6518 1606
rect 6210 1584 6518 1604
rect 6656 1562 6684 3538
rect 6840 3534 6868 3878
rect 7024 3602 7052 4218
rect 7392 4146 7420 4422
rect 7760 4380 8068 4400
rect 7760 4378 7766 4380
rect 7822 4378 7846 4380
rect 7902 4378 7926 4380
rect 7982 4378 8006 4380
rect 8062 4378 8068 4380
rect 7822 4326 7824 4378
rect 8004 4326 8006 4378
rect 7760 4324 7766 4326
rect 7822 4324 7846 4326
rect 7902 4324 7926 4326
rect 7982 4324 8006 4326
rect 8062 4324 8068 4326
rect 7760 4304 8068 4324
rect 8220 4282 8248 4558
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8220 3670 8248 4082
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 7024 3466 7052 3538
rect 7012 3460 7064 3466
rect 7012 3402 7064 3408
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6748 2650 6776 3334
rect 7024 3126 7052 3402
rect 7012 3120 7064 3126
rect 7012 3062 7064 3068
rect 7576 3058 7604 3402
rect 7760 3292 8068 3312
rect 7760 3290 7766 3292
rect 7822 3290 7846 3292
rect 7902 3290 7926 3292
rect 7982 3290 8006 3292
rect 8062 3290 8068 3292
rect 7822 3238 7824 3290
rect 8004 3238 8006 3290
rect 7760 3236 7766 3238
rect 7822 3236 7846 3238
rect 7902 3236 7926 3238
rect 7982 3236 8006 3238
rect 8062 3236 8068 3238
rect 7760 3216 8068 3236
rect 8128 3194 8156 3402
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6828 2916 6880 2922
rect 6828 2858 6880 2864
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6840 2514 6868 2858
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 6932 2038 6960 2926
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7208 2446 7236 2790
rect 8036 2582 8064 2994
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 8024 2576 8076 2582
rect 8024 2518 8076 2524
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 6920 2032 6972 2038
rect 6920 1974 6972 1980
rect 7024 1902 7052 2246
rect 7104 2100 7156 2106
rect 7104 2042 7156 2048
rect 7012 1896 7064 1902
rect 7012 1838 7064 1844
rect 6920 1828 6972 1834
rect 6920 1770 6972 1776
rect 6932 1562 6960 1770
rect 7012 1760 7064 1766
rect 7012 1702 7064 1708
rect 6644 1556 6696 1562
rect 6644 1498 6696 1504
rect 6920 1556 6972 1562
rect 6920 1498 6972 1504
rect 6656 1426 6684 1498
rect 6000 1420 6052 1426
rect 6000 1362 6052 1368
rect 6644 1420 6696 1426
rect 6644 1362 6696 1368
rect 6552 1352 6604 1358
rect 6552 1294 6604 1300
rect 6368 1284 6420 1290
rect 6368 1226 6420 1232
rect 6092 1216 6144 1222
rect 6092 1158 6144 1164
rect 5816 1012 5868 1018
rect 5816 954 5868 960
rect 5540 400 5592 406
rect 5540 342 5592 348
rect 6104 338 6132 1158
rect 6380 746 6408 1226
rect 6368 740 6420 746
rect 6368 682 6420 688
rect 6210 572 6518 592
rect 6210 570 6216 572
rect 6272 570 6296 572
rect 6352 570 6376 572
rect 6432 570 6456 572
rect 6512 570 6518 572
rect 6272 518 6274 570
rect 6454 518 6456 570
rect 6210 516 6216 518
rect 6272 516 6296 518
rect 6352 516 6376 518
rect 6432 516 6456 518
rect 6512 516 6518 518
rect 6210 496 6518 516
rect 6564 474 6592 1294
rect 7024 1222 7052 1702
rect 7116 1358 7144 2042
rect 7208 1601 7236 2382
rect 7668 1986 7696 2518
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 7760 2204 8068 2224
rect 7760 2202 7766 2204
rect 7822 2202 7846 2204
rect 7902 2202 7926 2204
rect 7982 2202 8006 2204
rect 8062 2202 8068 2204
rect 7822 2150 7824 2202
rect 8004 2150 8006 2202
rect 7760 2148 7766 2150
rect 7822 2148 7846 2150
rect 7902 2148 7926 2150
rect 7982 2148 8006 2150
rect 8062 2148 8068 2150
rect 7760 2128 8068 2148
rect 7300 1970 7696 1986
rect 8022 2000 8078 2009
rect 7288 1964 7708 1970
rect 7340 1958 7656 1964
rect 7288 1906 7340 1912
rect 7656 1906 7708 1912
rect 7932 1964 7984 1970
rect 8022 1935 8078 1944
rect 7932 1906 7984 1912
rect 7472 1828 7524 1834
rect 7472 1770 7524 1776
rect 7288 1760 7340 1766
rect 7288 1702 7340 1708
rect 7194 1592 7250 1601
rect 7194 1527 7250 1536
rect 7196 1488 7248 1494
rect 7196 1430 7248 1436
rect 7104 1352 7156 1358
rect 7104 1294 7156 1300
rect 6920 1216 6972 1222
rect 6920 1158 6972 1164
rect 7012 1216 7064 1222
rect 7012 1158 7064 1164
rect 6552 468 6604 474
rect 6552 410 6604 416
rect 3516 332 3568 338
rect 3516 274 3568 280
rect 6092 332 6144 338
rect 6092 274 6144 280
rect 1308 264 1360 270
rect 1308 206 1360 212
rect 2964 264 3016 270
rect 2964 206 3016 212
rect 6932 202 6960 1158
rect 7024 882 7052 1158
rect 7012 876 7064 882
rect 7012 818 7064 824
rect 7116 474 7144 1294
rect 7208 1290 7236 1430
rect 7196 1284 7248 1290
rect 7196 1226 7248 1232
rect 7104 468 7156 474
rect 7104 410 7156 416
rect 7300 270 7328 1702
rect 7380 1420 7432 1426
rect 7380 1362 7432 1368
rect 7392 1290 7420 1362
rect 7484 1358 7512 1770
rect 7944 1766 7972 1906
rect 8036 1902 8064 1935
rect 8024 1896 8076 1902
rect 8024 1838 8076 1844
rect 7840 1760 7892 1766
rect 7840 1702 7892 1708
rect 7932 1760 7984 1766
rect 7932 1702 7984 1708
rect 7852 1426 7880 1702
rect 8128 1494 8156 2382
rect 8220 2106 8248 3606
rect 8496 3534 8524 5306
rect 8588 5166 8616 6054
rect 8680 5710 8708 6054
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 9048 5234 9076 6054
rect 9232 5370 9260 10066
rect 10888 9994 10916 10678
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 10876 9988 10928 9994
rect 10876 9930 10928 9936
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 9864 9648 9916 9654
rect 9916 9608 9996 9636
rect 9864 9590 9916 9596
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9784 9382 9812 9522
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9310 9276 9618 9296
rect 9310 9274 9316 9276
rect 9372 9274 9396 9276
rect 9452 9274 9476 9276
rect 9532 9274 9556 9276
rect 9612 9274 9618 9276
rect 9372 9222 9374 9274
rect 9554 9222 9556 9274
rect 9310 9220 9316 9222
rect 9372 9220 9396 9222
rect 9452 9220 9476 9222
rect 9532 9220 9556 9222
rect 9612 9220 9618 9222
rect 9310 9200 9618 9220
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9416 8430 9444 8910
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9600 8498 9628 8570
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9310 8188 9618 8208
rect 9310 8186 9316 8188
rect 9372 8186 9396 8188
rect 9452 8186 9476 8188
rect 9532 8186 9556 8188
rect 9612 8186 9618 8188
rect 9372 8134 9374 8186
rect 9554 8134 9556 8186
rect 9310 8132 9316 8134
rect 9372 8132 9396 8134
rect 9452 8132 9476 8134
rect 9532 8132 9556 8134
rect 9612 8132 9618 8134
rect 9310 8112 9618 8132
rect 9784 8090 9812 9318
rect 9876 8906 9904 9386
rect 9968 9382 9996 9608
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9876 8498 9904 8842
rect 9968 8838 9996 9318
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 10152 8294 10180 8774
rect 10244 8634 10272 9862
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 10336 7342 10364 8978
rect 10520 8566 10548 9046
rect 10704 8634 10732 9862
rect 10860 9820 11168 9840
rect 10860 9818 10866 9820
rect 10922 9818 10946 9820
rect 11002 9818 11026 9820
rect 11082 9818 11106 9820
rect 11162 9818 11168 9820
rect 10922 9766 10924 9818
rect 11104 9766 11106 9818
rect 10860 9764 10866 9766
rect 10922 9764 10946 9766
rect 11002 9764 11026 9766
rect 11082 9764 11106 9766
rect 11162 9764 11168 9766
rect 10860 9744 11168 9764
rect 11256 9722 11284 10542
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11348 8974 11376 9318
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10600 8424 10652 8430
rect 10796 8412 10824 8910
rect 10860 8732 11168 8752
rect 10860 8730 10866 8732
rect 10922 8730 10946 8732
rect 11002 8730 11026 8732
rect 11082 8730 11106 8732
rect 11162 8730 11168 8732
rect 10922 8678 10924 8730
rect 11104 8678 11106 8730
rect 10860 8676 10866 8678
rect 10922 8676 10946 8678
rect 11002 8676 11026 8678
rect 11082 8676 11106 8678
rect 11162 8676 11168 8678
rect 10860 8656 11168 8676
rect 10652 8384 10824 8412
rect 10600 8366 10652 8372
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11164 7886 11192 8298
rect 11440 8294 11468 8978
rect 11532 8430 11560 10066
rect 11900 9178 11928 10610
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12410 10364 12718 10384
rect 12410 10362 12416 10364
rect 12472 10362 12496 10364
rect 12552 10362 12576 10364
rect 12632 10362 12656 10364
rect 12712 10362 12718 10364
rect 12472 10310 12474 10362
rect 12654 10310 12656 10362
rect 12410 10308 12416 10310
rect 12472 10308 12496 10310
rect 12552 10308 12576 10310
rect 12632 10308 12656 10310
rect 12712 10308 12718 10310
rect 12410 10288 12718 10308
rect 12820 10266 12848 10542
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12452 9722 12480 9862
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 11992 8498 12020 8842
rect 12084 8838 12112 9114
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11440 7954 11468 8230
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 10860 7644 11168 7664
rect 10860 7642 10866 7644
rect 10922 7642 10946 7644
rect 11002 7642 11026 7644
rect 11082 7642 11106 7644
rect 11162 7642 11168 7644
rect 10922 7590 10924 7642
rect 11104 7590 11106 7642
rect 10860 7588 10866 7590
rect 10922 7588 10946 7590
rect 11002 7588 11026 7590
rect 11082 7588 11106 7590
rect 11162 7588 11168 7590
rect 10860 7568 11168 7588
rect 11256 7546 11284 7686
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 9310 7100 9618 7120
rect 9310 7098 9316 7100
rect 9372 7098 9396 7100
rect 9452 7098 9476 7100
rect 9532 7098 9556 7100
rect 9612 7098 9618 7100
rect 9372 7046 9374 7098
rect 9554 7046 9556 7098
rect 9310 7044 9316 7046
rect 9372 7044 9396 7046
rect 9452 7044 9476 7046
rect 9532 7044 9556 7046
rect 9612 7044 9618 7046
rect 9310 7024 9618 7044
rect 10336 6798 10364 7278
rect 10784 7268 10836 7274
rect 10784 7210 10836 7216
rect 10796 7002 10824 7210
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10704 6118 10732 6666
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 9310 6012 9618 6032
rect 9310 6010 9316 6012
rect 9372 6010 9396 6012
rect 9452 6010 9476 6012
rect 9532 6010 9556 6012
rect 9612 6010 9618 6012
rect 9372 5958 9374 6010
rect 9554 5958 9556 6010
rect 9310 5956 9316 5958
rect 9372 5956 9396 5958
rect 9452 5956 9476 5958
rect 9532 5956 9556 5958
rect 9612 5956 9618 5958
rect 9310 5936 9618 5956
rect 10704 5574 10732 6054
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 9220 5364 9272 5370
rect 9140 5324 9220 5352
rect 8852 5228 8904 5234
rect 8852 5170 8904 5176
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8864 4826 8892 5170
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 9140 4690 9168 5324
rect 9220 5306 9272 5312
rect 9324 5302 9352 5510
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 10796 5234 10824 6938
rect 11072 6848 11100 7346
rect 11440 7342 11468 7890
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 10980 6820 11100 6848
rect 10980 6730 11008 6820
rect 11440 6798 11468 7142
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10860 6556 11168 6576
rect 10860 6554 10866 6556
rect 10922 6554 10946 6556
rect 11002 6554 11026 6556
rect 11082 6554 11106 6556
rect 11162 6554 11168 6556
rect 10922 6502 10924 6554
rect 11104 6502 11106 6554
rect 10860 6500 10866 6502
rect 10922 6500 10946 6502
rect 11002 6500 11026 6502
rect 11082 6500 11106 6502
rect 11162 6500 11168 6502
rect 10860 6480 11168 6500
rect 11440 5778 11468 6734
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 10860 5468 11168 5488
rect 10860 5466 10866 5468
rect 10922 5466 10946 5468
rect 11002 5466 11026 5468
rect 11082 5466 11106 5468
rect 11162 5466 11168 5468
rect 10922 5414 10924 5466
rect 11104 5414 11106 5466
rect 10860 5412 10866 5414
rect 10922 5412 10946 5414
rect 11002 5412 11026 5414
rect 11082 5412 11106 5414
rect 11162 5412 11168 5414
rect 10860 5392 11168 5412
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 9220 5092 9272 5098
rect 9220 5034 9272 5040
rect 9232 4690 9260 5034
rect 9310 4924 9618 4944
rect 9310 4922 9316 4924
rect 9372 4922 9396 4924
rect 9452 4922 9476 4924
rect 9532 4922 9556 4924
rect 9612 4922 9618 4924
rect 9372 4870 9374 4922
rect 9554 4870 9556 4922
rect 9310 4868 9316 4870
rect 9372 4868 9396 4870
rect 9452 4868 9476 4870
rect 9532 4868 9556 4870
rect 9612 4868 9618 4870
rect 9310 4848 9618 4868
rect 11348 4690 11376 5306
rect 11440 5234 11468 5714
rect 11532 5370 11560 8366
rect 11808 8090 11836 8434
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11900 7886 11928 8230
rect 12084 8022 12112 8774
rect 12176 8634 12204 9318
rect 12268 8838 12296 9454
rect 12410 9276 12718 9296
rect 12410 9274 12416 9276
rect 12472 9274 12496 9276
rect 12552 9274 12576 9276
rect 12632 9274 12656 9276
rect 12712 9274 12718 9276
rect 12472 9222 12474 9274
rect 12654 9222 12656 9274
rect 12410 9220 12416 9222
rect 12472 9220 12496 9222
rect 12552 9220 12576 9222
rect 12632 9220 12656 9222
rect 12712 9220 12718 9222
rect 12410 9200 12718 9220
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12348 8560 12400 8566
rect 12268 8520 12348 8548
rect 12072 8016 12124 8022
rect 12072 7958 12124 7964
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11716 7410 11744 7822
rect 12084 7546 12112 7958
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 12176 7410 12204 7754
rect 12268 7750 12296 8520
rect 12348 8502 12400 8508
rect 12452 8378 12480 9046
rect 12820 9042 12848 10202
rect 12912 9110 12940 10610
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12900 9104 12952 9110
rect 12900 9046 12952 9052
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12716 8968 12768 8974
rect 13004 8956 13032 9318
rect 12716 8910 12768 8916
rect 12912 8928 13032 8956
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12360 8362 12480 8378
rect 12636 8362 12664 8774
rect 12728 8634 12756 8910
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12912 8498 12940 8928
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12912 8362 12940 8434
rect 12348 8356 12480 8362
rect 12400 8350 12480 8356
rect 12624 8356 12676 8362
rect 12348 8298 12400 8304
rect 12624 8298 12676 8304
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12410 8188 12718 8208
rect 12410 8186 12416 8188
rect 12472 8186 12496 8188
rect 12552 8186 12576 8188
rect 12632 8186 12656 8188
rect 12712 8186 12718 8188
rect 12472 8134 12474 8186
rect 12654 8134 12656 8186
rect 12410 8132 12416 8134
rect 12472 8132 12496 8134
rect 12552 8132 12576 8134
rect 12632 8132 12656 8134
rect 12712 8132 12718 8134
rect 12410 8112 12718 8132
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 12268 7342 12296 7686
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12176 6390 12204 7142
rect 12268 7002 12296 7142
rect 12410 7100 12718 7120
rect 12410 7098 12416 7100
rect 12472 7098 12496 7100
rect 12552 7098 12576 7100
rect 12632 7098 12656 7100
rect 12712 7098 12718 7100
rect 12472 7046 12474 7098
rect 12654 7046 12656 7098
rect 12410 7044 12416 7046
rect 12472 7044 12496 7046
rect 12552 7044 12576 7046
rect 12632 7044 12656 7046
rect 12712 7044 12718 7046
rect 12410 7024 12718 7044
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12820 6866 12848 7278
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12820 6662 12848 6802
rect 12912 6798 12940 7346
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11716 5642 11744 6054
rect 12410 6012 12718 6032
rect 12410 6010 12416 6012
rect 12472 6010 12496 6012
rect 12552 6010 12576 6012
rect 12632 6010 12656 6012
rect 12712 6010 12718 6012
rect 12472 5958 12474 6010
rect 12654 5958 12656 6010
rect 12410 5956 12416 5958
rect 12472 5956 12496 5958
rect 12552 5956 12576 5958
rect 12632 5956 12656 5958
rect 12712 5956 12718 5958
rect 12410 5936 12718 5956
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 12820 5574 12848 6190
rect 12348 5568 12400 5574
rect 12808 5568 12860 5574
rect 12400 5516 12572 5522
rect 12348 5510 12572 5516
rect 12808 5510 12860 5516
rect 12360 5494 12572 5510
rect 12544 5370 12572 5494
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4690 11560 4966
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 8944 4548 8996 4554
rect 8944 4490 8996 4496
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8404 3194 8432 3470
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8680 2922 8708 2994
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 8680 2446 8708 2858
rect 8864 2650 8892 4082
rect 8956 4078 8984 4490
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 9140 3448 9168 4422
rect 10796 4146 10824 4422
rect 10860 4380 11168 4400
rect 10860 4378 10866 4380
rect 10922 4378 10946 4380
rect 11002 4378 11026 4380
rect 11082 4378 11106 4380
rect 11162 4378 11168 4380
rect 10922 4326 10924 4378
rect 11104 4326 11106 4378
rect 10860 4324 10866 4326
rect 10922 4324 10946 4326
rect 11002 4324 11026 4326
rect 11082 4324 11106 4326
rect 11162 4324 11168 4326
rect 10860 4304 11168 4324
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 9310 3836 9618 3856
rect 9310 3834 9316 3836
rect 9372 3834 9396 3836
rect 9452 3834 9476 3836
rect 9532 3834 9556 3836
rect 9612 3834 9618 3836
rect 9372 3782 9374 3834
rect 9554 3782 9556 3834
rect 9310 3780 9316 3782
rect 9372 3780 9396 3782
rect 9452 3780 9476 3782
rect 9532 3780 9556 3782
rect 9612 3780 9618 3782
rect 9310 3760 9618 3780
rect 11256 3738 11284 4082
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 9220 3460 9272 3466
rect 9140 3420 9220 3448
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8956 2922 8984 2994
rect 8944 2916 8996 2922
rect 8944 2858 8996 2864
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 8680 2106 8708 2382
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 8668 2100 8720 2106
rect 8668 2042 8720 2048
rect 8760 1964 8812 1970
rect 8760 1906 8812 1912
rect 8220 1834 8524 1850
rect 8220 1828 8536 1834
rect 8220 1822 8484 1828
rect 8116 1488 8168 1494
rect 8116 1430 8168 1436
rect 7840 1420 7892 1426
rect 7840 1362 7892 1368
rect 8128 1358 8156 1430
rect 7472 1352 7524 1358
rect 7472 1294 7524 1300
rect 8116 1352 8168 1358
rect 8116 1294 8168 1300
rect 7380 1284 7432 1290
rect 7380 1226 7432 1232
rect 7392 814 7420 1226
rect 7380 808 7432 814
rect 7380 750 7432 756
rect 7484 746 7512 1294
rect 8220 1222 8248 1822
rect 8484 1770 8536 1776
rect 8772 1766 8800 1906
rect 8760 1760 8812 1766
rect 8760 1702 8812 1708
rect 8208 1216 8260 1222
rect 8208 1158 8260 1164
rect 8576 1216 8628 1222
rect 8576 1158 8628 1164
rect 7760 1116 8068 1136
rect 7760 1114 7766 1116
rect 7822 1114 7846 1116
rect 7902 1114 7926 1116
rect 7982 1114 8006 1116
rect 8062 1114 8068 1116
rect 7822 1062 7824 1114
rect 8004 1062 8006 1114
rect 7760 1060 7766 1062
rect 7822 1060 7846 1062
rect 7902 1060 7926 1062
rect 7982 1060 8006 1062
rect 8062 1060 8068 1062
rect 7760 1040 8068 1060
rect 8392 944 8444 950
rect 8392 886 8444 892
rect 7472 740 7524 746
rect 7472 682 7524 688
rect 8404 474 8432 886
rect 8588 474 8616 1158
rect 8772 814 8800 1702
rect 8852 1352 8904 1358
rect 8852 1294 8904 1300
rect 8864 950 8892 1294
rect 8852 944 8904 950
rect 8852 886 8904 892
rect 8760 808 8812 814
rect 8760 750 8812 756
rect 8852 672 8904 678
rect 8852 614 8904 620
rect 8392 468 8444 474
rect 8392 410 8444 416
rect 8576 468 8628 474
rect 8576 410 8628 416
rect 8864 270 8892 614
rect 9048 338 9076 2450
rect 9140 1018 9168 3420
rect 9220 3402 9272 3408
rect 10060 3058 10088 3470
rect 11164 3380 11192 3674
rect 11164 3352 11284 3380
rect 10860 3292 11168 3312
rect 10860 3290 10866 3292
rect 10922 3290 10946 3292
rect 11002 3290 11026 3292
rect 11082 3290 11106 3292
rect 11162 3290 11168 3292
rect 10922 3238 10924 3290
rect 11104 3238 11106 3290
rect 10860 3236 10866 3238
rect 10922 3236 10946 3238
rect 11002 3236 11026 3238
rect 11082 3236 11106 3238
rect 11162 3236 11168 3238
rect 10860 3216 11168 3236
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 9310 2748 9618 2768
rect 9310 2746 9316 2748
rect 9372 2746 9396 2748
rect 9452 2746 9476 2748
rect 9532 2746 9556 2748
rect 9612 2746 9618 2748
rect 9372 2694 9374 2746
rect 9554 2694 9556 2746
rect 9310 2692 9316 2694
rect 9372 2692 9396 2694
rect 9452 2692 9476 2694
rect 9532 2692 9556 2694
rect 9612 2692 9618 2694
rect 9310 2672 9618 2692
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 9232 2310 9260 2450
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 9312 2372 9364 2378
rect 9312 2314 9364 2320
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9232 1970 9260 2246
rect 9324 2106 9352 2314
rect 9312 2100 9364 2106
rect 9312 2042 9364 2048
rect 9404 2032 9456 2038
rect 9402 2000 9404 2009
rect 9456 2000 9458 2009
rect 9220 1964 9272 1970
rect 9402 1935 9458 1944
rect 9220 1906 9272 1912
rect 9508 1902 9536 2382
rect 9772 1964 9824 1970
rect 9772 1906 9824 1912
rect 9496 1896 9548 1902
rect 9324 1844 9496 1850
rect 9324 1838 9548 1844
rect 9324 1834 9536 1838
rect 9312 1828 9536 1834
rect 9364 1822 9536 1828
rect 9312 1770 9364 1776
rect 9310 1660 9618 1680
rect 9310 1658 9316 1660
rect 9372 1658 9396 1660
rect 9452 1658 9476 1660
rect 9532 1658 9556 1660
rect 9612 1658 9618 1660
rect 9372 1606 9374 1658
rect 9554 1606 9556 1658
rect 9310 1604 9316 1606
rect 9372 1604 9396 1606
rect 9452 1604 9476 1606
rect 9532 1604 9556 1606
rect 9612 1604 9618 1606
rect 9310 1584 9618 1604
rect 9680 1556 9732 1562
rect 9680 1498 9732 1504
rect 9692 1290 9720 1498
rect 9784 1426 9812 1906
rect 9864 1760 9916 1766
rect 9864 1702 9916 1708
rect 9772 1420 9824 1426
rect 9772 1362 9824 1368
rect 9876 1358 9904 1702
rect 10060 1562 10088 2586
rect 11256 2446 11284 3352
rect 11348 2650 11376 4014
rect 11716 3942 11744 5170
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11808 4214 11836 4966
rect 12410 4924 12718 4944
rect 12410 4922 12416 4924
rect 12472 4922 12496 4924
rect 12552 4922 12576 4924
rect 12632 4922 12656 4924
rect 12712 4922 12718 4924
rect 12472 4870 12474 4922
rect 12654 4870 12656 4922
rect 12410 4868 12416 4870
rect 12472 4868 12496 4870
rect 12552 4868 12576 4870
rect 12632 4868 12656 4870
rect 12712 4868 12718 4870
rect 12410 4848 12718 4868
rect 13096 4690 13124 10678
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 13280 10130 13308 10406
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 13188 8634 13216 8842
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13648 8634 13676 8774
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13648 8022 13676 8570
rect 13832 8430 13860 10202
rect 14476 10130 14504 10406
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 13960 9820 14268 9840
rect 13960 9818 13966 9820
rect 14022 9818 14046 9820
rect 14102 9818 14126 9820
rect 14182 9818 14206 9820
rect 14262 9818 14268 9820
rect 14022 9766 14024 9818
rect 14204 9766 14206 9818
rect 13960 9764 13966 9766
rect 14022 9764 14046 9766
rect 14102 9764 14126 9766
rect 14182 9764 14206 9766
rect 14262 9764 14268 9766
rect 13960 9744 14268 9764
rect 14752 9586 14780 10406
rect 15120 10266 15148 10610
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15212 9586 15240 10406
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 14740 9444 14792 9450
rect 14740 9386 14792 9392
rect 14752 9042 14780 9386
rect 15292 9376 15344 9382
rect 15212 9336 15292 9364
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 13960 8732 14268 8752
rect 13960 8730 13966 8732
rect 14022 8730 14046 8732
rect 14102 8730 14126 8732
rect 14182 8730 14206 8732
rect 14262 8730 14268 8732
rect 14022 8678 14024 8730
rect 14204 8678 14206 8730
rect 13960 8676 13966 8678
rect 14022 8676 14046 8678
rect 14102 8676 14126 8678
rect 14182 8676 14206 8678
rect 14262 8676 14268 8678
rect 13960 8656 14268 8676
rect 14476 8634 14504 8978
rect 15212 8906 15240 9336
rect 15292 9318 15344 9324
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 14016 7886 14044 8298
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 13960 7644 14268 7664
rect 13960 7642 13966 7644
rect 14022 7642 14046 7644
rect 14102 7642 14126 7644
rect 14182 7642 14206 7644
rect 14262 7642 14268 7644
rect 14022 7590 14024 7642
rect 14204 7590 14206 7642
rect 13960 7588 13966 7590
rect 14022 7588 14046 7590
rect 14102 7588 14126 7590
rect 14182 7588 14206 7590
rect 14262 7588 14268 7590
rect 13960 7568 14268 7588
rect 14384 7478 14412 7890
rect 14188 7472 14240 7478
rect 14372 7472 14424 7478
rect 14240 7420 14320 7426
rect 14188 7414 14320 7420
rect 14372 7414 14424 7420
rect 14004 7404 14056 7410
rect 14200 7398 14320 7414
rect 14004 7346 14056 7352
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13556 6458 13584 6734
rect 14016 6730 14044 7346
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 14108 7002 14136 7210
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14292 6934 14320 7398
rect 14280 6928 14332 6934
rect 14280 6870 14332 6876
rect 14292 6746 14320 6870
rect 14384 6866 14412 7414
rect 14476 7410 14504 8570
rect 14936 8498 14964 8774
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14660 7886 14688 8298
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 14844 7886 14872 8230
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 14004 6724 14056 6730
rect 14292 6718 14412 6746
rect 14004 6666 14056 6672
rect 13960 6556 14268 6576
rect 13960 6554 13966 6556
rect 14022 6554 14046 6556
rect 14102 6554 14126 6556
rect 14182 6554 14206 6556
rect 14262 6554 14268 6556
rect 14022 6502 14024 6554
rect 14204 6502 14206 6554
rect 13960 6500 13966 6502
rect 14022 6500 14046 6502
rect 14102 6500 14126 6502
rect 14182 6500 14206 6502
rect 14262 6500 14268 6502
rect 13960 6480 14268 6500
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13832 5574 13860 6258
rect 14384 6254 14412 6718
rect 14476 6254 14504 7346
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14292 5778 14320 6054
rect 14476 5846 14504 6190
rect 14464 5840 14516 5846
rect 14464 5782 14516 5788
rect 14280 5772 14332 5778
rect 14280 5714 14332 5720
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 13960 5468 14268 5488
rect 13960 5466 13966 5468
rect 14022 5466 14046 5468
rect 14102 5466 14126 5468
rect 14182 5466 14206 5468
rect 14262 5466 14268 5468
rect 14022 5414 14024 5466
rect 14204 5414 14206 5466
rect 13960 5412 13966 5414
rect 14022 5412 14046 5414
rect 14102 5412 14126 5414
rect 14182 5412 14206 5414
rect 14262 5412 14268 5414
rect 13960 5392 14268 5412
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13268 5296 13320 5302
rect 13268 5238 13320 5244
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 12268 3738 12296 4150
rect 12452 4146 12480 4422
rect 13096 4162 13124 4626
rect 13280 4622 13308 5238
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 12440 4140 12492 4146
rect 13096 4134 13216 4162
rect 12440 4082 12492 4088
rect 13188 4078 13216 4134
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 12900 4004 12952 4010
rect 12900 3946 12952 3952
rect 12410 3836 12718 3856
rect 12410 3834 12416 3836
rect 12472 3834 12496 3836
rect 12552 3834 12576 3836
rect 12632 3834 12656 3836
rect 12712 3834 12718 3836
rect 12472 3782 12474 3834
rect 12654 3782 12656 3834
rect 12410 3780 12416 3782
rect 12472 3780 12496 3782
rect 12552 3780 12576 3782
rect 12632 3780 12656 3782
rect 12712 3780 12718 3782
rect 12410 3760 12718 3780
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 11796 3596 11848 3602
rect 11796 3538 11848 3544
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11716 2378 11744 3334
rect 11808 2854 11836 3538
rect 12912 3534 12940 3946
rect 13280 3602 13308 4558
rect 13464 4486 13492 5306
rect 14384 5030 14412 5510
rect 14476 5234 14504 5782
rect 14568 5710 14596 6598
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14660 5642 14688 6258
rect 14752 6118 14780 7754
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 15120 6458 15148 6598
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 14740 6112 14792 6118
rect 14740 6054 14792 6060
rect 15396 5914 15424 11206
rect 15580 11098 15608 11206
rect 15658 11200 15714 12000
rect 18510 11200 18566 12000
rect 18786 11248 18842 11257
rect 15672 11098 15700 11200
rect 15580 11070 15700 11098
rect 17060 10908 17368 10928
rect 17060 10906 17066 10908
rect 17122 10906 17146 10908
rect 17202 10906 17226 10908
rect 17282 10906 17306 10908
rect 17362 10906 17368 10908
rect 17122 10854 17124 10906
rect 17304 10854 17306 10906
rect 17060 10852 17066 10854
rect 17122 10852 17146 10854
rect 17202 10852 17226 10854
rect 17282 10852 17306 10854
rect 17362 10852 17368 10854
rect 17060 10832 17368 10852
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 15510 10364 15818 10384
rect 15510 10362 15516 10364
rect 15572 10362 15596 10364
rect 15652 10362 15676 10364
rect 15732 10362 15756 10364
rect 15812 10362 15818 10364
rect 15572 10310 15574 10362
rect 15754 10310 15756 10362
rect 15510 10308 15516 10310
rect 15572 10308 15596 10310
rect 15652 10308 15676 10310
rect 15732 10308 15756 10310
rect 15812 10308 15818 10310
rect 15510 10288 15818 10308
rect 16960 10130 16988 10406
rect 18064 10266 18092 10610
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16488 10056 16540 10062
rect 16540 10004 16620 10010
rect 16488 9998 16620 10004
rect 16500 9982 16620 9998
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16132 9654 16160 9862
rect 16592 9722 16620 9982
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 17060 9820 17368 9840
rect 17060 9818 17066 9820
rect 17122 9818 17146 9820
rect 17202 9818 17226 9820
rect 17282 9818 17306 9820
rect 17362 9818 17368 9820
rect 17122 9766 17124 9818
rect 17304 9766 17306 9818
rect 17060 9764 17066 9766
rect 17122 9764 17146 9766
rect 17202 9764 17226 9766
rect 17282 9764 17306 9766
rect 17362 9764 17368 9766
rect 17060 9744 17368 9764
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16120 9648 16172 9654
rect 16120 9590 16172 9596
rect 16132 9382 16160 9590
rect 18340 9518 18368 9862
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 15510 9276 15818 9296
rect 15510 9274 15516 9276
rect 15572 9274 15596 9276
rect 15652 9274 15676 9276
rect 15732 9274 15756 9276
rect 15812 9274 15818 9276
rect 15572 9222 15574 9274
rect 15754 9222 15756 9274
rect 15510 9220 15516 9222
rect 15572 9220 15596 9222
rect 15652 9220 15676 9222
rect 15732 9220 15756 9222
rect 15812 9220 15818 9222
rect 15510 9200 15818 9220
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15510 8188 15818 8208
rect 15510 8186 15516 8188
rect 15572 8186 15596 8188
rect 15652 8186 15676 8188
rect 15732 8186 15756 8188
rect 15812 8186 15818 8188
rect 15572 8134 15574 8186
rect 15754 8134 15756 8186
rect 15510 8132 15516 8134
rect 15572 8132 15596 8134
rect 15652 8132 15676 8134
rect 15732 8132 15756 8134
rect 15812 8132 15818 8134
rect 15510 8112 15818 8132
rect 15948 8022 15976 8910
rect 16132 8820 16160 9318
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 16212 8832 16264 8838
rect 16132 8792 16212 8820
rect 16212 8774 16264 8780
rect 16224 8566 16252 8774
rect 17060 8732 17368 8752
rect 17060 8730 17066 8732
rect 17122 8730 17146 8732
rect 17202 8730 17226 8732
rect 17282 8730 17306 8732
rect 17362 8730 17368 8732
rect 17122 8678 17124 8730
rect 17304 8678 17306 8730
rect 17060 8676 17066 8678
rect 17122 8676 17146 8678
rect 17202 8676 17226 8678
rect 17282 8676 17306 8678
rect 17362 8676 17368 8678
rect 17060 8656 17368 8676
rect 16212 8560 16264 8566
rect 16948 8560 17000 8566
rect 16264 8508 16344 8514
rect 16212 8502 16344 8508
rect 16948 8502 17000 8508
rect 16224 8486 16344 8502
rect 15936 8016 15988 8022
rect 15936 7958 15988 7964
rect 15510 7100 15818 7120
rect 15510 7098 15516 7100
rect 15572 7098 15596 7100
rect 15652 7098 15676 7100
rect 15732 7098 15756 7100
rect 15812 7098 15818 7100
rect 15572 7046 15574 7098
rect 15754 7046 15756 7098
rect 15510 7044 15516 7046
rect 15572 7044 15596 7046
rect 15652 7044 15676 7046
rect 15732 7044 15756 7046
rect 15812 7044 15818 7046
rect 15510 7024 15818 7044
rect 15844 6724 15896 6730
rect 15844 6666 15896 6672
rect 15856 6118 15884 6666
rect 15948 6662 15976 7958
rect 16316 7818 16344 8486
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16592 7954 16620 8366
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16776 7954 16804 8230
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16304 7812 16356 7818
rect 16304 7754 16356 7760
rect 16316 7206 16344 7754
rect 16960 7410 16988 8502
rect 17420 8430 17448 9114
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17880 7886 17908 8910
rect 18524 8090 18552 11200
rect 18786 11183 18842 11192
rect 18800 10674 18828 11183
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18616 9761 18644 9998
rect 18602 9752 18658 9761
rect 18602 9687 18658 9696
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18616 8265 18644 8434
rect 18602 8256 18658 8265
rect 18602 8191 18658 8200
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17060 7644 17368 7664
rect 17060 7642 17066 7644
rect 17122 7642 17146 7644
rect 17202 7642 17226 7644
rect 17282 7642 17306 7644
rect 17362 7642 17368 7644
rect 17122 7590 17124 7642
rect 17304 7590 17306 7642
rect 17060 7588 17066 7590
rect 17122 7588 17146 7590
rect 17202 7588 17226 7590
rect 17282 7588 17306 7590
rect 17362 7588 17368 7590
rect 17060 7568 17368 7588
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16316 6730 16344 7142
rect 17880 6866 17908 7822
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 16304 6724 16356 6730
rect 16304 6666 16356 6672
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16224 6186 16252 6394
rect 16316 6322 16344 6666
rect 16960 6458 16988 6802
rect 17500 6724 17552 6730
rect 17500 6666 17552 6672
rect 17060 6556 17368 6576
rect 17060 6554 17066 6556
rect 17122 6554 17146 6556
rect 17202 6554 17226 6556
rect 17282 6554 17306 6556
rect 17362 6554 17368 6556
rect 17122 6502 17124 6554
rect 17304 6502 17306 6554
rect 17060 6500 17066 6502
rect 17122 6500 17146 6502
rect 17202 6500 17226 6502
rect 17282 6500 17306 6502
rect 17362 6500 17368 6502
rect 17060 6480 17368 6500
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16212 6180 16264 6186
rect 16212 6122 16264 6128
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15510 6012 15818 6032
rect 15510 6010 15516 6012
rect 15572 6010 15596 6012
rect 15652 6010 15676 6012
rect 15732 6010 15756 6012
rect 15812 6010 15818 6012
rect 15572 5958 15574 6010
rect 15754 5958 15756 6010
rect 15510 5956 15516 5958
rect 15572 5956 15596 5958
rect 15652 5956 15676 5958
rect 15732 5956 15756 5958
rect 15812 5956 15818 5958
rect 15510 5936 15818 5956
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 15856 5778 15884 6054
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 16224 5710 16252 6122
rect 16500 5846 16528 6258
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 16488 5840 16540 5846
rect 16488 5782 16540 5788
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 14648 5636 14700 5642
rect 14648 5578 14700 5584
rect 16120 5636 16172 5642
rect 16120 5578 16172 5584
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 15028 5166 15056 5510
rect 16132 5302 16160 5578
rect 16224 5302 16252 5646
rect 16120 5296 16172 5302
rect 16120 5238 16172 5244
rect 16212 5296 16264 5302
rect 16212 5238 16264 5244
rect 15016 5160 15068 5166
rect 15016 5102 15068 5108
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 13452 4480 13504 4486
rect 13452 4422 13504 4428
rect 13464 4214 13492 4422
rect 13740 4282 13768 4490
rect 13960 4380 14268 4400
rect 13960 4378 13966 4380
rect 14022 4378 14046 4380
rect 14102 4378 14126 4380
rect 14182 4378 14206 4380
rect 14262 4378 14268 4380
rect 14022 4326 14024 4378
rect 14204 4326 14206 4378
rect 13960 4324 13966 4326
rect 14022 4324 14046 4326
rect 14102 4324 14126 4326
rect 14182 4324 14206 4326
rect 14262 4324 14268 4326
rect 13960 4304 14268 4324
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13452 4208 13504 4214
rect 13452 4150 13504 4156
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 12084 3058 12112 3334
rect 12544 3058 13032 3074
rect 12072 3052 12124 3058
rect 12072 2994 12124 3000
rect 12532 3052 13032 3058
rect 12584 3046 13032 3052
rect 12532 2994 12584 3000
rect 13004 2990 13032 3046
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 11992 2446 12020 2790
rect 12410 2748 12718 2768
rect 12410 2746 12416 2748
rect 12472 2746 12496 2748
rect 12552 2746 12576 2748
rect 12632 2746 12656 2748
rect 12712 2746 12718 2748
rect 12472 2694 12474 2746
rect 12654 2694 12656 2746
rect 12410 2692 12416 2694
rect 12472 2692 12496 2694
rect 12552 2692 12576 2694
rect 12632 2692 12656 2694
rect 12712 2692 12718 2694
rect 12410 2672 12718 2692
rect 12820 2650 12848 2926
rect 13004 2650 13032 2926
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 11336 2372 11388 2378
rect 11336 2314 11388 2320
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 11704 2372 11756 2378
rect 11704 2314 11756 2320
rect 10860 2204 11168 2224
rect 10860 2202 10866 2204
rect 10922 2202 10946 2204
rect 11002 2202 11026 2204
rect 11082 2202 11106 2204
rect 11162 2202 11168 2204
rect 10922 2150 10924 2202
rect 11104 2150 11106 2202
rect 10860 2148 10866 2150
rect 10922 2148 10946 2150
rect 11002 2148 11026 2150
rect 11082 2148 11106 2150
rect 11162 2148 11168 2150
rect 10860 2128 11168 2148
rect 11244 2100 11296 2106
rect 11244 2042 11296 2048
rect 10324 2032 10376 2038
rect 10138 2000 10194 2009
rect 10324 1974 10376 1980
rect 11150 2000 11206 2009
rect 10138 1935 10194 1944
rect 10152 1834 10180 1935
rect 10140 1828 10192 1834
rect 10140 1770 10192 1776
rect 10048 1556 10100 1562
rect 10048 1498 10100 1504
rect 10152 1358 10180 1770
rect 10336 1358 10364 1974
rect 10692 1964 10744 1970
rect 11150 1935 11152 1944
rect 10692 1906 10744 1912
rect 11204 1935 11206 1944
rect 11152 1906 11204 1912
rect 10704 1850 10732 1906
rect 11256 1873 11284 2042
rect 11348 2038 11376 2314
rect 11428 2304 11480 2310
rect 11428 2246 11480 2252
rect 11336 2032 11388 2038
rect 11336 1974 11388 1980
rect 11440 1970 11468 2246
rect 11624 2106 11652 2314
rect 11612 2100 11664 2106
rect 11612 2042 11664 2048
rect 11428 1964 11480 1970
rect 11428 1906 11480 1912
rect 11612 1964 11664 1970
rect 11612 1906 11664 1912
rect 11336 1896 11388 1902
rect 11242 1864 11298 1873
rect 10704 1822 11192 1850
rect 11060 1760 11112 1766
rect 11060 1702 11112 1708
rect 11072 1562 11100 1702
rect 11164 1562 11192 1822
rect 11336 1838 11388 1844
rect 11242 1799 11298 1808
rect 11348 1766 11376 1838
rect 11336 1760 11388 1766
rect 11336 1702 11388 1708
rect 11060 1556 11112 1562
rect 11060 1498 11112 1504
rect 11152 1556 11204 1562
rect 11152 1498 11204 1504
rect 11624 1494 11652 1906
rect 10784 1488 10836 1494
rect 10784 1430 10836 1436
rect 11612 1488 11664 1494
rect 11612 1430 11664 1436
rect 9864 1352 9916 1358
rect 9864 1294 9916 1300
rect 10140 1352 10192 1358
rect 10140 1294 10192 1300
rect 10324 1352 10376 1358
rect 10324 1294 10376 1300
rect 9680 1284 9732 1290
rect 9680 1226 9732 1232
rect 9128 1012 9180 1018
rect 9128 954 9180 960
rect 9312 1012 9364 1018
rect 9312 954 9364 960
rect 9324 814 9352 954
rect 9312 808 9364 814
rect 9312 750 9364 756
rect 9310 572 9618 592
rect 9310 570 9316 572
rect 9372 570 9396 572
rect 9452 570 9476 572
rect 9532 570 9556 572
rect 9612 570 9618 572
rect 9372 518 9374 570
rect 9554 518 9556 570
rect 9310 516 9316 518
rect 9372 516 9396 518
rect 9452 516 9476 518
rect 9532 516 9556 518
rect 9612 516 9618 518
rect 9310 496 9618 516
rect 9036 332 9088 338
rect 9036 274 9088 280
rect 9876 270 9904 1294
rect 10600 808 10652 814
rect 10600 750 10652 756
rect 10612 474 10640 750
rect 10600 468 10652 474
rect 10600 410 10652 416
rect 10796 270 10824 1430
rect 11336 1420 11388 1426
rect 11336 1362 11388 1368
rect 11244 1216 11296 1222
rect 11244 1158 11296 1164
rect 10860 1116 11168 1136
rect 10860 1114 10866 1116
rect 10922 1114 10946 1116
rect 11002 1114 11026 1116
rect 11082 1114 11106 1116
rect 11162 1114 11168 1116
rect 10922 1062 10924 1114
rect 11104 1062 11106 1114
rect 10860 1060 10866 1062
rect 10922 1060 10946 1062
rect 11002 1060 11026 1062
rect 11082 1060 11106 1062
rect 11162 1060 11168 1062
rect 10860 1040 11168 1060
rect 11256 338 11284 1158
rect 11348 762 11376 1362
rect 11716 762 11744 2314
rect 13188 2106 13216 2518
rect 13280 2514 13308 3538
rect 13464 3126 13492 4150
rect 13832 4078 13860 4150
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 13832 3058 13860 3334
rect 13960 3292 14268 3312
rect 13960 3290 13966 3292
rect 14022 3290 14046 3292
rect 14102 3290 14126 3292
rect 14182 3290 14206 3292
rect 14262 3290 14268 3292
rect 14022 3238 14024 3290
rect 14204 3238 14206 3290
rect 13960 3236 13966 3238
rect 14022 3236 14046 3238
rect 14102 3236 14126 3238
rect 14182 3236 14206 3238
rect 14262 3236 14268 3238
rect 13960 3216 14268 3236
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 13176 2100 13228 2106
rect 13176 2042 13228 2048
rect 12992 2032 13044 2038
rect 12992 1974 13044 1980
rect 12900 1964 12952 1970
rect 12900 1906 12952 1912
rect 12808 1760 12860 1766
rect 12808 1702 12860 1708
rect 12410 1660 12718 1680
rect 12410 1658 12416 1660
rect 12472 1658 12496 1660
rect 12552 1658 12576 1660
rect 12632 1658 12656 1660
rect 12712 1658 12718 1660
rect 12472 1606 12474 1658
rect 12654 1606 12656 1658
rect 12410 1604 12416 1606
rect 12472 1604 12496 1606
rect 12552 1604 12576 1606
rect 12632 1604 12656 1606
rect 12712 1604 12718 1606
rect 12410 1584 12718 1604
rect 11796 1488 11848 1494
rect 11796 1430 11848 1436
rect 12622 1456 12678 1465
rect 11348 734 11744 762
rect 11808 746 11836 1430
rect 12622 1391 12678 1400
rect 12256 1352 12308 1358
rect 12070 1320 12126 1329
rect 12256 1294 12308 1300
rect 12070 1255 12072 1264
rect 12124 1255 12126 1264
rect 12072 1226 12124 1232
rect 12268 1170 12296 1294
rect 12636 1222 12664 1391
rect 12820 1290 12848 1702
rect 12808 1284 12860 1290
rect 12808 1226 12860 1232
rect 12912 1222 12940 1906
rect 12176 1142 12296 1170
rect 12624 1216 12676 1222
rect 12624 1158 12676 1164
rect 12900 1216 12952 1222
rect 12900 1158 12952 1164
rect 12176 950 12204 1142
rect 12164 944 12216 950
rect 12164 886 12216 892
rect 12900 944 12952 950
rect 13004 932 13032 1974
rect 13084 1964 13136 1970
rect 13084 1906 13136 1912
rect 12952 904 13032 932
rect 12900 886 12952 892
rect 12348 876 12400 882
rect 12808 876 12860 882
rect 12400 836 12808 864
rect 12348 818 12400 824
rect 12808 818 12860 824
rect 11244 332 11296 338
rect 11244 274 11296 280
rect 7288 264 7340 270
rect 7288 206 7340 212
rect 8852 264 8904 270
rect 8852 206 8904 212
rect 9864 264 9916 270
rect 9864 206 9916 212
rect 10784 264 10836 270
rect 10784 206 10836 212
rect 11348 202 11376 734
rect 11716 678 11744 734
rect 11796 740 11848 746
rect 11796 682 11848 688
rect 11612 672 11664 678
rect 11612 614 11664 620
rect 11704 672 11756 678
rect 11704 614 11756 620
rect 11624 270 11652 614
rect 12410 572 12718 592
rect 12410 570 12416 572
rect 12472 570 12496 572
rect 12552 570 12576 572
rect 12632 570 12656 572
rect 12712 570 12718 572
rect 12472 518 12474 570
rect 12654 518 12656 570
rect 12410 516 12416 518
rect 12472 516 12496 518
rect 12552 516 12576 518
rect 12632 516 12656 518
rect 12712 516 12718 518
rect 12410 496 12718 516
rect 12820 270 12848 818
rect 13096 474 13124 1906
rect 13544 1352 13596 1358
rect 13542 1320 13544 1329
rect 13596 1320 13598 1329
rect 13176 1284 13228 1290
rect 13740 1290 13768 2450
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13832 2106 13860 2314
rect 13960 2204 14268 2224
rect 13960 2202 13966 2204
rect 14022 2202 14046 2204
rect 14102 2202 14126 2204
rect 14182 2202 14206 2204
rect 14262 2202 14268 2204
rect 14022 2150 14024 2202
rect 14204 2150 14206 2202
rect 13960 2148 13966 2150
rect 14022 2148 14046 2150
rect 14102 2148 14126 2150
rect 14182 2148 14206 2150
rect 14262 2148 14268 2150
rect 13960 2128 14268 2148
rect 13820 2100 13872 2106
rect 13820 2042 13872 2048
rect 14384 1970 14412 2790
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14372 1964 14424 1970
rect 14372 1906 14424 1912
rect 14476 1902 14504 2246
rect 13912 1896 13964 1902
rect 14464 1896 14516 1902
rect 13964 1844 14320 1850
rect 13912 1838 14320 1844
rect 14464 1838 14516 1844
rect 13924 1822 14320 1838
rect 14188 1760 14240 1766
rect 14188 1702 14240 1708
rect 14200 1494 14228 1702
rect 14292 1494 14320 1822
rect 14188 1488 14240 1494
rect 14188 1430 14240 1436
rect 14280 1488 14332 1494
rect 14568 1465 14596 4082
rect 15028 4078 15056 4558
rect 15212 4486 15240 4966
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15304 4146 15332 4966
rect 15396 4554 15424 5102
rect 15510 4924 15818 4944
rect 15510 4922 15516 4924
rect 15572 4922 15596 4924
rect 15652 4922 15676 4924
rect 15732 4922 15756 4924
rect 15812 4922 15818 4924
rect 15572 4870 15574 4922
rect 15754 4870 15756 4922
rect 15510 4868 15516 4870
rect 15572 4868 15596 4870
rect 15652 4868 15676 4870
rect 15732 4868 15756 4870
rect 15812 4868 15818 4870
rect 15510 4848 15818 4868
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14752 3602 14780 3878
rect 14740 3596 14792 3602
rect 14792 3556 14872 3584
rect 14740 3538 14792 3544
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14660 3058 14688 3334
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14752 2990 14780 3334
rect 14844 3058 14872 3556
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14740 2100 14792 2106
rect 14740 2042 14792 2048
rect 14752 1873 14780 2042
rect 14936 1970 14964 3470
rect 15028 3194 15056 4014
rect 15212 3738 15240 4014
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15016 3188 15068 3194
rect 15016 3130 15068 3136
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 15120 2446 15148 2586
rect 15108 2440 15160 2446
rect 15160 2400 15240 2428
rect 15108 2382 15160 2388
rect 15108 2100 15160 2106
rect 15108 2042 15160 2048
rect 14832 1964 14884 1970
rect 14832 1906 14884 1912
rect 14924 1964 14976 1970
rect 14924 1906 14976 1912
rect 14738 1864 14794 1873
rect 14738 1799 14794 1808
rect 14740 1760 14792 1766
rect 14740 1702 14792 1708
rect 14752 1578 14780 1702
rect 14660 1562 14780 1578
rect 14844 1562 14872 1906
rect 14648 1556 14780 1562
rect 14700 1550 14780 1556
rect 14832 1556 14884 1562
rect 14648 1498 14700 1504
rect 14832 1498 14884 1504
rect 14280 1430 14332 1436
rect 14554 1456 14610 1465
rect 15120 1426 15148 2042
rect 14554 1391 14610 1400
rect 15108 1420 15160 1426
rect 15108 1362 15160 1368
rect 14096 1352 14148 1358
rect 14148 1300 14412 1306
rect 14096 1294 14412 1300
rect 13542 1255 13598 1264
rect 13728 1284 13780 1290
rect 13176 1226 13228 1232
rect 14108 1278 14412 1294
rect 13728 1226 13780 1232
rect 13188 882 13216 1226
rect 13740 1018 13768 1226
rect 13820 1216 13872 1222
rect 13820 1158 13872 1164
rect 13728 1012 13780 1018
rect 13728 954 13780 960
rect 13832 950 13860 1158
rect 13960 1116 14268 1136
rect 13960 1114 13966 1116
rect 14022 1114 14046 1116
rect 14102 1114 14126 1116
rect 14182 1114 14206 1116
rect 14262 1114 14268 1116
rect 14022 1062 14024 1114
rect 14204 1062 14206 1114
rect 13960 1060 13966 1062
rect 14022 1060 14046 1062
rect 14102 1060 14126 1062
rect 14182 1060 14206 1062
rect 14262 1060 14268 1062
rect 13960 1040 14268 1060
rect 14384 1018 14412 1278
rect 14464 1216 14516 1222
rect 14464 1158 14516 1164
rect 15016 1216 15068 1222
rect 15016 1158 15068 1164
rect 14372 1012 14424 1018
rect 14372 954 14424 960
rect 13820 944 13872 950
rect 13820 886 13872 892
rect 14476 882 14504 1158
rect 13176 876 13228 882
rect 13176 818 13228 824
rect 14464 876 14516 882
rect 14464 818 14516 824
rect 13084 468 13136 474
rect 13084 410 13136 416
rect 13188 338 13216 818
rect 14740 672 14792 678
rect 14740 614 14792 620
rect 13176 332 13228 338
rect 13176 274 13228 280
rect 14752 270 14780 614
rect 15028 474 15056 1158
rect 15212 814 15240 2400
rect 15396 2038 15424 4490
rect 15510 3836 15818 3856
rect 15510 3834 15516 3836
rect 15572 3834 15596 3836
rect 15652 3834 15676 3836
rect 15732 3834 15756 3836
rect 15812 3834 15818 3836
rect 15572 3782 15574 3834
rect 15754 3782 15756 3834
rect 15510 3780 15516 3782
rect 15572 3780 15596 3782
rect 15652 3780 15676 3782
rect 15732 3780 15756 3782
rect 15812 3780 15818 3782
rect 15510 3760 15818 3780
rect 15856 3534 15884 4558
rect 16132 4486 16160 5238
rect 16592 5098 16620 6190
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 16960 5166 16988 5850
rect 17060 5468 17368 5488
rect 17060 5466 17066 5468
rect 17122 5466 17146 5468
rect 17202 5466 17226 5468
rect 17282 5466 17306 5468
rect 17362 5466 17368 5468
rect 17122 5414 17124 5466
rect 17304 5414 17306 5466
rect 17060 5412 17066 5414
rect 17122 5412 17146 5414
rect 17202 5412 17226 5414
rect 17282 5412 17306 5414
rect 17362 5412 17368 5414
rect 17060 5392 17368 5412
rect 17420 5234 17448 6190
rect 17512 5778 17540 6666
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 17880 5710 17908 6802
rect 18512 6792 18564 6798
rect 18510 6760 18512 6769
rect 18564 6760 18566 6769
rect 18510 6695 18566 6704
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18340 5778 18368 6598
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 16120 4480 16172 4486
rect 16120 4422 16172 4428
rect 16132 4214 16160 4422
rect 16120 4208 16172 4214
rect 16120 4150 16172 4156
rect 16592 4146 16620 4626
rect 17060 4380 17368 4400
rect 17060 4378 17066 4380
rect 17122 4378 17146 4380
rect 17202 4378 17226 4380
rect 17282 4378 17306 4380
rect 17362 4378 17368 4380
rect 17122 4326 17124 4378
rect 17304 4326 17306 4378
rect 17060 4324 17066 4326
rect 17122 4324 17146 4326
rect 17202 4324 17226 4326
rect 17282 4324 17306 4326
rect 17362 4324 17368 4326
rect 17060 4304 17368 4324
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15844 3392 15896 3398
rect 15948 3380 15976 4014
rect 16408 3466 16436 4014
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 16396 3460 16448 3466
rect 16396 3402 16448 3408
rect 17408 3460 17460 3466
rect 17408 3402 17460 3408
rect 15896 3352 15976 3380
rect 15844 3334 15896 3340
rect 15856 3126 15884 3334
rect 16132 3194 16160 3402
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 15844 3120 15896 3126
rect 15844 3062 15896 3068
rect 16408 2922 16436 3402
rect 16856 3392 16908 3398
rect 16856 3334 16908 3340
rect 16868 3058 16896 3334
rect 17060 3292 17368 3312
rect 17060 3290 17066 3292
rect 17122 3290 17146 3292
rect 17202 3290 17226 3292
rect 17282 3290 17306 3292
rect 17362 3290 17368 3292
rect 17122 3238 17124 3290
rect 17304 3238 17306 3290
rect 17060 3236 17066 3238
rect 17122 3236 17146 3238
rect 17202 3236 17226 3238
rect 17282 3236 17306 3238
rect 17362 3236 17368 3238
rect 17060 3216 17368 3236
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 17132 2848 17184 2854
rect 17132 2790 17184 2796
rect 15510 2748 15818 2768
rect 15510 2746 15516 2748
rect 15572 2746 15596 2748
rect 15652 2746 15676 2748
rect 15732 2746 15756 2748
rect 15812 2746 15818 2748
rect 15572 2694 15574 2746
rect 15754 2694 15756 2746
rect 15510 2692 15516 2694
rect 15572 2692 15596 2694
rect 15652 2692 15676 2694
rect 15732 2692 15756 2694
rect 15812 2692 15818 2694
rect 15510 2672 15818 2692
rect 17144 2650 17172 2790
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17144 2446 17172 2586
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 15384 2032 15436 2038
rect 15384 1974 15436 1980
rect 15488 1902 15516 2314
rect 17060 2204 17368 2224
rect 17060 2202 17066 2204
rect 17122 2202 17146 2204
rect 17202 2202 17226 2204
rect 17282 2202 17306 2204
rect 17362 2202 17368 2204
rect 17122 2150 17124 2202
rect 17304 2150 17306 2202
rect 17060 2148 17066 2150
rect 17122 2148 17146 2150
rect 17202 2148 17226 2150
rect 17282 2148 17306 2150
rect 17362 2148 17368 2150
rect 17060 2128 17368 2148
rect 17420 2038 17448 3402
rect 17512 2106 17540 4626
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17788 3058 17816 4422
rect 17972 4282 18000 5306
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 18064 4010 18092 5510
rect 18524 5273 18552 5646
rect 18510 5264 18566 5273
rect 18510 5199 18566 5208
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 18052 4004 18104 4010
rect 18052 3946 18104 3952
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17684 2984 17736 2990
rect 17684 2926 17736 2932
rect 17696 2650 17724 2926
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 17788 2582 17816 2994
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 17880 2446 17908 2790
rect 18156 2446 18184 2858
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 17880 2281 17908 2382
rect 18236 2372 18288 2378
rect 18236 2314 18288 2320
rect 17866 2272 17922 2281
rect 17866 2207 17922 2216
rect 18248 2106 18276 2314
rect 17500 2100 17552 2106
rect 17500 2042 17552 2048
rect 18236 2100 18288 2106
rect 18236 2042 18288 2048
rect 17408 2032 17460 2038
rect 17408 1974 17460 1980
rect 16488 1964 16540 1970
rect 16488 1906 16540 1912
rect 15476 1896 15528 1902
rect 15476 1838 15528 1844
rect 16120 1896 16172 1902
rect 16120 1838 16172 1844
rect 15510 1660 15818 1680
rect 15510 1658 15516 1660
rect 15572 1658 15596 1660
rect 15652 1658 15676 1660
rect 15732 1658 15756 1660
rect 15812 1658 15818 1660
rect 15572 1606 15574 1658
rect 15754 1606 15756 1658
rect 15510 1604 15516 1606
rect 15572 1604 15596 1606
rect 15652 1604 15676 1606
rect 15732 1604 15756 1606
rect 15812 1604 15818 1606
rect 15510 1584 15818 1604
rect 15660 1420 15712 1426
rect 15660 1362 15712 1368
rect 15200 808 15252 814
rect 15200 750 15252 756
rect 15672 746 15700 1362
rect 16132 1358 16160 1838
rect 16120 1352 16172 1358
rect 16120 1294 16172 1300
rect 16396 1284 16448 1290
rect 16396 1226 16448 1232
rect 15844 1216 15896 1222
rect 15844 1158 15896 1164
rect 15856 950 15884 1158
rect 16408 1018 16436 1226
rect 16500 1018 16528 1906
rect 16672 1760 16724 1766
rect 16672 1702 16724 1708
rect 16396 1012 16448 1018
rect 16396 954 16448 960
rect 16488 1012 16540 1018
rect 16488 954 16540 960
rect 15844 944 15896 950
rect 15844 886 15896 892
rect 16580 876 16632 882
rect 16580 818 16632 824
rect 15660 740 15712 746
rect 15660 682 15712 688
rect 15510 572 15818 592
rect 15510 570 15516 572
rect 15572 570 15596 572
rect 15652 570 15676 572
rect 15732 570 15756 572
rect 15812 570 15818 572
rect 15572 518 15574 570
rect 15754 518 15756 570
rect 15510 516 15516 518
rect 15572 516 15596 518
rect 15652 516 15676 518
rect 15732 516 15756 518
rect 15812 516 15818 518
rect 15510 496 15818 516
rect 15016 468 15068 474
rect 15016 410 15068 416
rect 16592 270 16620 818
rect 16684 338 16712 1702
rect 17060 1116 17368 1136
rect 17060 1114 17066 1116
rect 17122 1114 17146 1116
rect 17202 1114 17226 1116
rect 17282 1114 17306 1116
rect 17362 1114 17368 1116
rect 17122 1062 17124 1114
rect 17304 1062 17306 1114
rect 17060 1060 17066 1062
rect 17122 1060 17146 1062
rect 17202 1060 17226 1062
rect 17282 1060 17306 1062
rect 17362 1060 17368 1062
rect 17060 1040 17368 1060
rect 17420 1018 17448 1974
rect 17868 1216 17920 1222
rect 17868 1158 17920 1164
rect 17408 1012 17460 1018
rect 17408 954 17460 960
rect 17224 876 17276 882
rect 17224 818 17276 824
rect 16948 808 17000 814
rect 16948 750 17000 756
rect 16960 474 16988 750
rect 17236 474 17264 818
rect 16948 468 17000 474
rect 16948 410 17000 416
rect 17224 468 17276 474
rect 17224 410 17276 416
rect 16672 332 16724 338
rect 16672 274 16724 280
rect 17880 270 17908 1158
rect 18340 882 18368 4082
rect 18510 3768 18566 3777
rect 18510 3703 18566 3712
rect 18524 3534 18552 3703
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18328 876 18380 882
rect 18328 818 18380 824
rect 18512 808 18564 814
rect 18510 776 18512 785
rect 18564 776 18566 785
rect 18510 711 18566 720
rect 18524 474 18552 711
rect 18512 468 18564 474
rect 18512 410 18564 416
rect 11612 264 11664 270
rect 11612 206 11664 212
rect 12808 264 12860 270
rect 12808 206 12860 212
rect 14740 264 14792 270
rect 14740 206 14792 212
rect 16580 264 16632 270
rect 16580 206 16632 212
rect 17868 264 17920 270
rect 17868 206 17920 212
rect 6920 196 6972 202
rect 6920 138 6972 144
rect 11336 196 11388 202
rect 11336 138 11388 144
rect 4660 28 4968 48
rect 4660 26 4666 28
rect 4722 26 4746 28
rect 4802 26 4826 28
rect 4882 26 4906 28
rect 4962 26 4968 28
rect 4722 -26 4724 26
rect 4904 -26 4906 26
rect 4660 -28 4666 -26
rect 4722 -28 4746 -26
rect 4802 -28 4826 -26
rect 4882 -28 4906 -26
rect 4962 -28 4968 -26
rect 4660 -48 4968 -28
rect 7760 28 8068 48
rect 7760 26 7766 28
rect 7822 26 7846 28
rect 7902 26 7926 28
rect 7982 26 8006 28
rect 8062 26 8068 28
rect 7822 -26 7824 26
rect 8004 -26 8006 26
rect 7760 -28 7766 -26
rect 7822 -28 7846 -26
rect 7902 -28 7926 -26
rect 7982 -28 8006 -26
rect 8062 -28 8068 -26
rect 7760 -48 8068 -28
rect 10860 28 11168 48
rect 10860 26 10866 28
rect 10922 26 10946 28
rect 11002 26 11026 28
rect 11082 26 11106 28
rect 11162 26 11168 28
rect 10922 -26 10924 26
rect 11104 -26 11106 26
rect 10860 -28 10866 -26
rect 10922 -28 10946 -26
rect 11002 -28 11026 -26
rect 11082 -28 11106 -26
rect 11162 -28 11168 -26
rect 10860 -48 11168 -28
rect 13960 28 14268 48
rect 13960 26 13966 28
rect 14022 26 14046 28
rect 14102 26 14126 28
rect 14182 26 14206 28
rect 14262 26 14268 28
rect 14022 -26 14024 26
rect 14204 -26 14206 26
rect 13960 -28 13966 -26
rect 14022 -28 14046 -26
rect 14102 -28 14126 -26
rect 14182 -28 14206 -26
rect 14262 -28 14268 -26
rect 13960 -48 14268 -28
rect 17060 28 17368 48
rect 17060 26 17066 28
rect 17122 26 17146 28
rect 17202 26 17226 28
rect 17282 26 17306 28
rect 17362 26 17368 28
rect 17122 -26 17124 26
rect 17304 -26 17306 26
rect 17060 -28 17066 -26
rect 17122 -28 17146 -26
rect 17202 -28 17226 -26
rect 17282 -28 17306 -26
rect 17362 -28 17368 -26
rect 17060 -48 17368 -28
<< via2 >>
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 3276 10362 3332 10364
rect 3356 10362 3412 10364
rect 3116 10310 3162 10362
rect 3162 10310 3172 10362
rect 3196 10310 3226 10362
rect 3226 10310 3238 10362
rect 3238 10310 3252 10362
rect 3276 10310 3290 10362
rect 3290 10310 3302 10362
rect 3302 10310 3332 10362
rect 3356 10310 3366 10362
rect 3366 10310 3412 10362
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 3276 10308 3332 10310
rect 3356 10308 3412 10310
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 3276 9274 3332 9276
rect 3356 9274 3412 9276
rect 3116 9222 3162 9274
rect 3162 9222 3172 9274
rect 3196 9222 3226 9274
rect 3226 9222 3238 9274
rect 3238 9222 3252 9274
rect 3276 9222 3290 9274
rect 3290 9222 3302 9274
rect 3302 9222 3332 9274
rect 3356 9222 3366 9274
rect 3366 9222 3412 9274
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3276 9220 3332 9222
rect 3356 9220 3412 9222
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 3276 8186 3332 8188
rect 3356 8186 3412 8188
rect 3116 8134 3162 8186
rect 3162 8134 3172 8186
rect 3196 8134 3226 8186
rect 3226 8134 3238 8186
rect 3238 8134 3252 8186
rect 3276 8134 3290 8186
rect 3290 8134 3302 8186
rect 3302 8134 3332 8186
rect 3356 8134 3366 8186
rect 3366 8134 3412 8186
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 3276 8132 3332 8134
rect 3356 8132 3412 8134
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 3276 7098 3332 7100
rect 3356 7098 3412 7100
rect 3116 7046 3162 7098
rect 3162 7046 3172 7098
rect 3196 7046 3226 7098
rect 3226 7046 3238 7098
rect 3238 7046 3252 7098
rect 3276 7046 3290 7098
rect 3290 7046 3302 7098
rect 3302 7046 3332 7098
rect 3356 7046 3366 7098
rect 3366 7046 3412 7098
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3276 7044 3332 7046
rect 3356 7044 3412 7046
rect 3790 7420 3792 7440
rect 3792 7420 3844 7440
rect 3844 7420 3846 7440
rect 3790 7384 3846 7420
rect 4666 10906 4722 10908
rect 4746 10906 4802 10908
rect 4826 10906 4882 10908
rect 4906 10906 4962 10908
rect 4666 10854 4712 10906
rect 4712 10854 4722 10906
rect 4746 10854 4776 10906
rect 4776 10854 4788 10906
rect 4788 10854 4802 10906
rect 4826 10854 4840 10906
rect 4840 10854 4852 10906
rect 4852 10854 4882 10906
rect 4906 10854 4916 10906
rect 4916 10854 4962 10906
rect 4666 10852 4722 10854
rect 4746 10852 4802 10854
rect 4826 10852 4882 10854
rect 4906 10852 4962 10854
rect 7766 10906 7822 10908
rect 7846 10906 7902 10908
rect 7926 10906 7982 10908
rect 8006 10906 8062 10908
rect 7766 10854 7812 10906
rect 7812 10854 7822 10906
rect 7846 10854 7876 10906
rect 7876 10854 7888 10906
rect 7888 10854 7902 10906
rect 7926 10854 7940 10906
rect 7940 10854 7952 10906
rect 7952 10854 7982 10906
rect 8006 10854 8016 10906
rect 8016 10854 8062 10906
rect 7766 10852 7822 10854
rect 7846 10852 7902 10854
rect 7926 10852 7982 10854
rect 8006 10852 8062 10854
rect 10866 10906 10922 10908
rect 10946 10906 11002 10908
rect 11026 10906 11082 10908
rect 11106 10906 11162 10908
rect 10866 10854 10912 10906
rect 10912 10854 10922 10906
rect 10946 10854 10976 10906
rect 10976 10854 10988 10906
rect 10988 10854 11002 10906
rect 11026 10854 11040 10906
rect 11040 10854 11052 10906
rect 11052 10854 11082 10906
rect 11106 10854 11116 10906
rect 11116 10854 11162 10906
rect 10866 10852 10922 10854
rect 10946 10852 11002 10854
rect 11026 10852 11082 10854
rect 11106 10852 11162 10854
rect 13966 10906 14022 10908
rect 14046 10906 14102 10908
rect 14126 10906 14182 10908
rect 14206 10906 14262 10908
rect 13966 10854 14012 10906
rect 14012 10854 14022 10906
rect 14046 10854 14076 10906
rect 14076 10854 14088 10906
rect 14088 10854 14102 10906
rect 14126 10854 14140 10906
rect 14140 10854 14152 10906
rect 14152 10854 14182 10906
rect 14206 10854 14216 10906
rect 14216 10854 14262 10906
rect 13966 10852 14022 10854
rect 14046 10852 14102 10854
rect 14126 10852 14182 10854
rect 14206 10852 14262 10854
rect 4666 9818 4722 9820
rect 4746 9818 4802 9820
rect 4826 9818 4882 9820
rect 4906 9818 4962 9820
rect 4666 9766 4712 9818
rect 4712 9766 4722 9818
rect 4746 9766 4776 9818
rect 4776 9766 4788 9818
rect 4788 9766 4802 9818
rect 4826 9766 4840 9818
rect 4840 9766 4852 9818
rect 4852 9766 4882 9818
rect 4906 9766 4916 9818
rect 4916 9766 4962 9818
rect 4666 9764 4722 9766
rect 4746 9764 4802 9766
rect 4826 9764 4882 9766
rect 4906 9764 4962 9766
rect 4666 8730 4722 8732
rect 4746 8730 4802 8732
rect 4826 8730 4882 8732
rect 4906 8730 4962 8732
rect 4666 8678 4712 8730
rect 4712 8678 4722 8730
rect 4746 8678 4776 8730
rect 4776 8678 4788 8730
rect 4788 8678 4802 8730
rect 4826 8678 4840 8730
rect 4840 8678 4852 8730
rect 4852 8678 4882 8730
rect 4906 8678 4916 8730
rect 4916 8678 4962 8730
rect 4666 8676 4722 8678
rect 4746 8676 4802 8678
rect 4826 8676 4882 8678
rect 4906 8676 4962 8678
rect 4666 7642 4722 7644
rect 4746 7642 4802 7644
rect 4826 7642 4882 7644
rect 4906 7642 4962 7644
rect 4666 7590 4712 7642
rect 4712 7590 4722 7642
rect 4746 7590 4776 7642
rect 4776 7590 4788 7642
rect 4788 7590 4802 7642
rect 4826 7590 4840 7642
rect 4840 7590 4852 7642
rect 4852 7590 4882 7642
rect 4906 7590 4916 7642
rect 4916 7590 4962 7642
rect 4666 7588 4722 7590
rect 4746 7588 4802 7590
rect 4826 7588 4882 7590
rect 4906 7588 4962 7590
rect 4802 7384 4858 7440
rect 6216 10362 6272 10364
rect 6296 10362 6352 10364
rect 6376 10362 6432 10364
rect 6456 10362 6512 10364
rect 6216 10310 6262 10362
rect 6262 10310 6272 10362
rect 6296 10310 6326 10362
rect 6326 10310 6338 10362
rect 6338 10310 6352 10362
rect 6376 10310 6390 10362
rect 6390 10310 6402 10362
rect 6402 10310 6432 10362
rect 6456 10310 6466 10362
rect 6466 10310 6512 10362
rect 6216 10308 6272 10310
rect 6296 10308 6352 10310
rect 6376 10308 6432 10310
rect 6456 10308 6512 10310
rect 6216 9274 6272 9276
rect 6296 9274 6352 9276
rect 6376 9274 6432 9276
rect 6456 9274 6512 9276
rect 6216 9222 6262 9274
rect 6262 9222 6272 9274
rect 6296 9222 6326 9274
rect 6326 9222 6338 9274
rect 6338 9222 6352 9274
rect 6376 9222 6390 9274
rect 6390 9222 6402 9274
rect 6402 9222 6432 9274
rect 6456 9222 6466 9274
rect 6466 9222 6512 9274
rect 6216 9220 6272 9222
rect 6296 9220 6352 9222
rect 6376 9220 6432 9222
rect 6456 9220 6512 9222
rect 4666 6554 4722 6556
rect 4746 6554 4802 6556
rect 4826 6554 4882 6556
rect 4906 6554 4962 6556
rect 4666 6502 4712 6554
rect 4712 6502 4722 6554
rect 4746 6502 4776 6554
rect 4776 6502 4788 6554
rect 4788 6502 4802 6554
rect 4826 6502 4840 6554
rect 4840 6502 4852 6554
rect 4852 6502 4882 6554
rect 4906 6502 4916 6554
rect 4916 6502 4962 6554
rect 4666 6500 4722 6502
rect 4746 6500 4802 6502
rect 4826 6500 4882 6502
rect 4906 6500 4962 6502
rect 6216 8186 6272 8188
rect 6296 8186 6352 8188
rect 6376 8186 6432 8188
rect 6456 8186 6512 8188
rect 6216 8134 6262 8186
rect 6262 8134 6272 8186
rect 6296 8134 6326 8186
rect 6326 8134 6338 8186
rect 6338 8134 6352 8186
rect 6376 8134 6390 8186
rect 6390 8134 6402 8186
rect 6402 8134 6432 8186
rect 6456 8134 6466 8186
rect 6466 8134 6512 8186
rect 6216 8132 6272 8134
rect 6296 8132 6352 8134
rect 6376 8132 6432 8134
rect 6456 8132 6512 8134
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 3276 6010 3332 6012
rect 3356 6010 3412 6012
rect 3116 5958 3162 6010
rect 3162 5958 3172 6010
rect 3196 5958 3226 6010
rect 3226 5958 3238 6010
rect 3238 5958 3252 6010
rect 3276 5958 3290 6010
rect 3290 5958 3302 6010
rect 3302 5958 3332 6010
rect 3356 5958 3366 6010
rect 3366 5958 3412 6010
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 3276 5956 3332 5958
rect 3356 5956 3412 5958
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 3276 4922 3332 4924
rect 3356 4922 3412 4924
rect 3116 4870 3162 4922
rect 3162 4870 3172 4922
rect 3196 4870 3226 4922
rect 3226 4870 3238 4922
rect 3238 4870 3252 4922
rect 3276 4870 3290 4922
rect 3290 4870 3302 4922
rect 3302 4870 3332 4922
rect 3356 4870 3366 4922
rect 3366 4870 3412 4922
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 3276 4868 3332 4870
rect 3356 4868 3412 4870
rect 4666 5466 4722 5468
rect 4746 5466 4802 5468
rect 4826 5466 4882 5468
rect 4906 5466 4962 5468
rect 4666 5414 4712 5466
rect 4712 5414 4722 5466
rect 4746 5414 4776 5466
rect 4776 5414 4788 5466
rect 4788 5414 4802 5466
rect 4826 5414 4840 5466
rect 4840 5414 4852 5466
rect 4852 5414 4882 5466
rect 4906 5414 4916 5466
rect 4916 5414 4962 5466
rect 4666 5412 4722 5414
rect 4746 5412 4802 5414
rect 4826 5412 4882 5414
rect 4906 5412 4962 5414
rect 6216 7098 6272 7100
rect 6296 7098 6352 7100
rect 6376 7098 6432 7100
rect 6456 7098 6512 7100
rect 6216 7046 6262 7098
rect 6262 7046 6272 7098
rect 6296 7046 6326 7098
rect 6326 7046 6338 7098
rect 6338 7046 6352 7098
rect 6376 7046 6390 7098
rect 6390 7046 6402 7098
rect 6402 7046 6432 7098
rect 6456 7046 6466 7098
rect 6466 7046 6512 7098
rect 6216 7044 6272 7046
rect 6296 7044 6352 7046
rect 6376 7044 6432 7046
rect 6456 7044 6512 7046
rect 6216 6010 6272 6012
rect 6296 6010 6352 6012
rect 6376 6010 6432 6012
rect 6456 6010 6512 6012
rect 6216 5958 6262 6010
rect 6262 5958 6272 6010
rect 6296 5958 6326 6010
rect 6326 5958 6338 6010
rect 6338 5958 6352 6010
rect 6376 5958 6390 6010
rect 6390 5958 6402 6010
rect 6402 5958 6432 6010
rect 6456 5958 6466 6010
rect 6466 5958 6512 6010
rect 6216 5956 6272 5958
rect 6296 5956 6352 5958
rect 6376 5956 6432 5958
rect 6456 5956 6512 5958
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 3276 3834 3332 3836
rect 3356 3834 3412 3836
rect 3116 3782 3162 3834
rect 3162 3782 3172 3834
rect 3196 3782 3226 3834
rect 3226 3782 3238 3834
rect 3238 3782 3252 3834
rect 3276 3782 3290 3834
rect 3290 3782 3302 3834
rect 3302 3782 3332 3834
rect 3356 3782 3366 3834
rect 3366 3782 3412 3834
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 3276 3780 3332 3782
rect 3356 3780 3412 3782
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 3276 2746 3332 2748
rect 3356 2746 3412 2748
rect 3116 2694 3162 2746
rect 3162 2694 3172 2746
rect 3196 2694 3226 2746
rect 3226 2694 3238 2746
rect 3238 2694 3252 2746
rect 3276 2694 3290 2746
rect 3290 2694 3302 2746
rect 3302 2694 3332 2746
rect 3356 2694 3366 2746
rect 3366 2694 3412 2746
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 3276 2692 3332 2694
rect 3356 2692 3412 2694
rect 4666 4378 4722 4380
rect 4746 4378 4802 4380
rect 4826 4378 4882 4380
rect 4906 4378 4962 4380
rect 4666 4326 4712 4378
rect 4712 4326 4722 4378
rect 4746 4326 4776 4378
rect 4776 4326 4788 4378
rect 4788 4326 4802 4378
rect 4826 4326 4840 4378
rect 4840 4326 4852 4378
rect 4852 4326 4882 4378
rect 4906 4326 4916 4378
rect 4916 4326 4962 4378
rect 4666 4324 4722 4326
rect 4746 4324 4802 4326
rect 4826 4324 4882 4326
rect 4906 4324 4962 4326
rect 4666 3290 4722 3292
rect 4746 3290 4802 3292
rect 4826 3290 4882 3292
rect 4906 3290 4962 3292
rect 4666 3238 4712 3290
rect 4712 3238 4722 3290
rect 4746 3238 4776 3290
rect 4776 3238 4788 3290
rect 4788 3238 4802 3290
rect 4826 3238 4840 3290
rect 4840 3238 4852 3290
rect 4852 3238 4882 3290
rect 4906 3238 4916 3290
rect 4916 3238 4962 3290
rect 4666 3236 4722 3238
rect 4746 3236 4802 3238
rect 4826 3236 4882 3238
rect 4906 3236 4962 3238
rect 4666 2202 4722 2204
rect 4746 2202 4802 2204
rect 4826 2202 4882 2204
rect 4906 2202 4962 2204
rect 4666 2150 4712 2202
rect 4712 2150 4722 2202
rect 4746 2150 4776 2202
rect 4776 2150 4788 2202
rect 4788 2150 4802 2202
rect 4826 2150 4840 2202
rect 4840 2150 4852 2202
rect 4852 2150 4882 2202
rect 4906 2150 4916 2202
rect 4916 2150 4962 2202
rect 4666 2148 4722 2150
rect 4746 2148 4802 2150
rect 4826 2148 4882 2150
rect 4906 2148 4962 2150
rect 3116 1658 3172 1660
rect 3196 1658 3252 1660
rect 3276 1658 3332 1660
rect 3356 1658 3412 1660
rect 3116 1606 3162 1658
rect 3162 1606 3172 1658
rect 3196 1606 3226 1658
rect 3226 1606 3238 1658
rect 3238 1606 3252 1658
rect 3276 1606 3290 1658
rect 3290 1606 3302 1658
rect 3302 1606 3332 1658
rect 3356 1606 3366 1658
rect 3366 1606 3412 1658
rect 3116 1604 3172 1606
rect 3196 1604 3252 1606
rect 3276 1604 3332 1606
rect 3356 1604 3412 1606
rect 3116 570 3172 572
rect 3196 570 3252 572
rect 3276 570 3332 572
rect 3356 570 3412 572
rect 3116 518 3162 570
rect 3162 518 3172 570
rect 3196 518 3226 570
rect 3226 518 3238 570
rect 3238 518 3252 570
rect 3276 518 3290 570
rect 3290 518 3302 570
rect 3302 518 3332 570
rect 3356 518 3366 570
rect 3366 518 3412 570
rect 3116 516 3172 518
rect 3196 516 3252 518
rect 3276 516 3332 518
rect 3356 516 3412 518
rect 4666 1114 4722 1116
rect 4746 1114 4802 1116
rect 4826 1114 4882 1116
rect 4906 1114 4962 1116
rect 4666 1062 4712 1114
rect 4712 1062 4722 1114
rect 4746 1062 4776 1114
rect 4776 1062 4788 1114
rect 4788 1062 4802 1114
rect 4826 1062 4840 1114
rect 4840 1062 4852 1114
rect 4852 1062 4882 1114
rect 4906 1062 4916 1114
rect 4916 1062 4962 1114
rect 4666 1060 4722 1062
rect 4746 1060 4802 1062
rect 4826 1060 4882 1062
rect 4906 1060 4962 1062
rect 6216 4922 6272 4924
rect 6296 4922 6352 4924
rect 6376 4922 6432 4924
rect 6456 4922 6512 4924
rect 6216 4870 6262 4922
rect 6262 4870 6272 4922
rect 6296 4870 6326 4922
rect 6326 4870 6338 4922
rect 6338 4870 6352 4922
rect 6376 4870 6390 4922
rect 6390 4870 6402 4922
rect 6402 4870 6432 4922
rect 6456 4870 6466 4922
rect 6466 4870 6512 4922
rect 6216 4868 6272 4870
rect 6296 4868 6352 4870
rect 6376 4868 6432 4870
rect 6456 4868 6512 4870
rect 7766 9818 7822 9820
rect 7846 9818 7902 9820
rect 7926 9818 7982 9820
rect 8006 9818 8062 9820
rect 7766 9766 7812 9818
rect 7812 9766 7822 9818
rect 7846 9766 7876 9818
rect 7876 9766 7888 9818
rect 7888 9766 7902 9818
rect 7926 9766 7940 9818
rect 7940 9766 7952 9818
rect 7952 9766 7982 9818
rect 8006 9766 8016 9818
rect 8016 9766 8062 9818
rect 7766 9764 7822 9766
rect 7846 9764 7902 9766
rect 7926 9764 7982 9766
rect 8006 9764 8062 9766
rect 7766 8730 7822 8732
rect 7846 8730 7902 8732
rect 7926 8730 7982 8732
rect 8006 8730 8062 8732
rect 7766 8678 7812 8730
rect 7812 8678 7822 8730
rect 7846 8678 7876 8730
rect 7876 8678 7888 8730
rect 7888 8678 7902 8730
rect 7926 8678 7940 8730
rect 7940 8678 7952 8730
rect 7952 8678 7982 8730
rect 8006 8678 8016 8730
rect 8016 8678 8062 8730
rect 7766 8676 7822 8678
rect 7846 8676 7902 8678
rect 7926 8676 7982 8678
rect 8006 8676 8062 8678
rect 7766 7642 7822 7644
rect 7846 7642 7902 7644
rect 7926 7642 7982 7644
rect 8006 7642 8062 7644
rect 7766 7590 7812 7642
rect 7812 7590 7822 7642
rect 7846 7590 7876 7642
rect 7876 7590 7888 7642
rect 7888 7590 7902 7642
rect 7926 7590 7940 7642
rect 7940 7590 7952 7642
rect 7952 7590 7982 7642
rect 8006 7590 8016 7642
rect 8016 7590 8062 7642
rect 7766 7588 7822 7590
rect 7846 7588 7902 7590
rect 7926 7588 7982 7590
rect 8006 7588 8062 7590
rect 7766 6554 7822 6556
rect 7846 6554 7902 6556
rect 7926 6554 7982 6556
rect 8006 6554 8062 6556
rect 7766 6502 7812 6554
rect 7812 6502 7822 6554
rect 7846 6502 7876 6554
rect 7876 6502 7888 6554
rect 7888 6502 7902 6554
rect 7926 6502 7940 6554
rect 7940 6502 7952 6554
rect 7952 6502 7982 6554
rect 8006 6502 8016 6554
rect 8016 6502 8062 6554
rect 7766 6500 7822 6502
rect 7846 6500 7902 6502
rect 7926 6500 7982 6502
rect 8006 6500 8062 6502
rect 9316 10362 9372 10364
rect 9396 10362 9452 10364
rect 9476 10362 9532 10364
rect 9556 10362 9612 10364
rect 9316 10310 9362 10362
rect 9362 10310 9372 10362
rect 9396 10310 9426 10362
rect 9426 10310 9438 10362
rect 9438 10310 9452 10362
rect 9476 10310 9490 10362
rect 9490 10310 9502 10362
rect 9502 10310 9532 10362
rect 9556 10310 9566 10362
rect 9566 10310 9612 10362
rect 9316 10308 9372 10310
rect 9396 10308 9452 10310
rect 9476 10308 9532 10310
rect 9556 10308 9612 10310
rect 7766 5466 7822 5468
rect 7846 5466 7902 5468
rect 7926 5466 7982 5468
rect 8006 5466 8062 5468
rect 7766 5414 7812 5466
rect 7812 5414 7822 5466
rect 7846 5414 7876 5466
rect 7876 5414 7888 5466
rect 7888 5414 7902 5466
rect 7926 5414 7940 5466
rect 7940 5414 7952 5466
rect 7952 5414 7982 5466
rect 8006 5414 8016 5466
rect 8016 5414 8062 5466
rect 7766 5412 7822 5414
rect 7846 5412 7902 5414
rect 7926 5412 7982 5414
rect 8006 5412 8062 5414
rect 6216 3834 6272 3836
rect 6296 3834 6352 3836
rect 6376 3834 6432 3836
rect 6456 3834 6512 3836
rect 6216 3782 6262 3834
rect 6262 3782 6272 3834
rect 6296 3782 6326 3834
rect 6326 3782 6338 3834
rect 6338 3782 6352 3834
rect 6376 3782 6390 3834
rect 6390 3782 6402 3834
rect 6402 3782 6432 3834
rect 6456 3782 6466 3834
rect 6466 3782 6512 3834
rect 6216 3780 6272 3782
rect 6296 3780 6352 3782
rect 6376 3780 6432 3782
rect 6456 3780 6512 3782
rect 6216 2746 6272 2748
rect 6296 2746 6352 2748
rect 6376 2746 6432 2748
rect 6456 2746 6512 2748
rect 6216 2694 6262 2746
rect 6262 2694 6272 2746
rect 6296 2694 6326 2746
rect 6326 2694 6338 2746
rect 6338 2694 6352 2746
rect 6376 2694 6390 2746
rect 6390 2694 6402 2746
rect 6402 2694 6432 2746
rect 6456 2694 6466 2746
rect 6466 2694 6512 2746
rect 6216 2692 6272 2694
rect 6296 2692 6352 2694
rect 6376 2692 6432 2694
rect 6456 2692 6512 2694
rect 6216 1658 6272 1660
rect 6296 1658 6352 1660
rect 6376 1658 6432 1660
rect 6456 1658 6512 1660
rect 6216 1606 6262 1658
rect 6262 1606 6272 1658
rect 6296 1606 6326 1658
rect 6326 1606 6338 1658
rect 6338 1606 6352 1658
rect 6376 1606 6390 1658
rect 6390 1606 6402 1658
rect 6402 1606 6432 1658
rect 6456 1606 6466 1658
rect 6466 1606 6512 1658
rect 6216 1604 6272 1606
rect 6296 1604 6352 1606
rect 6376 1604 6432 1606
rect 6456 1604 6512 1606
rect 7766 4378 7822 4380
rect 7846 4378 7902 4380
rect 7926 4378 7982 4380
rect 8006 4378 8062 4380
rect 7766 4326 7812 4378
rect 7812 4326 7822 4378
rect 7846 4326 7876 4378
rect 7876 4326 7888 4378
rect 7888 4326 7902 4378
rect 7926 4326 7940 4378
rect 7940 4326 7952 4378
rect 7952 4326 7982 4378
rect 8006 4326 8016 4378
rect 8016 4326 8062 4378
rect 7766 4324 7822 4326
rect 7846 4324 7902 4326
rect 7926 4324 7982 4326
rect 8006 4324 8062 4326
rect 7766 3290 7822 3292
rect 7846 3290 7902 3292
rect 7926 3290 7982 3292
rect 8006 3290 8062 3292
rect 7766 3238 7812 3290
rect 7812 3238 7822 3290
rect 7846 3238 7876 3290
rect 7876 3238 7888 3290
rect 7888 3238 7902 3290
rect 7926 3238 7940 3290
rect 7940 3238 7952 3290
rect 7952 3238 7982 3290
rect 8006 3238 8016 3290
rect 8016 3238 8062 3290
rect 7766 3236 7822 3238
rect 7846 3236 7902 3238
rect 7926 3236 7982 3238
rect 8006 3236 8062 3238
rect 6216 570 6272 572
rect 6296 570 6352 572
rect 6376 570 6432 572
rect 6456 570 6512 572
rect 6216 518 6262 570
rect 6262 518 6272 570
rect 6296 518 6326 570
rect 6326 518 6338 570
rect 6338 518 6352 570
rect 6376 518 6390 570
rect 6390 518 6402 570
rect 6402 518 6432 570
rect 6456 518 6466 570
rect 6466 518 6512 570
rect 6216 516 6272 518
rect 6296 516 6352 518
rect 6376 516 6432 518
rect 6456 516 6512 518
rect 7766 2202 7822 2204
rect 7846 2202 7902 2204
rect 7926 2202 7982 2204
rect 8006 2202 8062 2204
rect 7766 2150 7812 2202
rect 7812 2150 7822 2202
rect 7846 2150 7876 2202
rect 7876 2150 7888 2202
rect 7888 2150 7902 2202
rect 7926 2150 7940 2202
rect 7940 2150 7952 2202
rect 7952 2150 7982 2202
rect 8006 2150 8016 2202
rect 8016 2150 8062 2202
rect 7766 2148 7822 2150
rect 7846 2148 7902 2150
rect 7926 2148 7982 2150
rect 8006 2148 8062 2150
rect 8022 1944 8078 2000
rect 7194 1536 7250 1592
rect 9316 9274 9372 9276
rect 9396 9274 9452 9276
rect 9476 9274 9532 9276
rect 9556 9274 9612 9276
rect 9316 9222 9362 9274
rect 9362 9222 9372 9274
rect 9396 9222 9426 9274
rect 9426 9222 9438 9274
rect 9438 9222 9452 9274
rect 9476 9222 9490 9274
rect 9490 9222 9502 9274
rect 9502 9222 9532 9274
rect 9556 9222 9566 9274
rect 9566 9222 9612 9274
rect 9316 9220 9372 9222
rect 9396 9220 9452 9222
rect 9476 9220 9532 9222
rect 9556 9220 9612 9222
rect 9316 8186 9372 8188
rect 9396 8186 9452 8188
rect 9476 8186 9532 8188
rect 9556 8186 9612 8188
rect 9316 8134 9362 8186
rect 9362 8134 9372 8186
rect 9396 8134 9426 8186
rect 9426 8134 9438 8186
rect 9438 8134 9452 8186
rect 9476 8134 9490 8186
rect 9490 8134 9502 8186
rect 9502 8134 9532 8186
rect 9556 8134 9566 8186
rect 9566 8134 9612 8186
rect 9316 8132 9372 8134
rect 9396 8132 9452 8134
rect 9476 8132 9532 8134
rect 9556 8132 9612 8134
rect 10866 9818 10922 9820
rect 10946 9818 11002 9820
rect 11026 9818 11082 9820
rect 11106 9818 11162 9820
rect 10866 9766 10912 9818
rect 10912 9766 10922 9818
rect 10946 9766 10976 9818
rect 10976 9766 10988 9818
rect 10988 9766 11002 9818
rect 11026 9766 11040 9818
rect 11040 9766 11052 9818
rect 11052 9766 11082 9818
rect 11106 9766 11116 9818
rect 11116 9766 11162 9818
rect 10866 9764 10922 9766
rect 10946 9764 11002 9766
rect 11026 9764 11082 9766
rect 11106 9764 11162 9766
rect 10866 8730 10922 8732
rect 10946 8730 11002 8732
rect 11026 8730 11082 8732
rect 11106 8730 11162 8732
rect 10866 8678 10912 8730
rect 10912 8678 10922 8730
rect 10946 8678 10976 8730
rect 10976 8678 10988 8730
rect 10988 8678 11002 8730
rect 11026 8678 11040 8730
rect 11040 8678 11052 8730
rect 11052 8678 11082 8730
rect 11106 8678 11116 8730
rect 11116 8678 11162 8730
rect 10866 8676 10922 8678
rect 10946 8676 11002 8678
rect 11026 8676 11082 8678
rect 11106 8676 11162 8678
rect 12416 10362 12472 10364
rect 12496 10362 12552 10364
rect 12576 10362 12632 10364
rect 12656 10362 12712 10364
rect 12416 10310 12462 10362
rect 12462 10310 12472 10362
rect 12496 10310 12526 10362
rect 12526 10310 12538 10362
rect 12538 10310 12552 10362
rect 12576 10310 12590 10362
rect 12590 10310 12602 10362
rect 12602 10310 12632 10362
rect 12656 10310 12666 10362
rect 12666 10310 12712 10362
rect 12416 10308 12472 10310
rect 12496 10308 12552 10310
rect 12576 10308 12632 10310
rect 12656 10308 12712 10310
rect 10866 7642 10922 7644
rect 10946 7642 11002 7644
rect 11026 7642 11082 7644
rect 11106 7642 11162 7644
rect 10866 7590 10912 7642
rect 10912 7590 10922 7642
rect 10946 7590 10976 7642
rect 10976 7590 10988 7642
rect 10988 7590 11002 7642
rect 11026 7590 11040 7642
rect 11040 7590 11052 7642
rect 11052 7590 11082 7642
rect 11106 7590 11116 7642
rect 11116 7590 11162 7642
rect 10866 7588 10922 7590
rect 10946 7588 11002 7590
rect 11026 7588 11082 7590
rect 11106 7588 11162 7590
rect 9316 7098 9372 7100
rect 9396 7098 9452 7100
rect 9476 7098 9532 7100
rect 9556 7098 9612 7100
rect 9316 7046 9362 7098
rect 9362 7046 9372 7098
rect 9396 7046 9426 7098
rect 9426 7046 9438 7098
rect 9438 7046 9452 7098
rect 9476 7046 9490 7098
rect 9490 7046 9502 7098
rect 9502 7046 9532 7098
rect 9556 7046 9566 7098
rect 9566 7046 9612 7098
rect 9316 7044 9372 7046
rect 9396 7044 9452 7046
rect 9476 7044 9532 7046
rect 9556 7044 9612 7046
rect 9316 6010 9372 6012
rect 9396 6010 9452 6012
rect 9476 6010 9532 6012
rect 9556 6010 9612 6012
rect 9316 5958 9362 6010
rect 9362 5958 9372 6010
rect 9396 5958 9426 6010
rect 9426 5958 9438 6010
rect 9438 5958 9452 6010
rect 9476 5958 9490 6010
rect 9490 5958 9502 6010
rect 9502 5958 9532 6010
rect 9556 5958 9566 6010
rect 9566 5958 9612 6010
rect 9316 5956 9372 5958
rect 9396 5956 9452 5958
rect 9476 5956 9532 5958
rect 9556 5956 9612 5958
rect 10866 6554 10922 6556
rect 10946 6554 11002 6556
rect 11026 6554 11082 6556
rect 11106 6554 11162 6556
rect 10866 6502 10912 6554
rect 10912 6502 10922 6554
rect 10946 6502 10976 6554
rect 10976 6502 10988 6554
rect 10988 6502 11002 6554
rect 11026 6502 11040 6554
rect 11040 6502 11052 6554
rect 11052 6502 11082 6554
rect 11106 6502 11116 6554
rect 11116 6502 11162 6554
rect 10866 6500 10922 6502
rect 10946 6500 11002 6502
rect 11026 6500 11082 6502
rect 11106 6500 11162 6502
rect 10866 5466 10922 5468
rect 10946 5466 11002 5468
rect 11026 5466 11082 5468
rect 11106 5466 11162 5468
rect 10866 5414 10912 5466
rect 10912 5414 10922 5466
rect 10946 5414 10976 5466
rect 10976 5414 10988 5466
rect 10988 5414 11002 5466
rect 11026 5414 11040 5466
rect 11040 5414 11052 5466
rect 11052 5414 11082 5466
rect 11106 5414 11116 5466
rect 11116 5414 11162 5466
rect 10866 5412 10922 5414
rect 10946 5412 11002 5414
rect 11026 5412 11082 5414
rect 11106 5412 11162 5414
rect 9316 4922 9372 4924
rect 9396 4922 9452 4924
rect 9476 4922 9532 4924
rect 9556 4922 9612 4924
rect 9316 4870 9362 4922
rect 9362 4870 9372 4922
rect 9396 4870 9426 4922
rect 9426 4870 9438 4922
rect 9438 4870 9452 4922
rect 9476 4870 9490 4922
rect 9490 4870 9502 4922
rect 9502 4870 9532 4922
rect 9556 4870 9566 4922
rect 9566 4870 9612 4922
rect 9316 4868 9372 4870
rect 9396 4868 9452 4870
rect 9476 4868 9532 4870
rect 9556 4868 9612 4870
rect 12416 9274 12472 9276
rect 12496 9274 12552 9276
rect 12576 9274 12632 9276
rect 12656 9274 12712 9276
rect 12416 9222 12462 9274
rect 12462 9222 12472 9274
rect 12496 9222 12526 9274
rect 12526 9222 12538 9274
rect 12538 9222 12552 9274
rect 12576 9222 12590 9274
rect 12590 9222 12602 9274
rect 12602 9222 12632 9274
rect 12656 9222 12666 9274
rect 12666 9222 12712 9274
rect 12416 9220 12472 9222
rect 12496 9220 12552 9222
rect 12576 9220 12632 9222
rect 12656 9220 12712 9222
rect 12416 8186 12472 8188
rect 12496 8186 12552 8188
rect 12576 8186 12632 8188
rect 12656 8186 12712 8188
rect 12416 8134 12462 8186
rect 12462 8134 12472 8186
rect 12496 8134 12526 8186
rect 12526 8134 12538 8186
rect 12538 8134 12552 8186
rect 12576 8134 12590 8186
rect 12590 8134 12602 8186
rect 12602 8134 12632 8186
rect 12656 8134 12666 8186
rect 12666 8134 12712 8186
rect 12416 8132 12472 8134
rect 12496 8132 12552 8134
rect 12576 8132 12632 8134
rect 12656 8132 12712 8134
rect 12416 7098 12472 7100
rect 12496 7098 12552 7100
rect 12576 7098 12632 7100
rect 12656 7098 12712 7100
rect 12416 7046 12462 7098
rect 12462 7046 12472 7098
rect 12496 7046 12526 7098
rect 12526 7046 12538 7098
rect 12538 7046 12552 7098
rect 12576 7046 12590 7098
rect 12590 7046 12602 7098
rect 12602 7046 12632 7098
rect 12656 7046 12666 7098
rect 12666 7046 12712 7098
rect 12416 7044 12472 7046
rect 12496 7044 12552 7046
rect 12576 7044 12632 7046
rect 12656 7044 12712 7046
rect 12416 6010 12472 6012
rect 12496 6010 12552 6012
rect 12576 6010 12632 6012
rect 12656 6010 12712 6012
rect 12416 5958 12462 6010
rect 12462 5958 12472 6010
rect 12496 5958 12526 6010
rect 12526 5958 12538 6010
rect 12538 5958 12552 6010
rect 12576 5958 12590 6010
rect 12590 5958 12602 6010
rect 12602 5958 12632 6010
rect 12656 5958 12666 6010
rect 12666 5958 12712 6010
rect 12416 5956 12472 5958
rect 12496 5956 12552 5958
rect 12576 5956 12632 5958
rect 12656 5956 12712 5958
rect 10866 4378 10922 4380
rect 10946 4378 11002 4380
rect 11026 4378 11082 4380
rect 11106 4378 11162 4380
rect 10866 4326 10912 4378
rect 10912 4326 10922 4378
rect 10946 4326 10976 4378
rect 10976 4326 10988 4378
rect 10988 4326 11002 4378
rect 11026 4326 11040 4378
rect 11040 4326 11052 4378
rect 11052 4326 11082 4378
rect 11106 4326 11116 4378
rect 11116 4326 11162 4378
rect 10866 4324 10922 4326
rect 10946 4324 11002 4326
rect 11026 4324 11082 4326
rect 11106 4324 11162 4326
rect 9316 3834 9372 3836
rect 9396 3834 9452 3836
rect 9476 3834 9532 3836
rect 9556 3834 9612 3836
rect 9316 3782 9362 3834
rect 9362 3782 9372 3834
rect 9396 3782 9426 3834
rect 9426 3782 9438 3834
rect 9438 3782 9452 3834
rect 9476 3782 9490 3834
rect 9490 3782 9502 3834
rect 9502 3782 9532 3834
rect 9556 3782 9566 3834
rect 9566 3782 9612 3834
rect 9316 3780 9372 3782
rect 9396 3780 9452 3782
rect 9476 3780 9532 3782
rect 9556 3780 9612 3782
rect 7766 1114 7822 1116
rect 7846 1114 7902 1116
rect 7926 1114 7982 1116
rect 8006 1114 8062 1116
rect 7766 1062 7812 1114
rect 7812 1062 7822 1114
rect 7846 1062 7876 1114
rect 7876 1062 7888 1114
rect 7888 1062 7902 1114
rect 7926 1062 7940 1114
rect 7940 1062 7952 1114
rect 7952 1062 7982 1114
rect 8006 1062 8016 1114
rect 8016 1062 8062 1114
rect 7766 1060 7822 1062
rect 7846 1060 7902 1062
rect 7926 1060 7982 1062
rect 8006 1060 8062 1062
rect 10866 3290 10922 3292
rect 10946 3290 11002 3292
rect 11026 3290 11082 3292
rect 11106 3290 11162 3292
rect 10866 3238 10912 3290
rect 10912 3238 10922 3290
rect 10946 3238 10976 3290
rect 10976 3238 10988 3290
rect 10988 3238 11002 3290
rect 11026 3238 11040 3290
rect 11040 3238 11052 3290
rect 11052 3238 11082 3290
rect 11106 3238 11116 3290
rect 11116 3238 11162 3290
rect 10866 3236 10922 3238
rect 10946 3236 11002 3238
rect 11026 3236 11082 3238
rect 11106 3236 11162 3238
rect 9316 2746 9372 2748
rect 9396 2746 9452 2748
rect 9476 2746 9532 2748
rect 9556 2746 9612 2748
rect 9316 2694 9362 2746
rect 9362 2694 9372 2746
rect 9396 2694 9426 2746
rect 9426 2694 9438 2746
rect 9438 2694 9452 2746
rect 9476 2694 9490 2746
rect 9490 2694 9502 2746
rect 9502 2694 9532 2746
rect 9556 2694 9566 2746
rect 9566 2694 9612 2746
rect 9316 2692 9372 2694
rect 9396 2692 9452 2694
rect 9476 2692 9532 2694
rect 9556 2692 9612 2694
rect 9402 1980 9404 2000
rect 9404 1980 9456 2000
rect 9456 1980 9458 2000
rect 9402 1944 9458 1980
rect 9316 1658 9372 1660
rect 9396 1658 9452 1660
rect 9476 1658 9532 1660
rect 9556 1658 9612 1660
rect 9316 1606 9362 1658
rect 9362 1606 9372 1658
rect 9396 1606 9426 1658
rect 9426 1606 9438 1658
rect 9438 1606 9452 1658
rect 9476 1606 9490 1658
rect 9490 1606 9502 1658
rect 9502 1606 9532 1658
rect 9556 1606 9566 1658
rect 9566 1606 9612 1658
rect 9316 1604 9372 1606
rect 9396 1604 9452 1606
rect 9476 1604 9532 1606
rect 9556 1604 9612 1606
rect 12416 4922 12472 4924
rect 12496 4922 12552 4924
rect 12576 4922 12632 4924
rect 12656 4922 12712 4924
rect 12416 4870 12462 4922
rect 12462 4870 12472 4922
rect 12496 4870 12526 4922
rect 12526 4870 12538 4922
rect 12538 4870 12552 4922
rect 12576 4870 12590 4922
rect 12590 4870 12602 4922
rect 12602 4870 12632 4922
rect 12656 4870 12666 4922
rect 12666 4870 12712 4922
rect 12416 4868 12472 4870
rect 12496 4868 12552 4870
rect 12576 4868 12632 4870
rect 12656 4868 12712 4870
rect 13966 9818 14022 9820
rect 14046 9818 14102 9820
rect 14126 9818 14182 9820
rect 14206 9818 14262 9820
rect 13966 9766 14012 9818
rect 14012 9766 14022 9818
rect 14046 9766 14076 9818
rect 14076 9766 14088 9818
rect 14088 9766 14102 9818
rect 14126 9766 14140 9818
rect 14140 9766 14152 9818
rect 14152 9766 14182 9818
rect 14206 9766 14216 9818
rect 14216 9766 14262 9818
rect 13966 9764 14022 9766
rect 14046 9764 14102 9766
rect 14126 9764 14182 9766
rect 14206 9764 14262 9766
rect 13966 8730 14022 8732
rect 14046 8730 14102 8732
rect 14126 8730 14182 8732
rect 14206 8730 14262 8732
rect 13966 8678 14012 8730
rect 14012 8678 14022 8730
rect 14046 8678 14076 8730
rect 14076 8678 14088 8730
rect 14088 8678 14102 8730
rect 14126 8678 14140 8730
rect 14140 8678 14152 8730
rect 14152 8678 14182 8730
rect 14206 8678 14216 8730
rect 14216 8678 14262 8730
rect 13966 8676 14022 8678
rect 14046 8676 14102 8678
rect 14126 8676 14182 8678
rect 14206 8676 14262 8678
rect 13966 7642 14022 7644
rect 14046 7642 14102 7644
rect 14126 7642 14182 7644
rect 14206 7642 14262 7644
rect 13966 7590 14012 7642
rect 14012 7590 14022 7642
rect 14046 7590 14076 7642
rect 14076 7590 14088 7642
rect 14088 7590 14102 7642
rect 14126 7590 14140 7642
rect 14140 7590 14152 7642
rect 14152 7590 14182 7642
rect 14206 7590 14216 7642
rect 14216 7590 14262 7642
rect 13966 7588 14022 7590
rect 14046 7588 14102 7590
rect 14126 7588 14182 7590
rect 14206 7588 14262 7590
rect 13966 6554 14022 6556
rect 14046 6554 14102 6556
rect 14126 6554 14182 6556
rect 14206 6554 14262 6556
rect 13966 6502 14012 6554
rect 14012 6502 14022 6554
rect 14046 6502 14076 6554
rect 14076 6502 14088 6554
rect 14088 6502 14102 6554
rect 14126 6502 14140 6554
rect 14140 6502 14152 6554
rect 14152 6502 14182 6554
rect 14206 6502 14216 6554
rect 14216 6502 14262 6554
rect 13966 6500 14022 6502
rect 14046 6500 14102 6502
rect 14126 6500 14182 6502
rect 14206 6500 14262 6502
rect 13966 5466 14022 5468
rect 14046 5466 14102 5468
rect 14126 5466 14182 5468
rect 14206 5466 14262 5468
rect 13966 5414 14012 5466
rect 14012 5414 14022 5466
rect 14046 5414 14076 5466
rect 14076 5414 14088 5466
rect 14088 5414 14102 5466
rect 14126 5414 14140 5466
rect 14140 5414 14152 5466
rect 14152 5414 14182 5466
rect 14206 5414 14216 5466
rect 14216 5414 14262 5466
rect 13966 5412 14022 5414
rect 14046 5412 14102 5414
rect 14126 5412 14182 5414
rect 14206 5412 14262 5414
rect 12416 3834 12472 3836
rect 12496 3834 12552 3836
rect 12576 3834 12632 3836
rect 12656 3834 12712 3836
rect 12416 3782 12462 3834
rect 12462 3782 12472 3834
rect 12496 3782 12526 3834
rect 12526 3782 12538 3834
rect 12538 3782 12552 3834
rect 12576 3782 12590 3834
rect 12590 3782 12602 3834
rect 12602 3782 12632 3834
rect 12656 3782 12666 3834
rect 12666 3782 12712 3834
rect 12416 3780 12472 3782
rect 12496 3780 12552 3782
rect 12576 3780 12632 3782
rect 12656 3780 12712 3782
rect 17066 10906 17122 10908
rect 17146 10906 17202 10908
rect 17226 10906 17282 10908
rect 17306 10906 17362 10908
rect 17066 10854 17112 10906
rect 17112 10854 17122 10906
rect 17146 10854 17176 10906
rect 17176 10854 17188 10906
rect 17188 10854 17202 10906
rect 17226 10854 17240 10906
rect 17240 10854 17252 10906
rect 17252 10854 17282 10906
rect 17306 10854 17316 10906
rect 17316 10854 17362 10906
rect 17066 10852 17122 10854
rect 17146 10852 17202 10854
rect 17226 10852 17282 10854
rect 17306 10852 17362 10854
rect 15516 10362 15572 10364
rect 15596 10362 15652 10364
rect 15676 10362 15732 10364
rect 15756 10362 15812 10364
rect 15516 10310 15562 10362
rect 15562 10310 15572 10362
rect 15596 10310 15626 10362
rect 15626 10310 15638 10362
rect 15638 10310 15652 10362
rect 15676 10310 15690 10362
rect 15690 10310 15702 10362
rect 15702 10310 15732 10362
rect 15756 10310 15766 10362
rect 15766 10310 15812 10362
rect 15516 10308 15572 10310
rect 15596 10308 15652 10310
rect 15676 10308 15732 10310
rect 15756 10308 15812 10310
rect 17066 9818 17122 9820
rect 17146 9818 17202 9820
rect 17226 9818 17282 9820
rect 17306 9818 17362 9820
rect 17066 9766 17112 9818
rect 17112 9766 17122 9818
rect 17146 9766 17176 9818
rect 17176 9766 17188 9818
rect 17188 9766 17202 9818
rect 17226 9766 17240 9818
rect 17240 9766 17252 9818
rect 17252 9766 17282 9818
rect 17306 9766 17316 9818
rect 17316 9766 17362 9818
rect 17066 9764 17122 9766
rect 17146 9764 17202 9766
rect 17226 9764 17282 9766
rect 17306 9764 17362 9766
rect 15516 9274 15572 9276
rect 15596 9274 15652 9276
rect 15676 9274 15732 9276
rect 15756 9274 15812 9276
rect 15516 9222 15562 9274
rect 15562 9222 15572 9274
rect 15596 9222 15626 9274
rect 15626 9222 15638 9274
rect 15638 9222 15652 9274
rect 15676 9222 15690 9274
rect 15690 9222 15702 9274
rect 15702 9222 15732 9274
rect 15756 9222 15766 9274
rect 15766 9222 15812 9274
rect 15516 9220 15572 9222
rect 15596 9220 15652 9222
rect 15676 9220 15732 9222
rect 15756 9220 15812 9222
rect 15516 8186 15572 8188
rect 15596 8186 15652 8188
rect 15676 8186 15732 8188
rect 15756 8186 15812 8188
rect 15516 8134 15562 8186
rect 15562 8134 15572 8186
rect 15596 8134 15626 8186
rect 15626 8134 15638 8186
rect 15638 8134 15652 8186
rect 15676 8134 15690 8186
rect 15690 8134 15702 8186
rect 15702 8134 15732 8186
rect 15756 8134 15766 8186
rect 15766 8134 15812 8186
rect 15516 8132 15572 8134
rect 15596 8132 15652 8134
rect 15676 8132 15732 8134
rect 15756 8132 15812 8134
rect 17066 8730 17122 8732
rect 17146 8730 17202 8732
rect 17226 8730 17282 8732
rect 17306 8730 17362 8732
rect 17066 8678 17112 8730
rect 17112 8678 17122 8730
rect 17146 8678 17176 8730
rect 17176 8678 17188 8730
rect 17188 8678 17202 8730
rect 17226 8678 17240 8730
rect 17240 8678 17252 8730
rect 17252 8678 17282 8730
rect 17306 8678 17316 8730
rect 17316 8678 17362 8730
rect 17066 8676 17122 8678
rect 17146 8676 17202 8678
rect 17226 8676 17282 8678
rect 17306 8676 17362 8678
rect 15516 7098 15572 7100
rect 15596 7098 15652 7100
rect 15676 7098 15732 7100
rect 15756 7098 15812 7100
rect 15516 7046 15562 7098
rect 15562 7046 15572 7098
rect 15596 7046 15626 7098
rect 15626 7046 15638 7098
rect 15638 7046 15652 7098
rect 15676 7046 15690 7098
rect 15690 7046 15702 7098
rect 15702 7046 15732 7098
rect 15756 7046 15766 7098
rect 15766 7046 15812 7098
rect 15516 7044 15572 7046
rect 15596 7044 15652 7046
rect 15676 7044 15732 7046
rect 15756 7044 15812 7046
rect 18786 11192 18842 11248
rect 18602 9696 18658 9752
rect 18602 8200 18658 8256
rect 17066 7642 17122 7644
rect 17146 7642 17202 7644
rect 17226 7642 17282 7644
rect 17306 7642 17362 7644
rect 17066 7590 17112 7642
rect 17112 7590 17122 7642
rect 17146 7590 17176 7642
rect 17176 7590 17188 7642
rect 17188 7590 17202 7642
rect 17226 7590 17240 7642
rect 17240 7590 17252 7642
rect 17252 7590 17282 7642
rect 17306 7590 17316 7642
rect 17316 7590 17362 7642
rect 17066 7588 17122 7590
rect 17146 7588 17202 7590
rect 17226 7588 17282 7590
rect 17306 7588 17362 7590
rect 17066 6554 17122 6556
rect 17146 6554 17202 6556
rect 17226 6554 17282 6556
rect 17306 6554 17362 6556
rect 17066 6502 17112 6554
rect 17112 6502 17122 6554
rect 17146 6502 17176 6554
rect 17176 6502 17188 6554
rect 17188 6502 17202 6554
rect 17226 6502 17240 6554
rect 17240 6502 17252 6554
rect 17252 6502 17282 6554
rect 17306 6502 17316 6554
rect 17316 6502 17362 6554
rect 17066 6500 17122 6502
rect 17146 6500 17202 6502
rect 17226 6500 17282 6502
rect 17306 6500 17362 6502
rect 15516 6010 15572 6012
rect 15596 6010 15652 6012
rect 15676 6010 15732 6012
rect 15756 6010 15812 6012
rect 15516 5958 15562 6010
rect 15562 5958 15572 6010
rect 15596 5958 15626 6010
rect 15626 5958 15638 6010
rect 15638 5958 15652 6010
rect 15676 5958 15690 6010
rect 15690 5958 15702 6010
rect 15702 5958 15732 6010
rect 15756 5958 15766 6010
rect 15766 5958 15812 6010
rect 15516 5956 15572 5958
rect 15596 5956 15652 5958
rect 15676 5956 15732 5958
rect 15756 5956 15812 5958
rect 13966 4378 14022 4380
rect 14046 4378 14102 4380
rect 14126 4378 14182 4380
rect 14206 4378 14262 4380
rect 13966 4326 14012 4378
rect 14012 4326 14022 4378
rect 14046 4326 14076 4378
rect 14076 4326 14088 4378
rect 14088 4326 14102 4378
rect 14126 4326 14140 4378
rect 14140 4326 14152 4378
rect 14152 4326 14182 4378
rect 14206 4326 14216 4378
rect 14216 4326 14262 4378
rect 13966 4324 14022 4326
rect 14046 4324 14102 4326
rect 14126 4324 14182 4326
rect 14206 4324 14262 4326
rect 12416 2746 12472 2748
rect 12496 2746 12552 2748
rect 12576 2746 12632 2748
rect 12656 2746 12712 2748
rect 12416 2694 12462 2746
rect 12462 2694 12472 2746
rect 12496 2694 12526 2746
rect 12526 2694 12538 2746
rect 12538 2694 12552 2746
rect 12576 2694 12590 2746
rect 12590 2694 12602 2746
rect 12602 2694 12632 2746
rect 12656 2694 12666 2746
rect 12666 2694 12712 2746
rect 12416 2692 12472 2694
rect 12496 2692 12552 2694
rect 12576 2692 12632 2694
rect 12656 2692 12712 2694
rect 10866 2202 10922 2204
rect 10946 2202 11002 2204
rect 11026 2202 11082 2204
rect 11106 2202 11162 2204
rect 10866 2150 10912 2202
rect 10912 2150 10922 2202
rect 10946 2150 10976 2202
rect 10976 2150 10988 2202
rect 10988 2150 11002 2202
rect 11026 2150 11040 2202
rect 11040 2150 11052 2202
rect 11052 2150 11082 2202
rect 11106 2150 11116 2202
rect 11116 2150 11162 2202
rect 10866 2148 10922 2150
rect 10946 2148 11002 2150
rect 11026 2148 11082 2150
rect 11106 2148 11162 2150
rect 10138 1944 10194 2000
rect 11150 1964 11206 2000
rect 11150 1944 11152 1964
rect 11152 1944 11204 1964
rect 11204 1944 11206 1964
rect 11242 1808 11298 1864
rect 9316 570 9372 572
rect 9396 570 9452 572
rect 9476 570 9532 572
rect 9556 570 9612 572
rect 9316 518 9362 570
rect 9362 518 9372 570
rect 9396 518 9426 570
rect 9426 518 9438 570
rect 9438 518 9452 570
rect 9476 518 9490 570
rect 9490 518 9502 570
rect 9502 518 9532 570
rect 9556 518 9566 570
rect 9566 518 9612 570
rect 9316 516 9372 518
rect 9396 516 9452 518
rect 9476 516 9532 518
rect 9556 516 9612 518
rect 10866 1114 10922 1116
rect 10946 1114 11002 1116
rect 11026 1114 11082 1116
rect 11106 1114 11162 1116
rect 10866 1062 10912 1114
rect 10912 1062 10922 1114
rect 10946 1062 10976 1114
rect 10976 1062 10988 1114
rect 10988 1062 11002 1114
rect 11026 1062 11040 1114
rect 11040 1062 11052 1114
rect 11052 1062 11082 1114
rect 11106 1062 11116 1114
rect 11116 1062 11162 1114
rect 10866 1060 10922 1062
rect 10946 1060 11002 1062
rect 11026 1060 11082 1062
rect 11106 1060 11162 1062
rect 13966 3290 14022 3292
rect 14046 3290 14102 3292
rect 14126 3290 14182 3292
rect 14206 3290 14262 3292
rect 13966 3238 14012 3290
rect 14012 3238 14022 3290
rect 14046 3238 14076 3290
rect 14076 3238 14088 3290
rect 14088 3238 14102 3290
rect 14126 3238 14140 3290
rect 14140 3238 14152 3290
rect 14152 3238 14182 3290
rect 14206 3238 14216 3290
rect 14216 3238 14262 3290
rect 13966 3236 14022 3238
rect 14046 3236 14102 3238
rect 14126 3236 14182 3238
rect 14206 3236 14262 3238
rect 12416 1658 12472 1660
rect 12496 1658 12552 1660
rect 12576 1658 12632 1660
rect 12656 1658 12712 1660
rect 12416 1606 12462 1658
rect 12462 1606 12472 1658
rect 12496 1606 12526 1658
rect 12526 1606 12538 1658
rect 12538 1606 12552 1658
rect 12576 1606 12590 1658
rect 12590 1606 12602 1658
rect 12602 1606 12632 1658
rect 12656 1606 12666 1658
rect 12666 1606 12712 1658
rect 12416 1604 12472 1606
rect 12496 1604 12552 1606
rect 12576 1604 12632 1606
rect 12656 1604 12712 1606
rect 12622 1400 12678 1456
rect 12070 1284 12126 1320
rect 12070 1264 12072 1284
rect 12072 1264 12124 1284
rect 12124 1264 12126 1284
rect 12416 570 12472 572
rect 12496 570 12552 572
rect 12576 570 12632 572
rect 12656 570 12712 572
rect 12416 518 12462 570
rect 12462 518 12472 570
rect 12496 518 12526 570
rect 12526 518 12538 570
rect 12538 518 12552 570
rect 12576 518 12590 570
rect 12590 518 12602 570
rect 12602 518 12632 570
rect 12656 518 12666 570
rect 12666 518 12712 570
rect 12416 516 12472 518
rect 12496 516 12552 518
rect 12576 516 12632 518
rect 12656 516 12712 518
rect 13542 1300 13544 1320
rect 13544 1300 13596 1320
rect 13596 1300 13598 1320
rect 13542 1264 13598 1300
rect 13966 2202 14022 2204
rect 14046 2202 14102 2204
rect 14126 2202 14182 2204
rect 14206 2202 14262 2204
rect 13966 2150 14012 2202
rect 14012 2150 14022 2202
rect 14046 2150 14076 2202
rect 14076 2150 14088 2202
rect 14088 2150 14102 2202
rect 14126 2150 14140 2202
rect 14140 2150 14152 2202
rect 14152 2150 14182 2202
rect 14206 2150 14216 2202
rect 14216 2150 14262 2202
rect 13966 2148 14022 2150
rect 14046 2148 14102 2150
rect 14126 2148 14182 2150
rect 14206 2148 14262 2150
rect 15516 4922 15572 4924
rect 15596 4922 15652 4924
rect 15676 4922 15732 4924
rect 15756 4922 15812 4924
rect 15516 4870 15562 4922
rect 15562 4870 15572 4922
rect 15596 4870 15626 4922
rect 15626 4870 15638 4922
rect 15638 4870 15652 4922
rect 15676 4870 15690 4922
rect 15690 4870 15702 4922
rect 15702 4870 15732 4922
rect 15756 4870 15766 4922
rect 15766 4870 15812 4922
rect 15516 4868 15572 4870
rect 15596 4868 15652 4870
rect 15676 4868 15732 4870
rect 15756 4868 15812 4870
rect 14738 1808 14794 1864
rect 14554 1400 14610 1456
rect 13966 1114 14022 1116
rect 14046 1114 14102 1116
rect 14126 1114 14182 1116
rect 14206 1114 14262 1116
rect 13966 1062 14012 1114
rect 14012 1062 14022 1114
rect 14046 1062 14076 1114
rect 14076 1062 14088 1114
rect 14088 1062 14102 1114
rect 14126 1062 14140 1114
rect 14140 1062 14152 1114
rect 14152 1062 14182 1114
rect 14206 1062 14216 1114
rect 14216 1062 14262 1114
rect 13966 1060 14022 1062
rect 14046 1060 14102 1062
rect 14126 1060 14182 1062
rect 14206 1060 14262 1062
rect 15516 3834 15572 3836
rect 15596 3834 15652 3836
rect 15676 3834 15732 3836
rect 15756 3834 15812 3836
rect 15516 3782 15562 3834
rect 15562 3782 15572 3834
rect 15596 3782 15626 3834
rect 15626 3782 15638 3834
rect 15638 3782 15652 3834
rect 15676 3782 15690 3834
rect 15690 3782 15702 3834
rect 15702 3782 15732 3834
rect 15756 3782 15766 3834
rect 15766 3782 15812 3834
rect 15516 3780 15572 3782
rect 15596 3780 15652 3782
rect 15676 3780 15732 3782
rect 15756 3780 15812 3782
rect 17066 5466 17122 5468
rect 17146 5466 17202 5468
rect 17226 5466 17282 5468
rect 17306 5466 17362 5468
rect 17066 5414 17112 5466
rect 17112 5414 17122 5466
rect 17146 5414 17176 5466
rect 17176 5414 17188 5466
rect 17188 5414 17202 5466
rect 17226 5414 17240 5466
rect 17240 5414 17252 5466
rect 17252 5414 17282 5466
rect 17306 5414 17316 5466
rect 17316 5414 17362 5466
rect 17066 5412 17122 5414
rect 17146 5412 17202 5414
rect 17226 5412 17282 5414
rect 17306 5412 17362 5414
rect 18510 6740 18512 6760
rect 18512 6740 18564 6760
rect 18564 6740 18566 6760
rect 18510 6704 18566 6740
rect 17066 4378 17122 4380
rect 17146 4378 17202 4380
rect 17226 4378 17282 4380
rect 17306 4378 17362 4380
rect 17066 4326 17112 4378
rect 17112 4326 17122 4378
rect 17146 4326 17176 4378
rect 17176 4326 17188 4378
rect 17188 4326 17202 4378
rect 17226 4326 17240 4378
rect 17240 4326 17252 4378
rect 17252 4326 17282 4378
rect 17306 4326 17316 4378
rect 17316 4326 17362 4378
rect 17066 4324 17122 4326
rect 17146 4324 17202 4326
rect 17226 4324 17282 4326
rect 17306 4324 17362 4326
rect 17066 3290 17122 3292
rect 17146 3290 17202 3292
rect 17226 3290 17282 3292
rect 17306 3290 17362 3292
rect 17066 3238 17112 3290
rect 17112 3238 17122 3290
rect 17146 3238 17176 3290
rect 17176 3238 17188 3290
rect 17188 3238 17202 3290
rect 17226 3238 17240 3290
rect 17240 3238 17252 3290
rect 17252 3238 17282 3290
rect 17306 3238 17316 3290
rect 17316 3238 17362 3290
rect 17066 3236 17122 3238
rect 17146 3236 17202 3238
rect 17226 3236 17282 3238
rect 17306 3236 17362 3238
rect 15516 2746 15572 2748
rect 15596 2746 15652 2748
rect 15676 2746 15732 2748
rect 15756 2746 15812 2748
rect 15516 2694 15562 2746
rect 15562 2694 15572 2746
rect 15596 2694 15626 2746
rect 15626 2694 15638 2746
rect 15638 2694 15652 2746
rect 15676 2694 15690 2746
rect 15690 2694 15702 2746
rect 15702 2694 15732 2746
rect 15756 2694 15766 2746
rect 15766 2694 15812 2746
rect 15516 2692 15572 2694
rect 15596 2692 15652 2694
rect 15676 2692 15732 2694
rect 15756 2692 15812 2694
rect 17066 2202 17122 2204
rect 17146 2202 17202 2204
rect 17226 2202 17282 2204
rect 17306 2202 17362 2204
rect 17066 2150 17112 2202
rect 17112 2150 17122 2202
rect 17146 2150 17176 2202
rect 17176 2150 17188 2202
rect 17188 2150 17202 2202
rect 17226 2150 17240 2202
rect 17240 2150 17252 2202
rect 17252 2150 17282 2202
rect 17306 2150 17316 2202
rect 17316 2150 17362 2202
rect 17066 2148 17122 2150
rect 17146 2148 17202 2150
rect 17226 2148 17282 2150
rect 17306 2148 17362 2150
rect 18510 5208 18566 5264
rect 17866 2216 17922 2272
rect 15516 1658 15572 1660
rect 15596 1658 15652 1660
rect 15676 1658 15732 1660
rect 15756 1658 15812 1660
rect 15516 1606 15562 1658
rect 15562 1606 15572 1658
rect 15596 1606 15626 1658
rect 15626 1606 15638 1658
rect 15638 1606 15652 1658
rect 15676 1606 15690 1658
rect 15690 1606 15702 1658
rect 15702 1606 15732 1658
rect 15756 1606 15766 1658
rect 15766 1606 15812 1658
rect 15516 1604 15572 1606
rect 15596 1604 15652 1606
rect 15676 1604 15732 1606
rect 15756 1604 15812 1606
rect 15516 570 15572 572
rect 15596 570 15652 572
rect 15676 570 15732 572
rect 15756 570 15812 572
rect 15516 518 15562 570
rect 15562 518 15572 570
rect 15596 518 15626 570
rect 15626 518 15638 570
rect 15638 518 15652 570
rect 15676 518 15690 570
rect 15690 518 15702 570
rect 15702 518 15732 570
rect 15756 518 15766 570
rect 15766 518 15812 570
rect 15516 516 15572 518
rect 15596 516 15652 518
rect 15676 516 15732 518
rect 15756 516 15812 518
rect 17066 1114 17122 1116
rect 17146 1114 17202 1116
rect 17226 1114 17282 1116
rect 17306 1114 17362 1116
rect 17066 1062 17112 1114
rect 17112 1062 17122 1114
rect 17146 1062 17176 1114
rect 17176 1062 17188 1114
rect 17188 1062 17202 1114
rect 17226 1062 17240 1114
rect 17240 1062 17252 1114
rect 17252 1062 17282 1114
rect 17306 1062 17316 1114
rect 17316 1062 17362 1114
rect 17066 1060 17122 1062
rect 17146 1060 17202 1062
rect 17226 1060 17282 1062
rect 17306 1060 17362 1062
rect 18510 3712 18566 3768
rect 18510 756 18512 776
rect 18512 756 18564 776
rect 18564 756 18566 776
rect 18510 720 18566 756
rect 4666 26 4722 28
rect 4746 26 4802 28
rect 4826 26 4882 28
rect 4906 26 4962 28
rect 4666 -26 4712 26
rect 4712 -26 4722 26
rect 4746 -26 4776 26
rect 4776 -26 4788 26
rect 4788 -26 4802 26
rect 4826 -26 4840 26
rect 4840 -26 4852 26
rect 4852 -26 4882 26
rect 4906 -26 4916 26
rect 4916 -26 4962 26
rect 4666 -28 4722 -26
rect 4746 -28 4802 -26
rect 4826 -28 4882 -26
rect 4906 -28 4962 -26
rect 7766 26 7822 28
rect 7846 26 7902 28
rect 7926 26 7982 28
rect 8006 26 8062 28
rect 7766 -26 7812 26
rect 7812 -26 7822 26
rect 7846 -26 7876 26
rect 7876 -26 7888 26
rect 7888 -26 7902 26
rect 7926 -26 7940 26
rect 7940 -26 7952 26
rect 7952 -26 7982 26
rect 8006 -26 8016 26
rect 8016 -26 8062 26
rect 7766 -28 7822 -26
rect 7846 -28 7902 -26
rect 7926 -28 7982 -26
rect 8006 -28 8062 -26
rect 10866 26 10922 28
rect 10946 26 11002 28
rect 11026 26 11082 28
rect 11106 26 11162 28
rect 10866 -26 10912 26
rect 10912 -26 10922 26
rect 10946 -26 10976 26
rect 10976 -26 10988 26
rect 10988 -26 11002 26
rect 11026 -26 11040 26
rect 11040 -26 11052 26
rect 11052 -26 11082 26
rect 11106 -26 11116 26
rect 11116 -26 11162 26
rect 10866 -28 10922 -26
rect 10946 -28 11002 -26
rect 11026 -28 11082 -26
rect 11106 -28 11162 -26
rect 13966 26 14022 28
rect 14046 26 14102 28
rect 14126 26 14182 28
rect 14206 26 14262 28
rect 13966 -26 14012 26
rect 14012 -26 14022 26
rect 14046 -26 14076 26
rect 14076 -26 14088 26
rect 14088 -26 14102 26
rect 14126 -26 14140 26
rect 14140 -26 14152 26
rect 14152 -26 14182 26
rect 14206 -26 14216 26
rect 14216 -26 14262 26
rect 13966 -28 14022 -26
rect 14046 -28 14102 -26
rect 14126 -28 14182 -26
rect 14206 -28 14262 -26
rect 17066 26 17122 28
rect 17146 26 17202 28
rect 17226 26 17282 28
rect 17306 26 17362 28
rect 17066 -26 17112 26
rect 17112 -26 17122 26
rect 17146 -26 17176 26
rect 17176 -26 17188 26
rect 17188 -26 17202 26
rect 17226 -26 17240 26
rect 17240 -26 17252 26
rect 17252 -26 17282 26
rect 17306 -26 17316 26
rect 17316 -26 17362 26
rect 17066 -28 17122 -26
rect 17146 -28 17202 -26
rect 17226 -28 17282 -26
rect 17306 -28 17362 -26
<< metal3 >>
rect 18781 11250 18847 11253
rect 19200 11250 20000 11280
rect 18781 11248 20000 11250
rect 18781 11192 18786 11248
rect 18842 11192 20000 11248
rect 18781 11190 20000 11192
rect 18781 11187 18847 11190
rect 19200 11160 20000 11190
rect 4654 10912 4974 10913
rect 4654 10848 4662 10912
rect 4726 10848 4742 10912
rect 4806 10848 4822 10912
rect 4886 10848 4902 10912
rect 4966 10848 4974 10912
rect 4654 10847 4974 10848
rect 7754 10912 8074 10913
rect 7754 10848 7762 10912
rect 7826 10848 7842 10912
rect 7906 10848 7922 10912
rect 7986 10848 8002 10912
rect 8066 10848 8074 10912
rect 7754 10847 8074 10848
rect 10854 10912 11174 10913
rect 10854 10848 10862 10912
rect 10926 10848 10942 10912
rect 11006 10848 11022 10912
rect 11086 10848 11102 10912
rect 11166 10848 11174 10912
rect 10854 10847 11174 10848
rect 13954 10912 14274 10913
rect 13954 10848 13962 10912
rect 14026 10848 14042 10912
rect 14106 10848 14122 10912
rect 14186 10848 14202 10912
rect 14266 10848 14274 10912
rect 13954 10847 14274 10848
rect 17054 10912 17374 10913
rect 17054 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17222 10912
rect 17286 10848 17302 10912
rect 17366 10848 17374 10912
rect 17054 10847 17374 10848
rect 3104 10368 3424 10369
rect 3104 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3272 10368
rect 3336 10304 3352 10368
rect 3416 10304 3424 10368
rect 3104 10303 3424 10304
rect 6204 10368 6524 10369
rect 6204 10304 6212 10368
rect 6276 10304 6292 10368
rect 6356 10304 6372 10368
rect 6436 10304 6452 10368
rect 6516 10304 6524 10368
rect 6204 10303 6524 10304
rect 9304 10368 9624 10369
rect 9304 10304 9312 10368
rect 9376 10304 9392 10368
rect 9456 10304 9472 10368
rect 9536 10304 9552 10368
rect 9616 10304 9624 10368
rect 9304 10303 9624 10304
rect 12404 10368 12724 10369
rect 12404 10304 12412 10368
rect 12476 10304 12492 10368
rect 12556 10304 12572 10368
rect 12636 10304 12652 10368
rect 12716 10304 12724 10368
rect 12404 10303 12724 10304
rect 15504 10368 15824 10369
rect 15504 10304 15512 10368
rect 15576 10304 15592 10368
rect 15656 10304 15672 10368
rect 15736 10304 15752 10368
rect 15816 10304 15824 10368
rect 15504 10303 15824 10304
rect 4654 9824 4974 9825
rect 4654 9760 4662 9824
rect 4726 9760 4742 9824
rect 4806 9760 4822 9824
rect 4886 9760 4902 9824
rect 4966 9760 4974 9824
rect 4654 9759 4974 9760
rect 7754 9824 8074 9825
rect 7754 9760 7762 9824
rect 7826 9760 7842 9824
rect 7906 9760 7922 9824
rect 7986 9760 8002 9824
rect 8066 9760 8074 9824
rect 7754 9759 8074 9760
rect 10854 9824 11174 9825
rect 10854 9760 10862 9824
rect 10926 9760 10942 9824
rect 11006 9760 11022 9824
rect 11086 9760 11102 9824
rect 11166 9760 11174 9824
rect 10854 9759 11174 9760
rect 13954 9824 14274 9825
rect 13954 9760 13962 9824
rect 14026 9760 14042 9824
rect 14106 9760 14122 9824
rect 14186 9760 14202 9824
rect 14266 9760 14274 9824
rect 13954 9759 14274 9760
rect 17054 9824 17374 9825
rect 17054 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17222 9824
rect 17286 9760 17302 9824
rect 17366 9760 17374 9824
rect 17054 9759 17374 9760
rect 18597 9754 18663 9757
rect 19200 9754 20000 9784
rect 18597 9752 20000 9754
rect 18597 9696 18602 9752
rect 18658 9696 20000 9752
rect 18597 9694 20000 9696
rect 18597 9691 18663 9694
rect 19200 9664 20000 9694
rect 3104 9280 3424 9281
rect 3104 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3272 9280
rect 3336 9216 3352 9280
rect 3416 9216 3424 9280
rect 3104 9215 3424 9216
rect 6204 9280 6524 9281
rect 6204 9216 6212 9280
rect 6276 9216 6292 9280
rect 6356 9216 6372 9280
rect 6436 9216 6452 9280
rect 6516 9216 6524 9280
rect 6204 9215 6524 9216
rect 9304 9280 9624 9281
rect 9304 9216 9312 9280
rect 9376 9216 9392 9280
rect 9456 9216 9472 9280
rect 9536 9216 9552 9280
rect 9616 9216 9624 9280
rect 9304 9215 9624 9216
rect 12404 9280 12724 9281
rect 12404 9216 12412 9280
rect 12476 9216 12492 9280
rect 12556 9216 12572 9280
rect 12636 9216 12652 9280
rect 12716 9216 12724 9280
rect 12404 9215 12724 9216
rect 15504 9280 15824 9281
rect 15504 9216 15512 9280
rect 15576 9216 15592 9280
rect 15656 9216 15672 9280
rect 15736 9216 15752 9280
rect 15816 9216 15824 9280
rect 15504 9215 15824 9216
rect 4654 8736 4974 8737
rect 4654 8672 4662 8736
rect 4726 8672 4742 8736
rect 4806 8672 4822 8736
rect 4886 8672 4902 8736
rect 4966 8672 4974 8736
rect 4654 8671 4974 8672
rect 7754 8736 8074 8737
rect 7754 8672 7762 8736
rect 7826 8672 7842 8736
rect 7906 8672 7922 8736
rect 7986 8672 8002 8736
rect 8066 8672 8074 8736
rect 7754 8671 8074 8672
rect 10854 8736 11174 8737
rect 10854 8672 10862 8736
rect 10926 8672 10942 8736
rect 11006 8672 11022 8736
rect 11086 8672 11102 8736
rect 11166 8672 11174 8736
rect 10854 8671 11174 8672
rect 13954 8736 14274 8737
rect 13954 8672 13962 8736
rect 14026 8672 14042 8736
rect 14106 8672 14122 8736
rect 14186 8672 14202 8736
rect 14266 8672 14274 8736
rect 13954 8671 14274 8672
rect 17054 8736 17374 8737
rect 17054 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17222 8736
rect 17286 8672 17302 8736
rect 17366 8672 17374 8736
rect 17054 8671 17374 8672
rect 18597 8258 18663 8261
rect 19200 8258 20000 8288
rect 18597 8256 20000 8258
rect 18597 8200 18602 8256
rect 18658 8200 20000 8256
rect 18597 8198 20000 8200
rect 18597 8195 18663 8198
rect 3104 8192 3424 8193
rect 3104 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3272 8192
rect 3336 8128 3352 8192
rect 3416 8128 3424 8192
rect 3104 8127 3424 8128
rect 6204 8192 6524 8193
rect 6204 8128 6212 8192
rect 6276 8128 6292 8192
rect 6356 8128 6372 8192
rect 6436 8128 6452 8192
rect 6516 8128 6524 8192
rect 6204 8127 6524 8128
rect 9304 8192 9624 8193
rect 9304 8128 9312 8192
rect 9376 8128 9392 8192
rect 9456 8128 9472 8192
rect 9536 8128 9552 8192
rect 9616 8128 9624 8192
rect 9304 8127 9624 8128
rect 12404 8192 12724 8193
rect 12404 8128 12412 8192
rect 12476 8128 12492 8192
rect 12556 8128 12572 8192
rect 12636 8128 12652 8192
rect 12716 8128 12724 8192
rect 12404 8127 12724 8128
rect 15504 8192 15824 8193
rect 15504 8128 15512 8192
rect 15576 8128 15592 8192
rect 15656 8128 15672 8192
rect 15736 8128 15752 8192
rect 15816 8128 15824 8192
rect 19200 8168 20000 8198
rect 15504 8127 15824 8128
rect 4654 7648 4974 7649
rect 4654 7584 4662 7648
rect 4726 7584 4742 7648
rect 4806 7584 4822 7648
rect 4886 7584 4902 7648
rect 4966 7584 4974 7648
rect 4654 7583 4974 7584
rect 7754 7648 8074 7649
rect 7754 7584 7762 7648
rect 7826 7584 7842 7648
rect 7906 7584 7922 7648
rect 7986 7584 8002 7648
rect 8066 7584 8074 7648
rect 7754 7583 8074 7584
rect 10854 7648 11174 7649
rect 10854 7584 10862 7648
rect 10926 7584 10942 7648
rect 11006 7584 11022 7648
rect 11086 7584 11102 7648
rect 11166 7584 11174 7648
rect 10854 7583 11174 7584
rect 13954 7648 14274 7649
rect 13954 7584 13962 7648
rect 14026 7584 14042 7648
rect 14106 7584 14122 7648
rect 14186 7584 14202 7648
rect 14266 7584 14274 7648
rect 13954 7583 14274 7584
rect 17054 7648 17374 7649
rect 17054 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17222 7648
rect 17286 7584 17302 7648
rect 17366 7584 17374 7648
rect 17054 7583 17374 7584
rect 3785 7442 3851 7445
rect 4797 7442 4863 7445
rect 3785 7440 4863 7442
rect 3785 7384 3790 7440
rect 3846 7384 4802 7440
rect 4858 7384 4863 7440
rect 3785 7382 4863 7384
rect 3785 7379 3851 7382
rect 4797 7379 4863 7382
rect 3104 7104 3424 7105
rect 3104 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3272 7104
rect 3336 7040 3352 7104
rect 3416 7040 3424 7104
rect 3104 7039 3424 7040
rect 6204 7104 6524 7105
rect 6204 7040 6212 7104
rect 6276 7040 6292 7104
rect 6356 7040 6372 7104
rect 6436 7040 6452 7104
rect 6516 7040 6524 7104
rect 6204 7039 6524 7040
rect 9304 7104 9624 7105
rect 9304 7040 9312 7104
rect 9376 7040 9392 7104
rect 9456 7040 9472 7104
rect 9536 7040 9552 7104
rect 9616 7040 9624 7104
rect 9304 7039 9624 7040
rect 12404 7104 12724 7105
rect 12404 7040 12412 7104
rect 12476 7040 12492 7104
rect 12556 7040 12572 7104
rect 12636 7040 12652 7104
rect 12716 7040 12724 7104
rect 12404 7039 12724 7040
rect 15504 7104 15824 7105
rect 15504 7040 15512 7104
rect 15576 7040 15592 7104
rect 15656 7040 15672 7104
rect 15736 7040 15752 7104
rect 15816 7040 15824 7104
rect 15504 7039 15824 7040
rect 18505 6762 18571 6765
rect 19200 6762 20000 6792
rect 18505 6760 20000 6762
rect 18505 6704 18510 6760
rect 18566 6704 20000 6760
rect 18505 6702 20000 6704
rect 18505 6699 18571 6702
rect 19200 6672 20000 6702
rect 4654 6560 4974 6561
rect 4654 6496 4662 6560
rect 4726 6496 4742 6560
rect 4806 6496 4822 6560
rect 4886 6496 4902 6560
rect 4966 6496 4974 6560
rect 4654 6495 4974 6496
rect 7754 6560 8074 6561
rect 7754 6496 7762 6560
rect 7826 6496 7842 6560
rect 7906 6496 7922 6560
rect 7986 6496 8002 6560
rect 8066 6496 8074 6560
rect 7754 6495 8074 6496
rect 10854 6560 11174 6561
rect 10854 6496 10862 6560
rect 10926 6496 10942 6560
rect 11006 6496 11022 6560
rect 11086 6496 11102 6560
rect 11166 6496 11174 6560
rect 10854 6495 11174 6496
rect 13954 6560 14274 6561
rect 13954 6496 13962 6560
rect 14026 6496 14042 6560
rect 14106 6496 14122 6560
rect 14186 6496 14202 6560
rect 14266 6496 14274 6560
rect 13954 6495 14274 6496
rect 17054 6560 17374 6561
rect 17054 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17222 6560
rect 17286 6496 17302 6560
rect 17366 6496 17374 6560
rect 17054 6495 17374 6496
rect 3104 6016 3424 6017
rect 3104 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3272 6016
rect 3336 5952 3352 6016
rect 3416 5952 3424 6016
rect 3104 5951 3424 5952
rect 6204 6016 6524 6017
rect 6204 5952 6212 6016
rect 6276 5952 6292 6016
rect 6356 5952 6372 6016
rect 6436 5952 6452 6016
rect 6516 5952 6524 6016
rect 6204 5951 6524 5952
rect 9304 6016 9624 6017
rect 9304 5952 9312 6016
rect 9376 5952 9392 6016
rect 9456 5952 9472 6016
rect 9536 5952 9552 6016
rect 9616 5952 9624 6016
rect 9304 5951 9624 5952
rect 12404 6016 12724 6017
rect 12404 5952 12412 6016
rect 12476 5952 12492 6016
rect 12556 5952 12572 6016
rect 12636 5952 12652 6016
rect 12716 5952 12724 6016
rect 12404 5951 12724 5952
rect 15504 6016 15824 6017
rect 15504 5952 15512 6016
rect 15576 5952 15592 6016
rect 15656 5952 15672 6016
rect 15736 5952 15752 6016
rect 15816 5952 15824 6016
rect 15504 5951 15824 5952
rect 4654 5472 4974 5473
rect 4654 5408 4662 5472
rect 4726 5408 4742 5472
rect 4806 5408 4822 5472
rect 4886 5408 4902 5472
rect 4966 5408 4974 5472
rect 4654 5407 4974 5408
rect 7754 5472 8074 5473
rect 7754 5408 7762 5472
rect 7826 5408 7842 5472
rect 7906 5408 7922 5472
rect 7986 5408 8002 5472
rect 8066 5408 8074 5472
rect 7754 5407 8074 5408
rect 10854 5472 11174 5473
rect 10854 5408 10862 5472
rect 10926 5408 10942 5472
rect 11006 5408 11022 5472
rect 11086 5408 11102 5472
rect 11166 5408 11174 5472
rect 10854 5407 11174 5408
rect 13954 5472 14274 5473
rect 13954 5408 13962 5472
rect 14026 5408 14042 5472
rect 14106 5408 14122 5472
rect 14186 5408 14202 5472
rect 14266 5408 14274 5472
rect 13954 5407 14274 5408
rect 17054 5472 17374 5473
rect 17054 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17222 5472
rect 17286 5408 17302 5472
rect 17366 5408 17374 5472
rect 17054 5407 17374 5408
rect 18505 5266 18571 5269
rect 19200 5266 20000 5296
rect 18505 5264 20000 5266
rect 18505 5208 18510 5264
rect 18566 5208 20000 5264
rect 18505 5206 20000 5208
rect 18505 5203 18571 5206
rect 19200 5176 20000 5206
rect 3104 4928 3424 4929
rect 3104 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3272 4928
rect 3336 4864 3352 4928
rect 3416 4864 3424 4928
rect 3104 4863 3424 4864
rect 6204 4928 6524 4929
rect 6204 4864 6212 4928
rect 6276 4864 6292 4928
rect 6356 4864 6372 4928
rect 6436 4864 6452 4928
rect 6516 4864 6524 4928
rect 6204 4863 6524 4864
rect 9304 4928 9624 4929
rect 9304 4864 9312 4928
rect 9376 4864 9392 4928
rect 9456 4864 9472 4928
rect 9536 4864 9552 4928
rect 9616 4864 9624 4928
rect 9304 4863 9624 4864
rect 12404 4928 12724 4929
rect 12404 4864 12412 4928
rect 12476 4864 12492 4928
rect 12556 4864 12572 4928
rect 12636 4864 12652 4928
rect 12716 4864 12724 4928
rect 12404 4863 12724 4864
rect 15504 4928 15824 4929
rect 15504 4864 15512 4928
rect 15576 4864 15592 4928
rect 15656 4864 15672 4928
rect 15736 4864 15752 4928
rect 15816 4864 15824 4928
rect 15504 4863 15824 4864
rect 4654 4384 4974 4385
rect 4654 4320 4662 4384
rect 4726 4320 4742 4384
rect 4806 4320 4822 4384
rect 4886 4320 4902 4384
rect 4966 4320 4974 4384
rect 4654 4319 4974 4320
rect 7754 4384 8074 4385
rect 7754 4320 7762 4384
rect 7826 4320 7842 4384
rect 7906 4320 7922 4384
rect 7986 4320 8002 4384
rect 8066 4320 8074 4384
rect 7754 4319 8074 4320
rect 10854 4384 11174 4385
rect 10854 4320 10862 4384
rect 10926 4320 10942 4384
rect 11006 4320 11022 4384
rect 11086 4320 11102 4384
rect 11166 4320 11174 4384
rect 10854 4319 11174 4320
rect 13954 4384 14274 4385
rect 13954 4320 13962 4384
rect 14026 4320 14042 4384
rect 14106 4320 14122 4384
rect 14186 4320 14202 4384
rect 14266 4320 14274 4384
rect 13954 4319 14274 4320
rect 17054 4384 17374 4385
rect 17054 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17222 4384
rect 17286 4320 17302 4384
rect 17366 4320 17374 4384
rect 17054 4319 17374 4320
rect 3104 3840 3424 3841
rect 3104 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3272 3840
rect 3336 3776 3352 3840
rect 3416 3776 3424 3840
rect 3104 3775 3424 3776
rect 6204 3840 6524 3841
rect 6204 3776 6212 3840
rect 6276 3776 6292 3840
rect 6356 3776 6372 3840
rect 6436 3776 6452 3840
rect 6516 3776 6524 3840
rect 6204 3775 6524 3776
rect 9304 3840 9624 3841
rect 9304 3776 9312 3840
rect 9376 3776 9392 3840
rect 9456 3776 9472 3840
rect 9536 3776 9552 3840
rect 9616 3776 9624 3840
rect 9304 3775 9624 3776
rect 12404 3840 12724 3841
rect 12404 3776 12412 3840
rect 12476 3776 12492 3840
rect 12556 3776 12572 3840
rect 12636 3776 12652 3840
rect 12716 3776 12724 3840
rect 12404 3775 12724 3776
rect 15504 3840 15824 3841
rect 15504 3776 15512 3840
rect 15576 3776 15592 3840
rect 15656 3776 15672 3840
rect 15736 3776 15752 3840
rect 15816 3776 15824 3840
rect 15504 3775 15824 3776
rect 18505 3770 18571 3773
rect 19200 3770 20000 3800
rect 18505 3768 20000 3770
rect 18505 3712 18510 3768
rect 18566 3712 20000 3768
rect 18505 3710 20000 3712
rect 18505 3707 18571 3710
rect 19200 3680 20000 3710
rect 4654 3296 4974 3297
rect 4654 3232 4662 3296
rect 4726 3232 4742 3296
rect 4806 3232 4822 3296
rect 4886 3232 4902 3296
rect 4966 3232 4974 3296
rect 4654 3231 4974 3232
rect 7754 3296 8074 3297
rect 7754 3232 7762 3296
rect 7826 3232 7842 3296
rect 7906 3232 7922 3296
rect 7986 3232 8002 3296
rect 8066 3232 8074 3296
rect 7754 3231 8074 3232
rect 10854 3296 11174 3297
rect 10854 3232 10862 3296
rect 10926 3232 10942 3296
rect 11006 3232 11022 3296
rect 11086 3232 11102 3296
rect 11166 3232 11174 3296
rect 10854 3231 11174 3232
rect 13954 3296 14274 3297
rect 13954 3232 13962 3296
rect 14026 3232 14042 3296
rect 14106 3232 14122 3296
rect 14186 3232 14202 3296
rect 14266 3232 14274 3296
rect 13954 3231 14274 3232
rect 17054 3296 17374 3297
rect 17054 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17222 3296
rect 17286 3232 17302 3296
rect 17366 3232 17374 3296
rect 17054 3231 17374 3232
rect 3104 2752 3424 2753
rect 3104 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3272 2752
rect 3336 2688 3352 2752
rect 3416 2688 3424 2752
rect 3104 2687 3424 2688
rect 6204 2752 6524 2753
rect 6204 2688 6212 2752
rect 6276 2688 6292 2752
rect 6356 2688 6372 2752
rect 6436 2688 6452 2752
rect 6516 2688 6524 2752
rect 6204 2687 6524 2688
rect 9304 2752 9624 2753
rect 9304 2688 9312 2752
rect 9376 2688 9392 2752
rect 9456 2688 9472 2752
rect 9536 2688 9552 2752
rect 9616 2688 9624 2752
rect 9304 2687 9624 2688
rect 12404 2752 12724 2753
rect 12404 2688 12412 2752
rect 12476 2688 12492 2752
rect 12556 2688 12572 2752
rect 12636 2688 12652 2752
rect 12716 2688 12724 2752
rect 12404 2687 12724 2688
rect 15504 2752 15824 2753
rect 15504 2688 15512 2752
rect 15576 2688 15592 2752
rect 15656 2688 15672 2752
rect 15736 2688 15752 2752
rect 15816 2688 15824 2752
rect 15504 2687 15824 2688
rect 17861 2274 17927 2277
rect 19200 2274 20000 2304
rect 17861 2272 20000 2274
rect 17861 2216 17866 2272
rect 17922 2216 20000 2272
rect 17861 2214 20000 2216
rect 17861 2211 17927 2214
rect 4654 2208 4974 2209
rect 4654 2144 4662 2208
rect 4726 2144 4742 2208
rect 4806 2144 4822 2208
rect 4886 2144 4902 2208
rect 4966 2144 4974 2208
rect 4654 2143 4974 2144
rect 7754 2208 8074 2209
rect 7754 2144 7762 2208
rect 7826 2144 7842 2208
rect 7906 2144 7922 2208
rect 7986 2144 8002 2208
rect 8066 2144 8074 2208
rect 7754 2143 8074 2144
rect 10854 2208 11174 2209
rect 10854 2144 10862 2208
rect 10926 2144 10942 2208
rect 11006 2144 11022 2208
rect 11086 2144 11102 2208
rect 11166 2144 11174 2208
rect 10854 2143 11174 2144
rect 13954 2208 14274 2209
rect 13954 2144 13962 2208
rect 14026 2144 14042 2208
rect 14106 2144 14122 2208
rect 14186 2144 14202 2208
rect 14266 2144 14274 2208
rect 13954 2143 14274 2144
rect 17054 2208 17374 2209
rect 17054 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17222 2208
rect 17286 2144 17302 2208
rect 17366 2144 17374 2208
rect 19200 2184 20000 2214
rect 17054 2143 17374 2144
rect 8017 2002 8083 2005
rect 9397 2002 9463 2005
rect 8017 2000 9463 2002
rect 8017 1944 8022 2000
rect 8078 1944 9402 2000
rect 9458 1944 9463 2000
rect 8017 1942 9463 1944
rect 8017 1939 8083 1942
rect 9397 1939 9463 1942
rect 10133 2002 10199 2005
rect 11145 2002 11211 2005
rect 10133 2000 11211 2002
rect 10133 1944 10138 2000
rect 10194 1944 11150 2000
rect 11206 1944 11211 2000
rect 10133 1942 11211 1944
rect 10133 1939 10199 1942
rect 11145 1939 11211 1942
rect 11237 1866 11303 1869
rect 14733 1866 14799 1869
rect 11237 1864 14799 1866
rect 11237 1808 11242 1864
rect 11298 1808 14738 1864
rect 14794 1808 14799 1864
rect 11237 1806 14799 1808
rect 11237 1803 11303 1806
rect 14733 1803 14799 1806
rect 3104 1664 3424 1665
rect 3104 1600 3112 1664
rect 3176 1600 3192 1664
rect 3256 1600 3272 1664
rect 3336 1600 3352 1664
rect 3416 1600 3424 1664
rect 3104 1599 3424 1600
rect 6204 1664 6524 1665
rect 6204 1600 6212 1664
rect 6276 1600 6292 1664
rect 6356 1600 6372 1664
rect 6436 1600 6452 1664
rect 6516 1600 6524 1664
rect 6204 1599 6524 1600
rect 9304 1664 9624 1665
rect 9304 1600 9312 1664
rect 9376 1600 9392 1664
rect 9456 1600 9472 1664
rect 9536 1600 9552 1664
rect 9616 1600 9624 1664
rect 9304 1599 9624 1600
rect 12404 1664 12724 1665
rect 12404 1600 12412 1664
rect 12476 1600 12492 1664
rect 12556 1600 12572 1664
rect 12636 1600 12652 1664
rect 12716 1600 12724 1664
rect 12404 1599 12724 1600
rect 15504 1664 15824 1665
rect 15504 1600 15512 1664
rect 15576 1600 15592 1664
rect 15656 1600 15672 1664
rect 15736 1600 15752 1664
rect 15816 1600 15824 1664
rect 15504 1599 15824 1600
rect 7189 1594 7255 1597
rect 7189 1592 7298 1594
rect 7189 1536 7194 1592
rect 7250 1536 7298 1592
rect 7189 1531 7298 1536
rect 7238 1458 7298 1531
rect 12617 1458 12683 1461
rect 14549 1458 14615 1461
rect 7238 1456 14615 1458
rect 7238 1400 12622 1456
rect 12678 1400 14554 1456
rect 14610 1400 14615 1456
rect 7238 1398 14615 1400
rect 12617 1395 12683 1398
rect 14549 1395 14615 1398
rect 12065 1322 12131 1325
rect 13537 1322 13603 1325
rect 12065 1320 13603 1322
rect 12065 1264 12070 1320
rect 12126 1264 13542 1320
rect 13598 1264 13603 1320
rect 12065 1262 13603 1264
rect 12065 1259 12131 1262
rect 13537 1259 13603 1262
rect 4654 1120 4974 1121
rect 4654 1056 4662 1120
rect 4726 1056 4742 1120
rect 4806 1056 4822 1120
rect 4886 1056 4902 1120
rect 4966 1056 4974 1120
rect 4654 1055 4974 1056
rect 7754 1120 8074 1121
rect 7754 1056 7762 1120
rect 7826 1056 7842 1120
rect 7906 1056 7922 1120
rect 7986 1056 8002 1120
rect 8066 1056 8074 1120
rect 7754 1055 8074 1056
rect 10854 1120 11174 1121
rect 10854 1056 10862 1120
rect 10926 1056 10942 1120
rect 11006 1056 11022 1120
rect 11086 1056 11102 1120
rect 11166 1056 11174 1120
rect 10854 1055 11174 1056
rect 13954 1120 14274 1121
rect 13954 1056 13962 1120
rect 14026 1056 14042 1120
rect 14106 1056 14122 1120
rect 14186 1056 14202 1120
rect 14266 1056 14274 1120
rect 13954 1055 14274 1056
rect 17054 1120 17374 1121
rect 17054 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17222 1120
rect 17286 1056 17302 1120
rect 17366 1056 17374 1120
rect 17054 1055 17374 1056
rect 18505 778 18571 781
rect 19200 778 20000 808
rect 18505 776 20000 778
rect 18505 720 18510 776
rect 18566 720 20000 776
rect 18505 718 20000 720
rect 18505 715 18571 718
rect 19200 688 20000 718
rect 3104 576 3424 577
rect 3104 512 3112 576
rect 3176 512 3192 576
rect 3256 512 3272 576
rect 3336 512 3352 576
rect 3416 512 3424 576
rect 3104 511 3424 512
rect 6204 576 6524 577
rect 6204 512 6212 576
rect 6276 512 6292 576
rect 6356 512 6372 576
rect 6436 512 6452 576
rect 6516 512 6524 576
rect 6204 511 6524 512
rect 9304 576 9624 577
rect 9304 512 9312 576
rect 9376 512 9392 576
rect 9456 512 9472 576
rect 9536 512 9552 576
rect 9616 512 9624 576
rect 9304 511 9624 512
rect 12404 576 12724 577
rect 12404 512 12412 576
rect 12476 512 12492 576
rect 12556 512 12572 576
rect 12636 512 12652 576
rect 12716 512 12724 576
rect 12404 511 12724 512
rect 15504 576 15824 577
rect 15504 512 15512 576
rect 15576 512 15592 576
rect 15656 512 15672 576
rect 15736 512 15752 576
rect 15816 512 15824 576
rect 15504 511 15824 512
rect 4654 32 4974 33
rect 4654 -32 4662 32
rect 4726 -32 4742 32
rect 4806 -32 4822 32
rect 4886 -32 4902 32
rect 4966 -32 4974 32
rect 4654 -33 4974 -32
rect 7754 32 8074 33
rect 7754 -32 7762 32
rect 7826 -32 7842 32
rect 7906 -32 7922 32
rect 7986 -32 8002 32
rect 8066 -32 8074 32
rect 7754 -33 8074 -32
rect 10854 32 11174 33
rect 10854 -32 10862 32
rect 10926 -32 10942 32
rect 11006 -32 11022 32
rect 11086 -32 11102 32
rect 11166 -32 11174 32
rect 10854 -33 11174 -32
rect 13954 32 14274 33
rect 13954 -32 13962 32
rect 14026 -32 14042 32
rect 14106 -32 14122 32
rect 14186 -32 14202 32
rect 14266 -32 14274 32
rect 13954 -33 14274 -32
rect 17054 32 17374 33
rect 17054 -32 17062 32
rect 17126 -32 17142 32
rect 17206 -32 17222 32
rect 17286 -32 17302 32
rect 17366 -32 17374 32
rect 17054 -33 17374 -32
<< via3 >>
rect 4662 10908 4726 10912
rect 4662 10852 4666 10908
rect 4666 10852 4722 10908
rect 4722 10852 4726 10908
rect 4662 10848 4726 10852
rect 4742 10908 4806 10912
rect 4742 10852 4746 10908
rect 4746 10852 4802 10908
rect 4802 10852 4806 10908
rect 4742 10848 4806 10852
rect 4822 10908 4886 10912
rect 4822 10852 4826 10908
rect 4826 10852 4882 10908
rect 4882 10852 4886 10908
rect 4822 10848 4886 10852
rect 4902 10908 4966 10912
rect 4902 10852 4906 10908
rect 4906 10852 4962 10908
rect 4962 10852 4966 10908
rect 4902 10848 4966 10852
rect 7762 10908 7826 10912
rect 7762 10852 7766 10908
rect 7766 10852 7822 10908
rect 7822 10852 7826 10908
rect 7762 10848 7826 10852
rect 7842 10908 7906 10912
rect 7842 10852 7846 10908
rect 7846 10852 7902 10908
rect 7902 10852 7906 10908
rect 7842 10848 7906 10852
rect 7922 10908 7986 10912
rect 7922 10852 7926 10908
rect 7926 10852 7982 10908
rect 7982 10852 7986 10908
rect 7922 10848 7986 10852
rect 8002 10908 8066 10912
rect 8002 10852 8006 10908
rect 8006 10852 8062 10908
rect 8062 10852 8066 10908
rect 8002 10848 8066 10852
rect 10862 10908 10926 10912
rect 10862 10852 10866 10908
rect 10866 10852 10922 10908
rect 10922 10852 10926 10908
rect 10862 10848 10926 10852
rect 10942 10908 11006 10912
rect 10942 10852 10946 10908
rect 10946 10852 11002 10908
rect 11002 10852 11006 10908
rect 10942 10848 11006 10852
rect 11022 10908 11086 10912
rect 11022 10852 11026 10908
rect 11026 10852 11082 10908
rect 11082 10852 11086 10908
rect 11022 10848 11086 10852
rect 11102 10908 11166 10912
rect 11102 10852 11106 10908
rect 11106 10852 11162 10908
rect 11162 10852 11166 10908
rect 11102 10848 11166 10852
rect 13962 10908 14026 10912
rect 13962 10852 13966 10908
rect 13966 10852 14022 10908
rect 14022 10852 14026 10908
rect 13962 10848 14026 10852
rect 14042 10908 14106 10912
rect 14042 10852 14046 10908
rect 14046 10852 14102 10908
rect 14102 10852 14106 10908
rect 14042 10848 14106 10852
rect 14122 10908 14186 10912
rect 14122 10852 14126 10908
rect 14126 10852 14182 10908
rect 14182 10852 14186 10908
rect 14122 10848 14186 10852
rect 14202 10908 14266 10912
rect 14202 10852 14206 10908
rect 14206 10852 14262 10908
rect 14262 10852 14266 10908
rect 14202 10848 14266 10852
rect 17062 10908 17126 10912
rect 17062 10852 17066 10908
rect 17066 10852 17122 10908
rect 17122 10852 17126 10908
rect 17062 10848 17126 10852
rect 17142 10908 17206 10912
rect 17142 10852 17146 10908
rect 17146 10852 17202 10908
rect 17202 10852 17206 10908
rect 17142 10848 17206 10852
rect 17222 10908 17286 10912
rect 17222 10852 17226 10908
rect 17226 10852 17282 10908
rect 17282 10852 17286 10908
rect 17222 10848 17286 10852
rect 17302 10908 17366 10912
rect 17302 10852 17306 10908
rect 17306 10852 17362 10908
rect 17362 10852 17366 10908
rect 17302 10848 17366 10852
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 3272 10364 3336 10368
rect 3272 10308 3276 10364
rect 3276 10308 3332 10364
rect 3332 10308 3336 10364
rect 3272 10304 3336 10308
rect 3352 10364 3416 10368
rect 3352 10308 3356 10364
rect 3356 10308 3412 10364
rect 3412 10308 3416 10364
rect 3352 10304 3416 10308
rect 6212 10364 6276 10368
rect 6212 10308 6216 10364
rect 6216 10308 6272 10364
rect 6272 10308 6276 10364
rect 6212 10304 6276 10308
rect 6292 10364 6356 10368
rect 6292 10308 6296 10364
rect 6296 10308 6352 10364
rect 6352 10308 6356 10364
rect 6292 10304 6356 10308
rect 6372 10364 6436 10368
rect 6372 10308 6376 10364
rect 6376 10308 6432 10364
rect 6432 10308 6436 10364
rect 6372 10304 6436 10308
rect 6452 10364 6516 10368
rect 6452 10308 6456 10364
rect 6456 10308 6512 10364
rect 6512 10308 6516 10364
rect 6452 10304 6516 10308
rect 9312 10364 9376 10368
rect 9312 10308 9316 10364
rect 9316 10308 9372 10364
rect 9372 10308 9376 10364
rect 9312 10304 9376 10308
rect 9392 10364 9456 10368
rect 9392 10308 9396 10364
rect 9396 10308 9452 10364
rect 9452 10308 9456 10364
rect 9392 10304 9456 10308
rect 9472 10364 9536 10368
rect 9472 10308 9476 10364
rect 9476 10308 9532 10364
rect 9532 10308 9536 10364
rect 9472 10304 9536 10308
rect 9552 10364 9616 10368
rect 9552 10308 9556 10364
rect 9556 10308 9612 10364
rect 9612 10308 9616 10364
rect 9552 10304 9616 10308
rect 12412 10364 12476 10368
rect 12412 10308 12416 10364
rect 12416 10308 12472 10364
rect 12472 10308 12476 10364
rect 12412 10304 12476 10308
rect 12492 10364 12556 10368
rect 12492 10308 12496 10364
rect 12496 10308 12552 10364
rect 12552 10308 12556 10364
rect 12492 10304 12556 10308
rect 12572 10364 12636 10368
rect 12572 10308 12576 10364
rect 12576 10308 12632 10364
rect 12632 10308 12636 10364
rect 12572 10304 12636 10308
rect 12652 10364 12716 10368
rect 12652 10308 12656 10364
rect 12656 10308 12712 10364
rect 12712 10308 12716 10364
rect 12652 10304 12716 10308
rect 15512 10364 15576 10368
rect 15512 10308 15516 10364
rect 15516 10308 15572 10364
rect 15572 10308 15576 10364
rect 15512 10304 15576 10308
rect 15592 10364 15656 10368
rect 15592 10308 15596 10364
rect 15596 10308 15652 10364
rect 15652 10308 15656 10364
rect 15592 10304 15656 10308
rect 15672 10364 15736 10368
rect 15672 10308 15676 10364
rect 15676 10308 15732 10364
rect 15732 10308 15736 10364
rect 15672 10304 15736 10308
rect 15752 10364 15816 10368
rect 15752 10308 15756 10364
rect 15756 10308 15812 10364
rect 15812 10308 15816 10364
rect 15752 10304 15816 10308
rect 4662 9820 4726 9824
rect 4662 9764 4666 9820
rect 4666 9764 4722 9820
rect 4722 9764 4726 9820
rect 4662 9760 4726 9764
rect 4742 9820 4806 9824
rect 4742 9764 4746 9820
rect 4746 9764 4802 9820
rect 4802 9764 4806 9820
rect 4742 9760 4806 9764
rect 4822 9820 4886 9824
rect 4822 9764 4826 9820
rect 4826 9764 4882 9820
rect 4882 9764 4886 9820
rect 4822 9760 4886 9764
rect 4902 9820 4966 9824
rect 4902 9764 4906 9820
rect 4906 9764 4962 9820
rect 4962 9764 4966 9820
rect 4902 9760 4966 9764
rect 7762 9820 7826 9824
rect 7762 9764 7766 9820
rect 7766 9764 7822 9820
rect 7822 9764 7826 9820
rect 7762 9760 7826 9764
rect 7842 9820 7906 9824
rect 7842 9764 7846 9820
rect 7846 9764 7902 9820
rect 7902 9764 7906 9820
rect 7842 9760 7906 9764
rect 7922 9820 7986 9824
rect 7922 9764 7926 9820
rect 7926 9764 7982 9820
rect 7982 9764 7986 9820
rect 7922 9760 7986 9764
rect 8002 9820 8066 9824
rect 8002 9764 8006 9820
rect 8006 9764 8062 9820
rect 8062 9764 8066 9820
rect 8002 9760 8066 9764
rect 10862 9820 10926 9824
rect 10862 9764 10866 9820
rect 10866 9764 10922 9820
rect 10922 9764 10926 9820
rect 10862 9760 10926 9764
rect 10942 9820 11006 9824
rect 10942 9764 10946 9820
rect 10946 9764 11002 9820
rect 11002 9764 11006 9820
rect 10942 9760 11006 9764
rect 11022 9820 11086 9824
rect 11022 9764 11026 9820
rect 11026 9764 11082 9820
rect 11082 9764 11086 9820
rect 11022 9760 11086 9764
rect 11102 9820 11166 9824
rect 11102 9764 11106 9820
rect 11106 9764 11162 9820
rect 11162 9764 11166 9820
rect 11102 9760 11166 9764
rect 13962 9820 14026 9824
rect 13962 9764 13966 9820
rect 13966 9764 14022 9820
rect 14022 9764 14026 9820
rect 13962 9760 14026 9764
rect 14042 9820 14106 9824
rect 14042 9764 14046 9820
rect 14046 9764 14102 9820
rect 14102 9764 14106 9820
rect 14042 9760 14106 9764
rect 14122 9820 14186 9824
rect 14122 9764 14126 9820
rect 14126 9764 14182 9820
rect 14182 9764 14186 9820
rect 14122 9760 14186 9764
rect 14202 9820 14266 9824
rect 14202 9764 14206 9820
rect 14206 9764 14262 9820
rect 14262 9764 14266 9820
rect 14202 9760 14266 9764
rect 17062 9820 17126 9824
rect 17062 9764 17066 9820
rect 17066 9764 17122 9820
rect 17122 9764 17126 9820
rect 17062 9760 17126 9764
rect 17142 9820 17206 9824
rect 17142 9764 17146 9820
rect 17146 9764 17202 9820
rect 17202 9764 17206 9820
rect 17142 9760 17206 9764
rect 17222 9820 17286 9824
rect 17222 9764 17226 9820
rect 17226 9764 17282 9820
rect 17282 9764 17286 9820
rect 17222 9760 17286 9764
rect 17302 9820 17366 9824
rect 17302 9764 17306 9820
rect 17306 9764 17362 9820
rect 17362 9764 17366 9820
rect 17302 9760 17366 9764
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 3272 9276 3336 9280
rect 3272 9220 3276 9276
rect 3276 9220 3332 9276
rect 3332 9220 3336 9276
rect 3272 9216 3336 9220
rect 3352 9276 3416 9280
rect 3352 9220 3356 9276
rect 3356 9220 3412 9276
rect 3412 9220 3416 9276
rect 3352 9216 3416 9220
rect 6212 9276 6276 9280
rect 6212 9220 6216 9276
rect 6216 9220 6272 9276
rect 6272 9220 6276 9276
rect 6212 9216 6276 9220
rect 6292 9276 6356 9280
rect 6292 9220 6296 9276
rect 6296 9220 6352 9276
rect 6352 9220 6356 9276
rect 6292 9216 6356 9220
rect 6372 9276 6436 9280
rect 6372 9220 6376 9276
rect 6376 9220 6432 9276
rect 6432 9220 6436 9276
rect 6372 9216 6436 9220
rect 6452 9276 6516 9280
rect 6452 9220 6456 9276
rect 6456 9220 6512 9276
rect 6512 9220 6516 9276
rect 6452 9216 6516 9220
rect 9312 9276 9376 9280
rect 9312 9220 9316 9276
rect 9316 9220 9372 9276
rect 9372 9220 9376 9276
rect 9312 9216 9376 9220
rect 9392 9276 9456 9280
rect 9392 9220 9396 9276
rect 9396 9220 9452 9276
rect 9452 9220 9456 9276
rect 9392 9216 9456 9220
rect 9472 9276 9536 9280
rect 9472 9220 9476 9276
rect 9476 9220 9532 9276
rect 9532 9220 9536 9276
rect 9472 9216 9536 9220
rect 9552 9276 9616 9280
rect 9552 9220 9556 9276
rect 9556 9220 9612 9276
rect 9612 9220 9616 9276
rect 9552 9216 9616 9220
rect 12412 9276 12476 9280
rect 12412 9220 12416 9276
rect 12416 9220 12472 9276
rect 12472 9220 12476 9276
rect 12412 9216 12476 9220
rect 12492 9276 12556 9280
rect 12492 9220 12496 9276
rect 12496 9220 12552 9276
rect 12552 9220 12556 9276
rect 12492 9216 12556 9220
rect 12572 9276 12636 9280
rect 12572 9220 12576 9276
rect 12576 9220 12632 9276
rect 12632 9220 12636 9276
rect 12572 9216 12636 9220
rect 12652 9276 12716 9280
rect 12652 9220 12656 9276
rect 12656 9220 12712 9276
rect 12712 9220 12716 9276
rect 12652 9216 12716 9220
rect 15512 9276 15576 9280
rect 15512 9220 15516 9276
rect 15516 9220 15572 9276
rect 15572 9220 15576 9276
rect 15512 9216 15576 9220
rect 15592 9276 15656 9280
rect 15592 9220 15596 9276
rect 15596 9220 15652 9276
rect 15652 9220 15656 9276
rect 15592 9216 15656 9220
rect 15672 9276 15736 9280
rect 15672 9220 15676 9276
rect 15676 9220 15732 9276
rect 15732 9220 15736 9276
rect 15672 9216 15736 9220
rect 15752 9276 15816 9280
rect 15752 9220 15756 9276
rect 15756 9220 15812 9276
rect 15812 9220 15816 9276
rect 15752 9216 15816 9220
rect 4662 8732 4726 8736
rect 4662 8676 4666 8732
rect 4666 8676 4722 8732
rect 4722 8676 4726 8732
rect 4662 8672 4726 8676
rect 4742 8732 4806 8736
rect 4742 8676 4746 8732
rect 4746 8676 4802 8732
rect 4802 8676 4806 8732
rect 4742 8672 4806 8676
rect 4822 8732 4886 8736
rect 4822 8676 4826 8732
rect 4826 8676 4882 8732
rect 4882 8676 4886 8732
rect 4822 8672 4886 8676
rect 4902 8732 4966 8736
rect 4902 8676 4906 8732
rect 4906 8676 4962 8732
rect 4962 8676 4966 8732
rect 4902 8672 4966 8676
rect 7762 8732 7826 8736
rect 7762 8676 7766 8732
rect 7766 8676 7822 8732
rect 7822 8676 7826 8732
rect 7762 8672 7826 8676
rect 7842 8732 7906 8736
rect 7842 8676 7846 8732
rect 7846 8676 7902 8732
rect 7902 8676 7906 8732
rect 7842 8672 7906 8676
rect 7922 8732 7986 8736
rect 7922 8676 7926 8732
rect 7926 8676 7982 8732
rect 7982 8676 7986 8732
rect 7922 8672 7986 8676
rect 8002 8732 8066 8736
rect 8002 8676 8006 8732
rect 8006 8676 8062 8732
rect 8062 8676 8066 8732
rect 8002 8672 8066 8676
rect 10862 8732 10926 8736
rect 10862 8676 10866 8732
rect 10866 8676 10922 8732
rect 10922 8676 10926 8732
rect 10862 8672 10926 8676
rect 10942 8732 11006 8736
rect 10942 8676 10946 8732
rect 10946 8676 11002 8732
rect 11002 8676 11006 8732
rect 10942 8672 11006 8676
rect 11022 8732 11086 8736
rect 11022 8676 11026 8732
rect 11026 8676 11082 8732
rect 11082 8676 11086 8732
rect 11022 8672 11086 8676
rect 11102 8732 11166 8736
rect 11102 8676 11106 8732
rect 11106 8676 11162 8732
rect 11162 8676 11166 8732
rect 11102 8672 11166 8676
rect 13962 8732 14026 8736
rect 13962 8676 13966 8732
rect 13966 8676 14022 8732
rect 14022 8676 14026 8732
rect 13962 8672 14026 8676
rect 14042 8732 14106 8736
rect 14042 8676 14046 8732
rect 14046 8676 14102 8732
rect 14102 8676 14106 8732
rect 14042 8672 14106 8676
rect 14122 8732 14186 8736
rect 14122 8676 14126 8732
rect 14126 8676 14182 8732
rect 14182 8676 14186 8732
rect 14122 8672 14186 8676
rect 14202 8732 14266 8736
rect 14202 8676 14206 8732
rect 14206 8676 14262 8732
rect 14262 8676 14266 8732
rect 14202 8672 14266 8676
rect 17062 8732 17126 8736
rect 17062 8676 17066 8732
rect 17066 8676 17122 8732
rect 17122 8676 17126 8732
rect 17062 8672 17126 8676
rect 17142 8732 17206 8736
rect 17142 8676 17146 8732
rect 17146 8676 17202 8732
rect 17202 8676 17206 8732
rect 17142 8672 17206 8676
rect 17222 8732 17286 8736
rect 17222 8676 17226 8732
rect 17226 8676 17282 8732
rect 17282 8676 17286 8732
rect 17222 8672 17286 8676
rect 17302 8732 17366 8736
rect 17302 8676 17306 8732
rect 17306 8676 17362 8732
rect 17362 8676 17366 8732
rect 17302 8672 17366 8676
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 3272 8188 3336 8192
rect 3272 8132 3276 8188
rect 3276 8132 3332 8188
rect 3332 8132 3336 8188
rect 3272 8128 3336 8132
rect 3352 8188 3416 8192
rect 3352 8132 3356 8188
rect 3356 8132 3412 8188
rect 3412 8132 3416 8188
rect 3352 8128 3416 8132
rect 6212 8188 6276 8192
rect 6212 8132 6216 8188
rect 6216 8132 6272 8188
rect 6272 8132 6276 8188
rect 6212 8128 6276 8132
rect 6292 8188 6356 8192
rect 6292 8132 6296 8188
rect 6296 8132 6352 8188
rect 6352 8132 6356 8188
rect 6292 8128 6356 8132
rect 6372 8188 6436 8192
rect 6372 8132 6376 8188
rect 6376 8132 6432 8188
rect 6432 8132 6436 8188
rect 6372 8128 6436 8132
rect 6452 8188 6516 8192
rect 6452 8132 6456 8188
rect 6456 8132 6512 8188
rect 6512 8132 6516 8188
rect 6452 8128 6516 8132
rect 9312 8188 9376 8192
rect 9312 8132 9316 8188
rect 9316 8132 9372 8188
rect 9372 8132 9376 8188
rect 9312 8128 9376 8132
rect 9392 8188 9456 8192
rect 9392 8132 9396 8188
rect 9396 8132 9452 8188
rect 9452 8132 9456 8188
rect 9392 8128 9456 8132
rect 9472 8188 9536 8192
rect 9472 8132 9476 8188
rect 9476 8132 9532 8188
rect 9532 8132 9536 8188
rect 9472 8128 9536 8132
rect 9552 8188 9616 8192
rect 9552 8132 9556 8188
rect 9556 8132 9612 8188
rect 9612 8132 9616 8188
rect 9552 8128 9616 8132
rect 12412 8188 12476 8192
rect 12412 8132 12416 8188
rect 12416 8132 12472 8188
rect 12472 8132 12476 8188
rect 12412 8128 12476 8132
rect 12492 8188 12556 8192
rect 12492 8132 12496 8188
rect 12496 8132 12552 8188
rect 12552 8132 12556 8188
rect 12492 8128 12556 8132
rect 12572 8188 12636 8192
rect 12572 8132 12576 8188
rect 12576 8132 12632 8188
rect 12632 8132 12636 8188
rect 12572 8128 12636 8132
rect 12652 8188 12716 8192
rect 12652 8132 12656 8188
rect 12656 8132 12712 8188
rect 12712 8132 12716 8188
rect 12652 8128 12716 8132
rect 15512 8188 15576 8192
rect 15512 8132 15516 8188
rect 15516 8132 15572 8188
rect 15572 8132 15576 8188
rect 15512 8128 15576 8132
rect 15592 8188 15656 8192
rect 15592 8132 15596 8188
rect 15596 8132 15652 8188
rect 15652 8132 15656 8188
rect 15592 8128 15656 8132
rect 15672 8188 15736 8192
rect 15672 8132 15676 8188
rect 15676 8132 15732 8188
rect 15732 8132 15736 8188
rect 15672 8128 15736 8132
rect 15752 8188 15816 8192
rect 15752 8132 15756 8188
rect 15756 8132 15812 8188
rect 15812 8132 15816 8188
rect 15752 8128 15816 8132
rect 4662 7644 4726 7648
rect 4662 7588 4666 7644
rect 4666 7588 4722 7644
rect 4722 7588 4726 7644
rect 4662 7584 4726 7588
rect 4742 7644 4806 7648
rect 4742 7588 4746 7644
rect 4746 7588 4802 7644
rect 4802 7588 4806 7644
rect 4742 7584 4806 7588
rect 4822 7644 4886 7648
rect 4822 7588 4826 7644
rect 4826 7588 4882 7644
rect 4882 7588 4886 7644
rect 4822 7584 4886 7588
rect 4902 7644 4966 7648
rect 4902 7588 4906 7644
rect 4906 7588 4962 7644
rect 4962 7588 4966 7644
rect 4902 7584 4966 7588
rect 7762 7644 7826 7648
rect 7762 7588 7766 7644
rect 7766 7588 7822 7644
rect 7822 7588 7826 7644
rect 7762 7584 7826 7588
rect 7842 7644 7906 7648
rect 7842 7588 7846 7644
rect 7846 7588 7902 7644
rect 7902 7588 7906 7644
rect 7842 7584 7906 7588
rect 7922 7644 7986 7648
rect 7922 7588 7926 7644
rect 7926 7588 7982 7644
rect 7982 7588 7986 7644
rect 7922 7584 7986 7588
rect 8002 7644 8066 7648
rect 8002 7588 8006 7644
rect 8006 7588 8062 7644
rect 8062 7588 8066 7644
rect 8002 7584 8066 7588
rect 10862 7644 10926 7648
rect 10862 7588 10866 7644
rect 10866 7588 10922 7644
rect 10922 7588 10926 7644
rect 10862 7584 10926 7588
rect 10942 7644 11006 7648
rect 10942 7588 10946 7644
rect 10946 7588 11002 7644
rect 11002 7588 11006 7644
rect 10942 7584 11006 7588
rect 11022 7644 11086 7648
rect 11022 7588 11026 7644
rect 11026 7588 11082 7644
rect 11082 7588 11086 7644
rect 11022 7584 11086 7588
rect 11102 7644 11166 7648
rect 11102 7588 11106 7644
rect 11106 7588 11162 7644
rect 11162 7588 11166 7644
rect 11102 7584 11166 7588
rect 13962 7644 14026 7648
rect 13962 7588 13966 7644
rect 13966 7588 14022 7644
rect 14022 7588 14026 7644
rect 13962 7584 14026 7588
rect 14042 7644 14106 7648
rect 14042 7588 14046 7644
rect 14046 7588 14102 7644
rect 14102 7588 14106 7644
rect 14042 7584 14106 7588
rect 14122 7644 14186 7648
rect 14122 7588 14126 7644
rect 14126 7588 14182 7644
rect 14182 7588 14186 7644
rect 14122 7584 14186 7588
rect 14202 7644 14266 7648
rect 14202 7588 14206 7644
rect 14206 7588 14262 7644
rect 14262 7588 14266 7644
rect 14202 7584 14266 7588
rect 17062 7644 17126 7648
rect 17062 7588 17066 7644
rect 17066 7588 17122 7644
rect 17122 7588 17126 7644
rect 17062 7584 17126 7588
rect 17142 7644 17206 7648
rect 17142 7588 17146 7644
rect 17146 7588 17202 7644
rect 17202 7588 17206 7644
rect 17142 7584 17206 7588
rect 17222 7644 17286 7648
rect 17222 7588 17226 7644
rect 17226 7588 17282 7644
rect 17282 7588 17286 7644
rect 17222 7584 17286 7588
rect 17302 7644 17366 7648
rect 17302 7588 17306 7644
rect 17306 7588 17362 7644
rect 17362 7588 17366 7644
rect 17302 7584 17366 7588
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 3272 7100 3336 7104
rect 3272 7044 3276 7100
rect 3276 7044 3332 7100
rect 3332 7044 3336 7100
rect 3272 7040 3336 7044
rect 3352 7100 3416 7104
rect 3352 7044 3356 7100
rect 3356 7044 3412 7100
rect 3412 7044 3416 7100
rect 3352 7040 3416 7044
rect 6212 7100 6276 7104
rect 6212 7044 6216 7100
rect 6216 7044 6272 7100
rect 6272 7044 6276 7100
rect 6212 7040 6276 7044
rect 6292 7100 6356 7104
rect 6292 7044 6296 7100
rect 6296 7044 6352 7100
rect 6352 7044 6356 7100
rect 6292 7040 6356 7044
rect 6372 7100 6436 7104
rect 6372 7044 6376 7100
rect 6376 7044 6432 7100
rect 6432 7044 6436 7100
rect 6372 7040 6436 7044
rect 6452 7100 6516 7104
rect 6452 7044 6456 7100
rect 6456 7044 6512 7100
rect 6512 7044 6516 7100
rect 6452 7040 6516 7044
rect 9312 7100 9376 7104
rect 9312 7044 9316 7100
rect 9316 7044 9372 7100
rect 9372 7044 9376 7100
rect 9312 7040 9376 7044
rect 9392 7100 9456 7104
rect 9392 7044 9396 7100
rect 9396 7044 9452 7100
rect 9452 7044 9456 7100
rect 9392 7040 9456 7044
rect 9472 7100 9536 7104
rect 9472 7044 9476 7100
rect 9476 7044 9532 7100
rect 9532 7044 9536 7100
rect 9472 7040 9536 7044
rect 9552 7100 9616 7104
rect 9552 7044 9556 7100
rect 9556 7044 9612 7100
rect 9612 7044 9616 7100
rect 9552 7040 9616 7044
rect 12412 7100 12476 7104
rect 12412 7044 12416 7100
rect 12416 7044 12472 7100
rect 12472 7044 12476 7100
rect 12412 7040 12476 7044
rect 12492 7100 12556 7104
rect 12492 7044 12496 7100
rect 12496 7044 12552 7100
rect 12552 7044 12556 7100
rect 12492 7040 12556 7044
rect 12572 7100 12636 7104
rect 12572 7044 12576 7100
rect 12576 7044 12632 7100
rect 12632 7044 12636 7100
rect 12572 7040 12636 7044
rect 12652 7100 12716 7104
rect 12652 7044 12656 7100
rect 12656 7044 12712 7100
rect 12712 7044 12716 7100
rect 12652 7040 12716 7044
rect 15512 7100 15576 7104
rect 15512 7044 15516 7100
rect 15516 7044 15572 7100
rect 15572 7044 15576 7100
rect 15512 7040 15576 7044
rect 15592 7100 15656 7104
rect 15592 7044 15596 7100
rect 15596 7044 15652 7100
rect 15652 7044 15656 7100
rect 15592 7040 15656 7044
rect 15672 7100 15736 7104
rect 15672 7044 15676 7100
rect 15676 7044 15732 7100
rect 15732 7044 15736 7100
rect 15672 7040 15736 7044
rect 15752 7100 15816 7104
rect 15752 7044 15756 7100
rect 15756 7044 15812 7100
rect 15812 7044 15816 7100
rect 15752 7040 15816 7044
rect 4662 6556 4726 6560
rect 4662 6500 4666 6556
rect 4666 6500 4722 6556
rect 4722 6500 4726 6556
rect 4662 6496 4726 6500
rect 4742 6556 4806 6560
rect 4742 6500 4746 6556
rect 4746 6500 4802 6556
rect 4802 6500 4806 6556
rect 4742 6496 4806 6500
rect 4822 6556 4886 6560
rect 4822 6500 4826 6556
rect 4826 6500 4882 6556
rect 4882 6500 4886 6556
rect 4822 6496 4886 6500
rect 4902 6556 4966 6560
rect 4902 6500 4906 6556
rect 4906 6500 4962 6556
rect 4962 6500 4966 6556
rect 4902 6496 4966 6500
rect 7762 6556 7826 6560
rect 7762 6500 7766 6556
rect 7766 6500 7822 6556
rect 7822 6500 7826 6556
rect 7762 6496 7826 6500
rect 7842 6556 7906 6560
rect 7842 6500 7846 6556
rect 7846 6500 7902 6556
rect 7902 6500 7906 6556
rect 7842 6496 7906 6500
rect 7922 6556 7986 6560
rect 7922 6500 7926 6556
rect 7926 6500 7982 6556
rect 7982 6500 7986 6556
rect 7922 6496 7986 6500
rect 8002 6556 8066 6560
rect 8002 6500 8006 6556
rect 8006 6500 8062 6556
rect 8062 6500 8066 6556
rect 8002 6496 8066 6500
rect 10862 6556 10926 6560
rect 10862 6500 10866 6556
rect 10866 6500 10922 6556
rect 10922 6500 10926 6556
rect 10862 6496 10926 6500
rect 10942 6556 11006 6560
rect 10942 6500 10946 6556
rect 10946 6500 11002 6556
rect 11002 6500 11006 6556
rect 10942 6496 11006 6500
rect 11022 6556 11086 6560
rect 11022 6500 11026 6556
rect 11026 6500 11082 6556
rect 11082 6500 11086 6556
rect 11022 6496 11086 6500
rect 11102 6556 11166 6560
rect 11102 6500 11106 6556
rect 11106 6500 11162 6556
rect 11162 6500 11166 6556
rect 11102 6496 11166 6500
rect 13962 6556 14026 6560
rect 13962 6500 13966 6556
rect 13966 6500 14022 6556
rect 14022 6500 14026 6556
rect 13962 6496 14026 6500
rect 14042 6556 14106 6560
rect 14042 6500 14046 6556
rect 14046 6500 14102 6556
rect 14102 6500 14106 6556
rect 14042 6496 14106 6500
rect 14122 6556 14186 6560
rect 14122 6500 14126 6556
rect 14126 6500 14182 6556
rect 14182 6500 14186 6556
rect 14122 6496 14186 6500
rect 14202 6556 14266 6560
rect 14202 6500 14206 6556
rect 14206 6500 14262 6556
rect 14262 6500 14266 6556
rect 14202 6496 14266 6500
rect 17062 6556 17126 6560
rect 17062 6500 17066 6556
rect 17066 6500 17122 6556
rect 17122 6500 17126 6556
rect 17062 6496 17126 6500
rect 17142 6556 17206 6560
rect 17142 6500 17146 6556
rect 17146 6500 17202 6556
rect 17202 6500 17206 6556
rect 17142 6496 17206 6500
rect 17222 6556 17286 6560
rect 17222 6500 17226 6556
rect 17226 6500 17282 6556
rect 17282 6500 17286 6556
rect 17222 6496 17286 6500
rect 17302 6556 17366 6560
rect 17302 6500 17306 6556
rect 17306 6500 17362 6556
rect 17362 6500 17366 6556
rect 17302 6496 17366 6500
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 3272 6012 3336 6016
rect 3272 5956 3276 6012
rect 3276 5956 3332 6012
rect 3332 5956 3336 6012
rect 3272 5952 3336 5956
rect 3352 6012 3416 6016
rect 3352 5956 3356 6012
rect 3356 5956 3412 6012
rect 3412 5956 3416 6012
rect 3352 5952 3416 5956
rect 6212 6012 6276 6016
rect 6212 5956 6216 6012
rect 6216 5956 6272 6012
rect 6272 5956 6276 6012
rect 6212 5952 6276 5956
rect 6292 6012 6356 6016
rect 6292 5956 6296 6012
rect 6296 5956 6352 6012
rect 6352 5956 6356 6012
rect 6292 5952 6356 5956
rect 6372 6012 6436 6016
rect 6372 5956 6376 6012
rect 6376 5956 6432 6012
rect 6432 5956 6436 6012
rect 6372 5952 6436 5956
rect 6452 6012 6516 6016
rect 6452 5956 6456 6012
rect 6456 5956 6512 6012
rect 6512 5956 6516 6012
rect 6452 5952 6516 5956
rect 9312 6012 9376 6016
rect 9312 5956 9316 6012
rect 9316 5956 9372 6012
rect 9372 5956 9376 6012
rect 9312 5952 9376 5956
rect 9392 6012 9456 6016
rect 9392 5956 9396 6012
rect 9396 5956 9452 6012
rect 9452 5956 9456 6012
rect 9392 5952 9456 5956
rect 9472 6012 9536 6016
rect 9472 5956 9476 6012
rect 9476 5956 9532 6012
rect 9532 5956 9536 6012
rect 9472 5952 9536 5956
rect 9552 6012 9616 6016
rect 9552 5956 9556 6012
rect 9556 5956 9612 6012
rect 9612 5956 9616 6012
rect 9552 5952 9616 5956
rect 12412 6012 12476 6016
rect 12412 5956 12416 6012
rect 12416 5956 12472 6012
rect 12472 5956 12476 6012
rect 12412 5952 12476 5956
rect 12492 6012 12556 6016
rect 12492 5956 12496 6012
rect 12496 5956 12552 6012
rect 12552 5956 12556 6012
rect 12492 5952 12556 5956
rect 12572 6012 12636 6016
rect 12572 5956 12576 6012
rect 12576 5956 12632 6012
rect 12632 5956 12636 6012
rect 12572 5952 12636 5956
rect 12652 6012 12716 6016
rect 12652 5956 12656 6012
rect 12656 5956 12712 6012
rect 12712 5956 12716 6012
rect 12652 5952 12716 5956
rect 15512 6012 15576 6016
rect 15512 5956 15516 6012
rect 15516 5956 15572 6012
rect 15572 5956 15576 6012
rect 15512 5952 15576 5956
rect 15592 6012 15656 6016
rect 15592 5956 15596 6012
rect 15596 5956 15652 6012
rect 15652 5956 15656 6012
rect 15592 5952 15656 5956
rect 15672 6012 15736 6016
rect 15672 5956 15676 6012
rect 15676 5956 15732 6012
rect 15732 5956 15736 6012
rect 15672 5952 15736 5956
rect 15752 6012 15816 6016
rect 15752 5956 15756 6012
rect 15756 5956 15812 6012
rect 15812 5956 15816 6012
rect 15752 5952 15816 5956
rect 4662 5468 4726 5472
rect 4662 5412 4666 5468
rect 4666 5412 4722 5468
rect 4722 5412 4726 5468
rect 4662 5408 4726 5412
rect 4742 5468 4806 5472
rect 4742 5412 4746 5468
rect 4746 5412 4802 5468
rect 4802 5412 4806 5468
rect 4742 5408 4806 5412
rect 4822 5468 4886 5472
rect 4822 5412 4826 5468
rect 4826 5412 4882 5468
rect 4882 5412 4886 5468
rect 4822 5408 4886 5412
rect 4902 5468 4966 5472
rect 4902 5412 4906 5468
rect 4906 5412 4962 5468
rect 4962 5412 4966 5468
rect 4902 5408 4966 5412
rect 7762 5468 7826 5472
rect 7762 5412 7766 5468
rect 7766 5412 7822 5468
rect 7822 5412 7826 5468
rect 7762 5408 7826 5412
rect 7842 5468 7906 5472
rect 7842 5412 7846 5468
rect 7846 5412 7902 5468
rect 7902 5412 7906 5468
rect 7842 5408 7906 5412
rect 7922 5468 7986 5472
rect 7922 5412 7926 5468
rect 7926 5412 7982 5468
rect 7982 5412 7986 5468
rect 7922 5408 7986 5412
rect 8002 5468 8066 5472
rect 8002 5412 8006 5468
rect 8006 5412 8062 5468
rect 8062 5412 8066 5468
rect 8002 5408 8066 5412
rect 10862 5468 10926 5472
rect 10862 5412 10866 5468
rect 10866 5412 10922 5468
rect 10922 5412 10926 5468
rect 10862 5408 10926 5412
rect 10942 5468 11006 5472
rect 10942 5412 10946 5468
rect 10946 5412 11002 5468
rect 11002 5412 11006 5468
rect 10942 5408 11006 5412
rect 11022 5468 11086 5472
rect 11022 5412 11026 5468
rect 11026 5412 11082 5468
rect 11082 5412 11086 5468
rect 11022 5408 11086 5412
rect 11102 5468 11166 5472
rect 11102 5412 11106 5468
rect 11106 5412 11162 5468
rect 11162 5412 11166 5468
rect 11102 5408 11166 5412
rect 13962 5468 14026 5472
rect 13962 5412 13966 5468
rect 13966 5412 14022 5468
rect 14022 5412 14026 5468
rect 13962 5408 14026 5412
rect 14042 5468 14106 5472
rect 14042 5412 14046 5468
rect 14046 5412 14102 5468
rect 14102 5412 14106 5468
rect 14042 5408 14106 5412
rect 14122 5468 14186 5472
rect 14122 5412 14126 5468
rect 14126 5412 14182 5468
rect 14182 5412 14186 5468
rect 14122 5408 14186 5412
rect 14202 5468 14266 5472
rect 14202 5412 14206 5468
rect 14206 5412 14262 5468
rect 14262 5412 14266 5468
rect 14202 5408 14266 5412
rect 17062 5468 17126 5472
rect 17062 5412 17066 5468
rect 17066 5412 17122 5468
rect 17122 5412 17126 5468
rect 17062 5408 17126 5412
rect 17142 5468 17206 5472
rect 17142 5412 17146 5468
rect 17146 5412 17202 5468
rect 17202 5412 17206 5468
rect 17142 5408 17206 5412
rect 17222 5468 17286 5472
rect 17222 5412 17226 5468
rect 17226 5412 17282 5468
rect 17282 5412 17286 5468
rect 17222 5408 17286 5412
rect 17302 5468 17366 5472
rect 17302 5412 17306 5468
rect 17306 5412 17362 5468
rect 17362 5412 17366 5468
rect 17302 5408 17366 5412
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 3272 4924 3336 4928
rect 3272 4868 3276 4924
rect 3276 4868 3332 4924
rect 3332 4868 3336 4924
rect 3272 4864 3336 4868
rect 3352 4924 3416 4928
rect 3352 4868 3356 4924
rect 3356 4868 3412 4924
rect 3412 4868 3416 4924
rect 3352 4864 3416 4868
rect 6212 4924 6276 4928
rect 6212 4868 6216 4924
rect 6216 4868 6272 4924
rect 6272 4868 6276 4924
rect 6212 4864 6276 4868
rect 6292 4924 6356 4928
rect 6292 4868 6296 4924
rect 6296 4868 6352 4924
rect 6352 4868 6356 4924
rect 6292 4864 6356 4868
rect 6372 4924 6436 4928
rect 6372 4868 6376 4924
rect 6376 4868 6432 4924
rect 6432 4868 6436 4924
rect 6372 4864 6436 4868
rect 6452 4924 6516 4928
rect 6452 4868 6456 4924
rect 6456 4868 6512 4924
rect 6512 4868 6516 4924
rect 6452 4864 6516 4868
rect 9312 4924 9376 4928
rect 9312 4868 9316 4924
rect 9316 4868 9372 4924
rect 9372 4868 9376 4924
rect 9312 4864 9376 4868
rect 9392 4924 9456 4928
rect 9392 4868 9396 4924
rect 9396 4868 9452 4924
rect 9452 4868 9456 4924
rect 9392 4864 9456 4868
rect 9472 4924 9536 4928
rect 9472 4868 9476 4924
rect 9476 4868 9532 4924
rect 9532 4868 9536 4924
rect 9472 4864 9536 4868
rect 9552 4924 9616 4928
rect 9552 4868 9556 4924
rect 9556 4868 9612 4924
rect 9612 4868 9616 4924
rect 9552 4864 9616 4868
rect 12412 4924 12476 4928
rect 12412 4868 12416 4924
rect 12416 4868 12472 4924
rect 12472 4868 12476 4924
rect 12412 4864 12476 4868
rect 12492 4924 12556 4928
rect 12492 4868 12496 4924
rect 12496 4868 12552 4924
rect 12552 4868 12556 4924
rect 12492 4864 12556 4868
rect 12572 4924 12636 4928
rect 12572 4868 12576 4924
rect 12576 4868 12632 4924
rect 12632 4868 12636 4924
rect 12572 4864 12636 4868
rect 12652 4924 12716 4928
rect 12652 4868 12656 4924
rect 12656 4868 12712 4924
rect 12712 4868 12716 4924
rect 12652 4864 12716 4868
rect 15512 4924 15576 4928
rect 15512 4868 15516 4924
rect 15516 4868 15572 4924
rect 15572 4868 15576 4924
rect 15512 4864 15576 4868
rect 15592 4924 15656 4928
rect 15592 4868 15596 4924
rect 15596 4868 15652 4924
rect 15652 4868 15656 4924
rect 15592 4864 15656 4868
rect 15672 4924 15736 4928
rect 15672 4868 15676 4924
rect 15676 4868 15732 4924
rect 15732 4868 15736 4924
rect 15672 4864 15736 4868
rect 15752 4924 15816 4928
rect 15752 4868 15756 4924
rect 15756 4868 15812 4924
rect 15812 4868 15816 4924
rect 15752 4864 15816 4868
rect 4662 4380 4726 4384
rect 4662 4324 4666 4380
rect 4666 4324 4722 4380
rect 4722 4324 4726 4380
rect 4662 4320 4726 4324
rect 4742 4380 4806 4384
rect 4742 4324 4746 4380
rect 4746 4324 4802 4380
rect 4802 4324 4806 4380
rect 4742 4320 4806 4324
rect 4822 4380 4886 4384
rect 4822 4324 4826 4380
rect 4826 4324 4882 4380
rect 4882 4324 4886 4380
rect 4822 4320 4886 4324
rect 4902 4380 4966 4384
rect 4902 4324 4906 4380
rect 4906 4324 4962 4380
rect 4962 4324 4966 4380
rect 4902 4320 4966 4324
rect 7762 4380 7826 4384
rect 7762 4324 7766 4380
rect 7766 4324 7822 4380
rect 7822 4324 7826 4380
rect 7762 4320 7826 4324
rect 7842 4380 7906 4384
rect 7842 4324 7846 4380
rect 7846 4324 7902 4380
rect 7902 4324 7906 4380
rect 7842 4320 7906 4324
rect 7922 4380 7986 4384
rect 7922 4324 7926 4380
rect 7926 4324 7982 4380
rect 7982 4324 7986 4380
rect 7922 4320 7986 4324
rect 8002 4380 8066 4384
rect 8002 4324 8006 4380
rect 8006 4324 8062 4380
rect 8062 4324 8066 4380
rect 8002 4320 8066 4324
rect 10862 4380 10926 4384
rect 10862 4324 10866 4380
rect 10866 4324 10922 4380
rect 10922 4324 10926 4380
rect 10862 4320 10926 4324
rect 10942 4380 11006 4384
rect 10942 4324 10946 4380
rect 10946 4324 11002 4380
rect 11002 4324 11006 4380
rect 10942 4320 11006 4324
rect 11022 4380 11086 4384
rect 11022 4324 11026 4380
rect 11026 4324 11082 4380
rect 11082 4324 11086 4380
rect 11022 4320 11086 4324
rect 11102 4380 11166 4384
rect 11102 4324 11106 4380
rect 11106 4324 11162 4380
rect 11162 4324 11166 4380
rect 11102 4320 11166 4324
rect 13962 4380 14026 4384
rect 13962 4324 13966 4380
rect 13966 4324 14022 4380
rect 14022 4324 14026 4380
rect 13962 4320 14026 4324
rect 14042 4380 14106 4384
rect 14042 4324 14046 4380
rect 14046 4324 14102 4380
rect 14102 4324 14106 4380
rect 14042 4320 14106 4324
rect 14122 4380 14186 4384
rect 14122 4324 14126 4380
rect 14126 4324 14182 4380
rect 14182 4324 14186 4380
rect 14122 4320 14186 4324
rect 14202 4380 14266 4384
rect 14202 4324 14206 4380
rect 14206 4324 14262 4380
rect 14262 4324 14266 4380
rect 14202 4320 14266 4324
rect 17062 4380 17126 4384
rect 17062 4324 17066 4380
rect 17066 4324 17122 4380
rect 17122 4324 17126 4380
rect 17062 4320 17126 4324
rect 17142 4380 17206 4384
rect 17142 4324 17146 4380
rect 17146 4324 17202 4380
rect 17202 4324 17206 4380
rect 17142 4320 17206 4324
rect 17222 4380 17286 4384
rect 17222 4324 17226 4380
rect 17226 4324 17282 4380
rect 17282 4324 17286 4380
rect 17222 4320 17286 4324
rect 17302 4380 17366 4384
rect 17302 4324 17306 4380
rect 17306 4324 17362 4380
rect 17362 4324 17366 4380
rect 17302 4320 17366 4324
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 3272 3836 3336 3840
rect 3272 3780 3276 3836
rect 3276 3780 3332 3836
rect 3332 3780 3336 3836
rect 3272 3776 3336 3780
rect 3352 3836 3416 3840
rect 3352 3780 3356 3836
rect 3356 3780 3412 3836
rect 3412 3780 3416 3836
rect 3352 3776 3416 3780
rect 6212 3836 6276 3840
rect 6212 3780 6216 3836
rect 6216 3780 6272 3836
rect 6272 3780 6276 3836
rect 6212 3776 6276 3780
rect 6292 3836 6356 3840
rect 6292 3780 6296 3836
rect 6296 3780 6352 3836
rect 6352 3780 6356 3836
rect 6292 3776 6356 3780
rect 6372 3836 6436 3840
rect 6372 3780 6376 3836
rect 6376 3780 6432 3836
rect 6432 3780 6436 3836
rect 6372 3776 6436 3780
rect 6452 3836 6516 3840
rect 6452 3780 6456 3836
rect 6456 3780 6512 3836
rect 6512 3780 6516 3836
rect 6452 3776 6516 3780
rect 9312 3836 9376 3840
rect 9312 3780 9316 3836
rect 9316 3780 9372 3836
rect 9372 3780 9376 3836
rect 9312 3776 9376 3780
rect 9392 3836 9456 3840
rect 9392 3780 9396 3836
rect 9396 3780 9452 3836
rect 9452 3780 9456 3836
rect 9392 3776 9456 3780
rect 9472 3836 9536 3840
rect 9472 3780 9476 3836
rect 9476 3780 9532 3836
rect 9532 3780 9536 3836
rect 9472 3776 9536 3780
rect 9552 3836 9616 3840
rect 9552 3780 9556 3836
rect 9556 3780 9612 3836
rect 9612 3780 9616 3836
rect 9552 3776 9616 3780
rect 12412 3836 12476 3840
rect 12412 3780 12416 3836
rect 12416 3780 12472 3836
rect 12472 3780 12476 3836
rect 12412 3776 12476 3780
rect 12492 3836 12556 3840
rect 12492 3780 12496 3836
rect 12496 3780 12552 3836
rect 12552 3780 12556 3836
rect 12492 3776 12556 3780
rect 12572 3836 12636 3840
rect 12572 3780 12576 3836
rect 12576 3780 12632 3836
rect 12632 3780 12636 3836
rect 12572 3776 12636 3780
rect 12652 3836 12716 3840
rect 12652 3780 12656 3836
rect 12656 3780 12712 3836
rect 12712 3780 12716 3836
rect 12652 3776 12716 3780
rect 15512 3836 15576 3840
rect 15512 3780 15516 3836
rect 15516 3780 15572 3836
rect 15572 3780 15576 3836
rect 15512 3776 15576 3780
rect 15592 3836 15656 3840
rect 15592 3780 15596 3836
rect 15596 3780 15652 3836
rect 15652 3780 15656 3836
rect 15592 3776 15656 3780
rect 15672 3836 15736 3840
rect 15672 3780 15676 3836
rect 15676 3780 15732 3836
rect 15732 3780 15736 3836
rect 15672 3776 15736 3780
rect 15752 3836 15816 3840
rect 15752 3780 15756 3836
rect 15756 3780 15812 3836
rect 15812 3780 15816 3836
rect 15752 3776 15816 3780
rect 4662 3292 4726 3296
rect 4662 3236 4666 3292
rect 4666 3236 4722 3292
rect 4722 3236 4726 3292
rect 4662 3232 4726 3236
rect 4742 3292 4806 3296
rect 4742 3236 4746 3292
rect 4746 3236 4802 3292
rect 4802 3236 4806 3292
rect 4742 3232 4806 3236
rect 4822 3292 4886 3296
rect 4822 3236 4826 3292
rect 4826 3236 4882 3292
rect 4882 3236 4886 3292
rect 4822 3232 4886 3236
rect 4902 3292 4966 3296
rect 4902 3236 4906 3292
rect 4906 3236 4962 3292
rect 4962 3236 4966 3292
rect 4902 3232 4966 3236
rect 7762 3292 7826 3296
rect 7762 3236 7766 3292
rect 7766 3236 7822 3292
rect 7822 3236 7826 3292
rect 7762 3232 7826 3236
rect 7842 3292 7906 3296
rect 7842 3236 7846 3292
rect 7846 3236 7902 3292
rect 7902 3236 7906 3292
rect 7842 3232 7906 3236
rect 7922 3292 7986 3296
rect 7922 3236 7926 3292
rect 7926 3236 7982 3292
rect 7982 3236 7986 3292
rect 7922 3232 7986 3236
rect 8002 3292 8066 3296
rect 8002 3236 8006 3292
rect 8006 3236 8062 3292
rect 8062 3236 8066 3292
rect 8002 3232 8066 3236
rect 10862 3292 10926 3296
rect 10862 3236 10866 3292
rect 10866 3236 10922 3292
rect 10922 3236 10926 3292
rect 10862 3232 10926 3236
rect 10942 3292 11006 3296
rect 10942 3236 10946 3292
rect 10946 3236 11002 3292
rect 11002 3236 11006 3292
rect 10942 3232 11006 3236
rect 11022 3292 11086 3296
rect 11022 3236 11026 3292
rect 11026 3236 11082 3292
rect 11082 3236 11086 3292
rect 11022 3232 11086 3236
rect 11102 3292 11166 3296
rect 11102 3236 11106 3292
rect 11106 3236 11162 3292
rect 11162 3236 11166 3292
rect 11102 3232 11166 3236
rect 13962 3292 14026 3296
rect 13962 3236 13966 3292
rect 13966 3236 14022 3292
rect 14022 3236 14026 3292
rect 13962 3232 14026 3236
rect 14042 3292 14106 3296
rect 14042 3236 14046 3292
rect 14046 3236 14102 3292
rect 14102 3236 14106 3292
rect 14042 3232 14106 3236
rect 14122 3292 14186 3296
rect 14122 3236 14126 3292
rect 14126 3236 14182 3292
rect 14182 3236 14186 3292
rect 14122 3232 14186 3236
rect 14202 3292 14266 3296
rect 14202 3236 14206 3292
rect 14206 3236 14262 3292
rect 14262 3236 14266 3292
rect 14202 3232 14266 3236
rect 17062 3292 17126 3296
rect 17062 3236 17066 3292
rect 17066 3236 17122 3292
rect 17122 3236 17126 3292
rect 17062 3232 17126 3236
rect 17142 3292 17206 3296
rect 17142 3236 17146 3292
rect 17146 3236 17202 3292
rect 17202 3236 17206 3292
rect 17142 3232 17206 3236
rect 17222 3292 17286 3296
rect 17222 3236 17226 3292
rect 17226 3236 17282 3292
rect 17282 3236 17286 3292
rect 17222 3232 17286 3236
rect 17302 3292 17366 3296
rect 17302 3236 17306 3292
rect 17306 3236 17362 3292
rect 17362 3236 17366 3292
rect 17302 3232 17366 3236
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 3272 2748 3336 2752
rect 3272 2692 3276 2748
rect 3276 2692 3332 2748
rect 3332 2692 3336 2748
rect 3272 2688 3336 2692
rect 3352 2748 3416 2752
rect 3352 2692 3356 2748
rect 3356 2692 3412 2748
rect 3412 2692 3416 2748
rect 3352 2688 3416 2692
rect 6212 2748 6276 2752
rect 6212 2692 6216 2748
rect 6216 2692 6272 2748
rect 6272 2692 6276 2748
rect 6212 2688 6276 2692
rect 6292 2748 6356 2752
rect 6292 2692 6296 2748
rect 6296 2692 6352 2748
rect 6352 2692 6356 2748
rect 6292 2688 6356 2692
rect 6372 2748 6436 2752
rect 6372 2692 6376 2748
rect 6376 2692 6432 2748
rect 6432 2692 6436 2748
rect 6372 2688 6436 2692
rect 6452 2748 6516 2752
rect 6452 2692 6456 2748
rect 6456 2692 6512 2748
rect 6512 2692 6516 2748
rect 6452 2688 6516 2692
rect 9312 2748 9376 2752
rect 9312 2692 9316 2748
rect 9316 2692 9372 2748
rect 9372 2692 9376 2748
rect 9312 2688 9376 2692
rect 9392 2748 9456 2752
rect 9392 2692 9396 2748
rect 9396 2692 9452 2748
rect 9452 2692 9456 2748
rect 9392 2688 9456 2692
rect 9472 2748 9536 2752
rect 9472 2692 9476 2748
rect 9476 2692 9532 2748
rect 9532 2692 9536 2748
rect 9472 2688 9536 2692
rect 9552 2748 9616 2752
rect 9552 2692 9556 2748
rect 9556 2692 9612 2748
rect 9612 2692 9616 2748
rect 9552 2688 9616 2692
rect 12412 2748 12476 2752
rect 12412 2692 12416 2748
rect 12416 2692 12472 2748
rect 12472 2692 12476 2748
rect 12412 2688 12476 2692
rect 12492 2748 12556 2752
rect 12492 2692 12496 2748
rect 12496 2692 12552 2748
rect 12552 2692 12556 2748
rect 12492 2688 12556 2692
rect 12572 2748 12636 2752
rect 12572 2692 12576 2748
rect 12576 2692 12632 2748
rect 12632 2692 12636 2748
rect 12572 2688 12636 2692
rect 12652 2748 12716 2752
rect 12652 2692 12656 2748
rect 12656 2692 12712 2748
rect 12712 2692 12716 2748
rect 12652 2688 12716 2692
rect 15512 2748 15576 2752
rect 15512 2692 15516 2748
rect 15516 2692 15572 2748
rect 15572 2692 15576 2748
rect 15512 2688 15576 2692
rect 15592 2748 15656 2752
rect 15592 2692 15596 2748
rect 15596 2692 15652 2748
rect 15652 2692 15656 2748
rect 15592 2688 15656 2692
rect 15672 2748 15736 2752
rect 15672 2692 15676 2748
rect 15676 2692 15732 2748
rect 15732 2692 15736 2748
rect 15672 2688 15736 2692
rect 15752 2748 15816 2752
rect 15752 2692 15756 2748
rect 15756 2692 15812 2748
rect 15812 2692 15816 2748
rect 15752 2688 15816 2692
rect 4662 2204 4726 2208
rect 4662 2148 4666 2204
rect 4666 2148 4722 2204
rect 4722 2148 4726 2204
rect 4662 2144 4726 2148
rect 4742 2204 4806 2208
rect 4742 2148 4746 2204
rect 4746 2148 4802 2204
rect 4802 2148 4806 2204
rect 4742 2144 4806 2148
rect 4822 2204 4886 2208
rect 4822 2148 4826 2204
rect 4826 2148 4882 2204
rect 4882 2148 4886 2204
rect 4822 2144 4886 2148
rect 4902 2204 4966 2208
rect 4902 2148 4906 2204
rect 4906 2148 4962 2204
rect 4962 2148 4966 2204
rect 4902 2144 4966 2148
rect 7762 2204 7826 2208
rect 7762 2148 7766 2204
rect 7766 2148 7822 2204
rect 7822 2148 7826 2204
rect 7762 2144 7826 2148
rect 7842 2204 7906 2208
rect 7842 2148 7846 2204
rect 7846 2148 7902 2204
rect 7902 2148 7906 2204
rect 7842 2144 7906 2148
rect 7922 2204 7986 2208
rect 7922 2148 7926 2204
rect 7926 2148 7982 2204
rect 7982 2148 7986 2204
rect 7922 2144 7986 2148
rect 8002 2204 8066 2208
rect 8002 2148 8006 2204
rect 8006 2148 8062 2204
rect 8062 2148 8066 2204
rect 8002 2144 8066 2148
rect 10862 2204 10926 2208
rect 10862 2148 10866 2204
rect 10866 2148 10922 2204
rect 10922 2148 10926 2204
rect 10862 2144 10926 2148
rect 10942 2204 11006 2208
rect 10942 2148 10946 2204
rect 10946 2148 11002 2204
rect 11002 2148 11006 2204
rect 10942 2144 11006 2148
rect 11022 2204 11086 2208
rect 11022 2148 11026 2204
rect 11026 2148 11082 2204
rect 11082 2148 11086 2204
rect 11022 2144 11086 2148
rect 11102 2204 11166 2208
rect 11102 2148 11106 2204
rect 11106 2148 11162 2204
rect 11162 2148 11166 2204
rect 11102 2144 11166 2148
rect 13962 2204 14026 2208
rect 13962 2148 13966 2204
rect 13966 2148 14022 2204
rect 14022 2148 14026 2204
rect 13962 2144 14026 2148
rect 14042 2204 14106 2208
rect 14042 2148 14046 2204
rect 14046 2148 14102 2204
rect 14102 2148 14106 2204
rect 14042 2144 14106 2148
rect 14122 2204 14186 2208
rect 14122 2148 14126 2204
rect 14126 2148 14182 2204
rect 14182 2148 14186 2204
rect 14122 2144 14186 2148
rect 14202 2204 14266 2208
rect 14202 2148 14206 2204
rect 14206 2148 14262 2204
rect 14262 2148 14266 2204
rect 14202 2144 14266 2148
rect 17062 2204 17126 2208
rect 17062 2148 17066 2204
rect 17066 2148 17122 2204
rect 17122 2148 17126 2204
rect 17062 2144 17126 2148
rect 17142 2204 17206 2208
rect 17142 2148 17146 2204
rect 17146 2148 17202 2204
rect 17202 2148 17206 2204
rect 17142 2144 17206 2148
rect 17222 2204 17286 2208
rect 17222 2148 17226 2204
rect 17226 2148 17282 2204
rect 17282 2148 17286 2204
rect 17222 2144 17286 2148
rect 17302 2204 17366 2208
rect 17302 2148 17306 2204
rect 17306 2148 17362 2204
rect 17362 2148 17366 2204
rect 17302 2144 17366 2148
rect 3112 1660 3176 1664
rect 3112 1604 3116 1660
rect 3116 1604 3172 1660
rect 3172 1604 3176 1660
rect 3112 1600 3176 1604
rect 3192 1660 3256 1664
rect 3192 1604 3196 1660
rect 3196 1604 3252 1660
rect 3252 1604 3256 1660
rect 3192 1600 3256 1604
rect 3272 1660 3336 1664
rect 3272 1604 3276 1660
rect 3276 1604 3332 1660
rect 3332 1604 3336 1660
rect 3272 1600 3336 1604
rect 3352 1660 3416 1664
rect 3352 1604 3356 1660
rect 3356 1604 3412 1660
rect 3412 1604 3416 1660
rect 3352 1600 3416 1604
rect 6212 1660 6276 1664
rect 6212 1604 6216 1660
rect 6216 1604 6272 1660
rect 6272 1604 6276 1660
rect 6212 1600 6276 1604
rect 6292 1660 6356 1664
rect 6292 1604 6296 1660
rect 6296 1604 6352 1660
rect 6352 1604 6356 1660
rect 6292 1600 6356 1604
rect 6372 1660 6436 1664
rect 6372 1604 6376 1660
rect 6376 1604 6432 1660
rect 6432 1604 6436 1660
rect 6372 1600 6436 1604
rect 6452 1660 6516 1664
rect 6452 1604 6456 1660
rect 6456 1604 6512 1660
rect 6512 1604 6516 1660
rect 6452 1600 6516 1604
rect 9312 1660 9376 1664
rect 9312 1604 9316 1660
rect 9316 1604 9372 1660
rect 9372 1604 9376 1660
rect 9312 1600 9376 1604
rect 9392 1660 9456 1664
rect 9392 1604 9396 1660
rect 9396 1604 9452 1660
rect 9452 1604 9456 1660
rect 9392 1600 9456 1604
rect 9472 1660 9536 1664
rect 9472 1604 9476 1660
rect 9476 1604 9532 1660
rect 9532 1604 9536 1660
rect 9472 1600 9536 1604
rect 9552 1660 9616 1664
rect 9552 1604 9556 1660
rect 9556 1604 9612 1660
rect 9612 1604 9616 1660
rect 9552 1600 9616 1604
rect 12412 1660 12476 1664
rect 12412 1604 12416 1660
rect 12416 1604 12472 1660
rect 12472 1604 12476 1660
rect 12412 1600 12476 1604
rect 12492 1660 12556 1664
rect 12492 1604 12496 1660
rect 12496 1604 12552 1660
rect 12552 1604 12556 1660
rect 12492 1600 12556 1604
rect 12572 1660 12636 1664
rect 12572 1604 12576 1660
rect 12576 1604 12632 1660
rect 12632 1604 12636 1660
rect 12572 1600 12636 1604
rect 12652 1660 12716 1664
rect 12652 1604 12656 1660
rect 12656 1604 12712 1660
rect 12712 1604 12716 1660
rect 12652 1600 12716 1604
rect 15512 1660 15576 1664
rect 15512 1604 15516 1660
rect 15516 1604 15572 1660
rect 15572 1604 15576 1660
rect 15512 1600 15576 1604
rect 15592 1660 15656 1664
rect 15592 1604 15596 1660
rect 15596 1604 15652 1660
rect 15652 1604 15656 1660
rect 15592 1600 15656 1604
rect 15672 1660 15736 1664
rect 15672 1604 15676 1660
rect 15676 1604 15732 1660
rect 15732 1604 15736 1660
rect 15672 1600 15736 1604
rect 15752 1660 15816 1664
rect 15752 1604 15756 1660
rect 15756 1604 15812 1660
rect 15812 1604 15816 1660
rect 15752 1600 15816 1604
rect 4662 1116 4726 1120
rect 4662 1060 4666 1116
rect 4666 1060 4722 1116
rect 4722 1060 4726 1116
rect 4662 1056 4726 1060
rect 4742 1116 4806 1120
rect 4742 1060 4746 1116
rect 4746 1060 4802 1116
rect 4802 1060 4806 1116
rect 4742 1056 4806 1060
rect 4822 1116 4886 1120
rect 4822 1060 4826 1116
rect 4826 1060 4882 1116
rect 4882 1060 4886 1116
rect 4822 1056 4886 1060
rect 4902 1116 4966 1120
rect 4902 1060 4906 1116
rect 4906 1060 4962 1116
rect 4962 1060 4966 1116
rect 4902 1056 4966 1060
rect 7762 1116 7826 1120
rect 7762 1060 7766 1116
rect 7766 1060 7822 1116
rect 7822 1060 7826 1116
rect 7762 1056 7826 1060
rect 7842 1116 7906 1120
rect 7842 1060 7846 1116
rect 7846 1060 7902 1116
rect 7902 1060 7906 1116
rect 7842 1056 7906 1060
rect 7922 1116 7986 1120
rect 7922 1060 7926 1116
rect 7926 1060 7982 1116
rect 7982 1060 7986 1116
rect 7922 1056 7986 1060
rect 8002 1116 8066 1120
rect 8002 1060 8006 1116
rect 8006 1060 8062 1116
rect 8062 1060 8066 1116
rect 8002 1056 8066 1060
rect 10862 1116 10926 1120
rect 10862 1060 10866 1116
rect 10866 1060 10922 1116
rect 10922 1060 10926 1116
rect 10862 1056 10926 1060
rect 10942 1116 11006 1120
rect 10942 1060 10946 1116
rect 10946 1060 11002 1116
rect 11002 1060 11006 1116
rect 10942 1056 11006 1060
rect 11022 1116 11086 1120
rect 11022 1060 11026 1116
rect 11026 1060 11082 1116
rect 11082 1060 11086 1116
rect 11022 1056 11086 1060
rect 11102 1116 11166 1120
rect 11102 1060 11106 1116
rect 11106 1060 11162 1116
rect 11162 1060 11166 1116
rect 11102 1056 11166 1060
rect 13962 1116 14026 1120
rect 13962 1060 13966 1116
rect 13966 1060 14022 1116
rect 14022 1060 14026 1116
rect 13962 1056 14026 1060
rect 14042 1116 14106 1120
rect 14042 1060 14046 1116
rect 14046 1060 14102 1116
rect 14102 1060 14106 1116
rect 14042 1056 14106 1060
rect 14122 1116 14186 1120
rect 14122 1060 14126 1116
rect 14126 1060 14182 1116
rect 14182 1060 14186 1116
rect 14122 1056 14186 1060
rect 14202 1116 14266 1120
rect 14202 1060 14206 1116
rect 14206 1060 14262 1116
rect 14262 1060 14266 1116
rect 14202 1056 14266 1060
rect 17062 1116 17126 1120
rect 17062 1060 17066 1116
rect 17066 1060 17122 1116
rect 17122 1060 17126 1116
rect 17062 1056 17126 1060
rect 17142 1116 17206 1120
rect 17142 1060 17146 1116
rect 17146 1060 17202 1116
rect 17202 1060 17206 1116
rect 17142 1056 17206 1060
rect 17222 1116 17286 1120
rect 17222 1060 17226 1116
rect 17226 1060 17282 1116
rect 17282 1060 17286 1116
rect 17222 1056 17286 1060
rect 17302 1116 17366 1120
rect 17302 1060 17306 1116
rect 17306 1060 17362 1116
rect 17362 1060 17366 1116
rect 17302 1056 17366 1060
rect 3112 572 3176 576
rect 3112 516 3116 572
rect 3116 516 3172 572
rect 3172 516 3176 572
rect 3112 512 3176 516
rect 3192 572 3256 576
rect 3192 516 3196 572
rect 3196 516 3252 572
rect 3252 516 3256 572
rect 3192 512 3256 516
rect 3272 572 3336 576
rect 3272 516 3276 572
rect 3276 516 3332 572
rect 3332 516 3336 572
rect 3272 512 3336 516
rect 3352 572 3416 576
rect 3352 516 3356 572
rect 3356 516 3412 572
rect 3412 516 3416 572
rect 3352 512 3416 516
rect 6212 572 6276 576
rect 6212 516 6216 572
rect 6216 516 6272 572
rect 6272 516 6276 572
rect 6212 512 6276 516
rect 6292 572 6356 576
rect 6292 516 6296 572
rect 6296 516 6352 572
rect 6352 516 6356 572
rect 6292 512 6356 516
rect 6372 572 6436 576
rect 6372 516 6376 572
rect 6376 516 6432 572
rect 6432 516 6436 572
rect 6372 512 6436 516
rect 6452 572 6516 576
rect 6452 516 6456 572
rect 6456 516 6512 572
rect 6512 516 6516 572
rect 6452 512 6516 516
rect 9312 572 9376 576
rect 9312 516 9316 572
rect 9316 516 9372 572
rect 9372 516 9376 572
rect 9312 512 9376 516
rect 9392 572 9456 576
rect 9392 516 9396 572
rect 9396 516 9452 572
rect 9452 516 9456 572
rect 9392 512 9456 516
rect 9472 572 9536 576
rect 9472 516 9476 572
rect 9476 516 9532 572
rect 9532 516 9536 572
rect 9472 512 9536 516
rect 9552 572 9616 576
rect 9552 516 9556 572
rect 9556 516 9612 572
rect 9612 516 9616 572
rect 9552 512 9616 516
rect 12412 572 12476 576
rect 12412 516 12416 572
rect 12416 516 12472 572
rect 12472 516 12476 572
rect 12412 512 12476 516
rect 12492 572 12556 576
rect 12492 516 12496 572
rect 12496 516 12552 572
rect 12552 516 12556 572
rect 12492 512 12556 516
rect 12572 572 12636 576
rect 12572 516 12576 572
rect 12576 516 12632 572
rect 12632 516 12636 572
rect 12572 512 12636 516
rect 12652 572 12716 576
rect 12652 516 12656 572
rect 12656 516 12712 572
rect 12712 516 12716 572
rect 12652 512 12716 516
rect 15512 572 15576 576
rect 15512 516 15516 572
rect 15516 516 15572 572
rect 15572 516 15576 572
rect 15512 512 15576 516
rect 15592 572 15656 576
rect 15592 516 15596 572
rect 15596 516 15652 572
rect 15652 516 15656 572
rect 15592 512 15656 516
rect 15672 572 15736 576
rect 15672 516 15676 572
rect 15676 516 15732 572
rect 15732 516 15736 572
rect 15672 512 15736 516
rect 15752 572 15816 576
rect 15752 516 15756 572
rect 15756 516 15812 572
rect 15812 516 15816 572
rect 15752 512 15816 516
rect 4662 28 4726 32
rect 4662 -28 4666 28
rect 4666 -28 4722 28
rect 4722 -28 4726 28
rect 4662 -32 4726 -28
rect 4742 28 4806 32
rect 4742 -28 4746 28
rect 4746 -28 4802 28
rect 4802 -28 4806 28
rect 4742 -32 4806 -28
rect 4822 28 4886 32
rect 4822 -28 4826 28
rect 4826 -28 4882 28
rect 4882 -28 4886 28
rect 4822 -32 4886 -28
rect 4902 28 4966 32
rect 4902 -28 4906 28
rect 4906 -28 4962 28
rect 4962 -28 4966 28
rect 4902 -32 4966 -28
rect 7762 28 7826 32
rect 7762 -28 7766 28
rect 7766 -28 7822 28
rect 7822 -28 7826 28
rect 7762 -32 7826 -28
rect 7842 28 7906 32
rect 7842 -28 7846 28
rect 7846 -28 7902 28
rect 7902 -28 7906 28
rect 7842 -32 7906 -28
rect 7922 28 7986 32
rect 7922 -28 7926 28
rect 7926 -28 7982 28
rect 7982 -28 7986 28
rect 7922 -32 7986 -28
rect 8002 28 8066 32
rect 8002 -28 8006 28
rect 8006 -28 8062 28
rect 8062 -28 8066 28
rect 8002 -32 8066 -28
rect 10862 28 10926 32
rect 10862 -28 10866 28
rect 10866 -28 10922 28
rect 10922 -28 10926 28
rect 10862 -32 10926 -28
rect 10942 28 11006 32
rect 10942 -28 10946 28
rect 10946 -28 11002 28
rect 11002 -28 11006 28
rect 10942 -32 11006 -28
rect 11022 28 11086 32
rect 11022 -28 11026 28
rect 11026 -28 11082 28
rect 11082 -28 11086 28
rect 11022 -32 11086 -28
rect 11102 28 11166 32
rect 11102 -28 11106 28
rect 11106 -28 11162 28
rect 11162 -28 11166 28
rect 11102 -32 11166 -28
rect 13962 28 14026 32
rect 13962 -28 13966 28
rect 13966 -28 14022 28
rect 14022 -28 14026 28
rect 13962 -32 14026 -28
rect 14042 28 14106 32
rect 14042 -28 14046 28
rect 14046 -28 14102 28
rect 14102 -28 14106 28
rect 14042 -32 14106 -28
rect 14122 28 14186 32
rect 14122 -28 14126 28
rect 14126 -28 14182 28
rect 14182 -28 14186 28
rect 14122 -32 14186 -28
rect 14202 28 14266 32
rect 14202 -28 14206 28
rect 14206 -28 14262 28
rect 14262 -28 14266 28
rect 14202 -32 14266 -28
rect 17062 28 17126 32
rect 17062 -28 17066 28
rect 17066 -28 17122 28
rect 17122 -28 17126 28
rect 17062 -32 17126 -28
rect 17142 28 17206 32
rect 17142 -28 17146 28
rect 17146 -28 17202 28
rect 17202 -28 17206 28
rect 17142 -32 17206 -28
rect 17222 28 17286 32
rect 17222 -28 17226 28
rect 17226 -28 17282 28
rect 17282 -28 17286 28
rect 17222 -32 17286 -28
rect 17302 28 17366 32
rect 17302 -28 17306 28
rect 17306 -28 17362 28
rect 17362 -28 17366 28
rect 17302 -32 17366 -28
<< metal4 >>
rect 3104 10368 3424 10928
rect 3104 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3272 10368
rect 3336 10304 3352 10368
rect 3416 10304 3424 10368
rect 3104 10160 3424 10304
rect 3104 9924 3146 10160
rect 3382 9924 3424 10160
rect 3104 9280 3424 9924
rect 3104 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3272 9280
rect 3336 9216 3352 9280
rect 3416 9216 3424 9280
rect 3104 8192 3424 9216
rect 3104 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3272 8192
rect 3336 8128 3352 8192
rect 3416 8128 3424 8192
rect 3104 7104 3424 8128
rect 3104 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3272 7104
rect 3336 7040 3352 7104
rect 3416 7040 3424 7104
rect 3104 6780 3424 7040
rect 3104 6544 3146 6780
rect 3382 6544 3424 6780
rect 3104 6016 3424 6544
rect 3104 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3272 6016
rect 3336 5952 3352 6016
rect 3416 5952 3424 6016
rect 3104 4928 3424 5952
rect 3104 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3272 4928
rect 3336 4864 3352 4928
rect 3416 4864 3424 4928
rect 3104 3840 3424 4864
rect 3104 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3272 3840
rect 3336 3776 3352 3840
rect 3416 3776 3424 3840
rect 3104 3400 3424 3776
rect 3104 3164 3146 3400
rect 3382 3164 3424 3400
rect 3104 2752 3424 3164
rect 3104 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3272 2752
rect 3336 2688 3352 2752
rect 3416 2688 3424 2752
rect 3104 1664 3424 2688
rect 3104 1600 3112 1664
rect 3176 1600 3192 1664
rect 3256 1600 3272 1664
rect 3336 1600 3352 1664
rect 3416 1600 3424 1664
rect 3104 576 3424 1600
rect 3104 512 3112 576
rect 3176 512 3192 576
rect 3256 512 3272 576
rect 3336 512 3352 576
rect 3416 512 3424 576
rect 3104 -48 3424 512
rect 4654 10912 4974 10928
rect 4654 10848 4662 10912
rect 4726 10848 4742 10912
rect 4806 10848 4822 10912
rect 4886 10848 4902 10912
rect 4966 10848 4974 10912
rect 4654 9824 4974 10848
rect 4654 9760 4662 9824
rect 4726 9760 4742 9824
rect 4806 9760 4822 9824
rect 4886 9760 4902 9824
rect 4966 9760 4974 9824
rect 4654 8736 4974 9760
rect 4654 8672 4662 8736
rect 4726 8672 4742 8736
rect 4806 8672 4822 8736
rect 4886 8672 4902 8736
rect 4966 8672 4974 8736
rect 4654 8470 4974 8672
rect 4654 8234 4696 8470
rect 4932 8234 4974 8470
rect 4654 7648 4974 8234
rect 4654 7584 4662 7648
rect 4726 7584 4742 7648
rect 4806 7584 4822 7648
rect 4886 7584 4902 7648
rect 4966 7584 4974 7648
rect 4654 6560 4974 7584
rect 4654 6496 4662 6560
rect 4726 6496 4742 6560
rect 4806 6496 4822 6560
rect 4886 6496 4902 6560
rect 4966 6496 4974 6560
rect 4654 5472 4974 6496
rect 4654 5408 4662 5472
rect 4726 5408 4742 5472
rect 4806 5408 4822 5472
rect 4886 5408 4902 5472
rect 4966 5408 4974 5472
rect 4654 5090 4974 5408
rect 4654 4854 4696 5090
rect 4932 4854 4974 5090
rect 4654 4384 4974 4854
rect 4654 4320 4662 4384
rect 4726 4320 4742 4384
rect 4806 4320 4822 4384
rect 4886 4320 4902 4384
rect 4966 4320 4974 4384
rect 4654 3296 4974 4320
rect 4654 3232 4662 3296
rect 4726 3232 4742 3296
rect 4806 3232 4822 3296
rect 4886 3232 4902 3296
rect 4966 3232 4974 3296
rect 4654 2208 4974 3232
rect 4654 2144 4662 2208
rect 4726 2144 4742 2208
rect 4806 2144 4822 2208
rect 4886 2144 4902 2208
rect 4966 2144 4974 2208
rect 4654 1120 4974 2144
rect 4654 1056 4662 1120
rect 4726 1056 4742 1120
rect 4806 1056 4822 1120
rect 4886 1056 4902 1120
rect 4966 1056 4974 1120
rect 4654 32 4974 1056
rect 4654 -32 4662 32
rect 4726 -32 4742 32
rect 4806 -32 4822 32
rect 4886 -32 4902 32
rect 4966 -32 4974 32
rect 4654 -48 4974 -32
rect 6204 10368 6524 10928
rect 6204 10304 6212 10368
rect 6276 10304 6292 10368
rect 6356 10304 6372 10368
rect 6436 10304 6452 10368
rect 6516 10304 6524 10368
rect 6204 10160 6524 10304
rect 6204 9924 6246 10160
rect 6482 9924 6524 10160
rect 6204 9280 6524 9924
rect 6204 9216 6212 9280
rect 6276 9216 6292 9280
rect 6356 9216 6372 9280
rect 6436 9216 6452 9280
rect 6516 9216 6524 9280
rect 6204 8192 6524 9216
rect 6204 8128 6212 8192
rect 6276 8128 6292 8192
rect 6356 8128 6372 8192
rect 6436 8128 6452 8192
rect 6516 8128 6524 8192
rect 6204 7104 6524 8128
rect 6204 7040 6212 7104
rect 6276 7040 6292 7104
rect 6356 7040 6372 7104
rect 6436 7040 6452 7104
rect 6516 7040 6524 7104
rect 6204 6780 6524 7040
rect 6204 6544 6246 6780
rect 6482 6544 6524 6780
rect 6204 6016 6524 6544
rect 6204 5952 6212 6016
rect 6276 5952 6292 6016
rect 6356 5952 6372 6016
rect 6436 5952 6452 6016
rect 6516 5952 6524 6016
rect 6204 4928 6524 5952
rect 6204 4864 6212 4928
rect 6276 4864 6292 4928
rect 6356 4864 6372 4928
rect 6436 4864 6452 4928
rect 6516 4864 6524 4928
rect 6204 3840 6524 4864
rect 6204 3776 6212 3840
rect 6276 3776 6292 3840
rect 6356 3776 6372 3840
rect 6436 3776 6452 3840
rect 6516 3776 6524 3840
rect 6204 3400 6524 3776
rect 6204 3164 6246 3400
rect 6482 3164 6524 3400
rect 6204 2752 6524 3164
rect 6204 2688 6212 2752
rect 6276 2688 6292 2752
rect 6356 2688 6372 2752
rect 6436 2688 6452 2752
rect 6516 2688 6524 2752
rect 6204 1664 6524 2688
rect 6204 1600 6212 1664
rect 6276 1600 6292 1664
rect 6356 1600 6372 1664
rect 6436 1600 6452 1664
rect 6516 1600 6524 1664
rect 6204 576 6524 1600
rect 6204 512 6212 576
rect 6276 512 6292 576
rect 6356 512 6372 576
rect 6436 512 6452 576
rect 6516 512 6524 576
rect 6204 -48 6524 512
rect 7754 10912 8074 10928
rect 7754 10848 7762 10912
rect 7826 10848 7842 10912
rect 7906 10848 7922 10912
rect 7986 10848 8002 10912
rect 8066 10848 8074 10912
rect 7754 9824 8074 10848
rect 7754 9760 7762 9824
rect 7826 9760 7842 9824
rect 7906 9760 7922 9824
rect 7986 9760 8002 9824
rect 8066 9760 8074 9824
rect 7754 8736 8074 9760
rect 7754 8672 7762 8736
rect 7826 8672 7842 8736
rect 7906 8672 7922 8736
rect 7986 8672 8002 8736
rect 8066 8672 8074 8736
rect 7754 8470 8074 8672
rect 7754 8234 7796 8470
rect 8032 8234 8074 8470
rect 7754 7648 8074 8234
rect 7754 7584 7762 7648
rect 7826 7584 7842 7648
rect 7906 7584 7922 7648
rect 7986 7584 8002 7648
rect 8066 7584 8074 7648
rect 7754 6560 8074 7584
rect 7754 6496 7762 6560
rect 7826 6496 7842 6560
rect 7906 6496 7922 6560
rect 7986 6496 8002 6560
rect 8066 6496 8074 6560
rect 7754 5472 8074 6496
rect 7754 5408 7762 5472
rect 7826 5408 7842 5472
rect 7906 5408 7922 5472
rect 7986 5408 8002 5472
rect 8066 5408 8074 5472
rect 7754 5090 8074 5408
rect 7754 4854 7796 5090
rect 8032 4854 8074 5090
rect 7754 4384 8074 4854
rect 7754 4320 7762 4384
rect 7826 4320 7842 4384
rect 7906 4320 7922 4384
rect 7986 4320 8002 4384
rect 8066 4320 8074 4384
rect 7754 3296 8074 4320
rect 7754 3232 7762 3296
rect 7826 3232 7842 3296
rect 7906 3232 7922 3296
rect 7986 3232 8002 3296
rect 8066 3232 8074 3296
rect 7754 2208 8074 3232
rect 7754 2144 7762 2208
rect 7826 2144 7842 2208
rect 7906 2144 7922 2208
rect 7986 2144 8002 2208
rect 8066 2144 8074 2208
rect 7754 1120 8074 2144
rect 7754 1056 7762 1120
rect 7826 1056 7842 1120
rect 7906 1056 7922 1120
rect 7986 1056 8002 1120
rect 8066 1056 8074 1120
rect 7754 32 8074 1056
rect 7754 -32 7762 32
rect 7826 -32 7842 32
rect 7906 -32 7922 32
rect 7986 -32 8002 32
rect 8066 -32 8074 32
rect 7754 -48 8074 -32
rect 9304 10368 9624 10928
rect 9304 10304 9312 10368
rect 9376 10304 9392 10368
rect 9456 10304 9472 10368
rect 9536 10304 9552 10368
rect 9616 10304 9624 10368
rect 9304 10160 9624 10304
rect 9304 9924 9346 10160
rect 9582 9924 9624 10160
rect 9304 9280 9624 9924
rect 9304 9216 9312 9280
rect 9376 9216 9392 9280
rect 9456 9216 9472 9280
rect 9536 9216 9552 9280
rect 9616 9216 9624 9280
rect 9304 8192 9624 9216
rect 9304 8128 9312 8192
rect 9376 8128 9392 8192
rect 9456 8128 9472 8192
rect 9536 8128 9552 8192
rect 9616 8128 9624 8192
rect 9304 7104 9624 8128
rect 9304 7040 9312 7104
rect 9376 7040 9392 7104
rect 9456 7040 9472 7104
rect 9536 7040 9552 7104
rect 9616 7040 9624 7104
rect 9304 6780 9624 7040
rect 9304 6544 9346 6780
rect 9582 6544 9624 6780
rect 9304 6016 9624 6544
rect 9304 5952 9312 6016
rect 9376 5952 9392 6016
rect 9456 5952 9472 6016
rect 9536 5952 9552 6016
rect 9616 5952 9624 6016
rect 9304 4928 9624 5952
rect 9304 4864 9312 4928
rect 9376 4864 9392 4928
rect 9456 4864 9472 4928
rect 9536 4864 9552 4928
rect 9616 4864 9624 4928
rect 9304 3840 9624 4864
rect 9304 3776 9312 3840
rect 9376 3776 9392 3840
rect 9456 3776 9472 3840
rect 9536 3776 9552 3840
rect 9616 3776 9624 3840
rect 9304 3400 9624 3776
rect 9304 3164 9346 3400
rect 9582 3164 9624 3400
rect 9304 2752 9624 3164
rect 9304 2688 9312 2752
rect 9376 2688 9392 2752
rect 9456 2688 9472 2752
rect 9536 2688 9552 2752
rect 9616 2688 9624 2752
rect 9304 1664 9624 2688
rect 9304 1600 9312 1664
rect 9376 1600 9392 1664
rect 9456 1600 9472 1664
rect 9536 1600 9552 1664
rect 9616 1600 9624 1664
rect 9304 576 9624 1600
rect 9304 512 9312 576
rect 9376 512 9392 576
rect 9456 512 9472 576
rect 9536 512 9552 576
rect 9616 512 9624 576
rect 9304 -48 9624 512
rect 10854 10912 11174 10928
rect 10854 10848 10862 10912
rect 10926 10848 10942 10912
rect 11006 10848 11022 10912
rect 11086 10848 11102 10912
rect 11166 10848 11174 10912
rect 10854 9824 11174 10848
rect 10854 9760 10862 9824
rect 10926 9760 10942 9824
rect 11006 9760 11022 9824
rect 11086 9760 11102 9824
rect 11166 9760 11174 9824
rect 10854 8736 11174 9760
rect 10854 8672 10862 8736
rect 10926 8672 10942 8736
rect 11006 8672 11022 8736
rect 11086 8672 11102 8736
rect 11166 8672 11174 8736
rect 10854 8470 11174 8672
rect 10854 8234 10896 8470
rect 11132 8234 11174 8470
rect 10854 7648 11174 8234
rect 10854 7584 10862 7648
rect 10926 7584 10942 7648
rect 11006 7584 11022 7648
rect 11086 7584 11102 7648
rect 11166 7584 11174 7648
rect 10854 6560 11174 7584
rect 10854 6496 10862 6560
rect 10926 6496 10942 6560
rect 11006 6496 11022 6560
rect 11086 6496 11102 6560
rect 11166 6496 11174 6560
rect 10854 5472 11174 6496
rect 10854 5408 10862 5472
rect 10926 5408 10942 5472
rect 11006 5408 11022 5472
rect 11086 5408 11102 5472
rect 11166 5408 11174 5472
rect 10854 5090 11174 5408
rect 10854 4854 10896 5090
rect 11132 4854 11174 5090
rect 10854 4384 11174 4854
rect 10854 4320 10862 4384
rect 10926 4320 10942 4384
rect 11006 4320 11022 4384
rect 11086 4320 11102 4384
rect 11166 4320 11174 4384
rect 10854 3296 11174 4320
rect 10854 3232 10862 3296
rect 10926 3232 10942 3296
rect 11006 3232 11022 3296
rect 11086 3232 11102 3296
rect 11166 3232 11174 3296
rect 10854 2208 11174 3232
rect 10854 2144 10862 2208
rect 10926 2144 10942 2208
rect 11006 2144 11022 2208
rect 11086 2144 11102 2208
rect 11166 2144 11174 2208
rect 10854 1120 11174 2144
rect 10854 1056 10862 1120
rect 10926 1056 10942 1120
rect 11006 1056 11022 1120
rect 11086 1056 11102 1120
rect 11166 1056 11174 1120
rect 10854 32 11174 1056
rect 10854 -32 10862 32
rect 10926 -32 10942 32
rect 11006 -32 11022 32
rect 11086 -32 11102 32
rect 11166 -32 11174 32
rect 10854 -48 11174 -32
rect 12404 10368 12724 10928
rect 12404 10304 12412 10368
rect 12476 10304 12492 10368
rect 12556 10304 12572 10368
rect 12636 10304 12652 10368
rect 12716 10304 12724 10368
rect 12404 10160 12724 10304
rect 12404 9924 12446 10160
rect 12682 9924 12724 10160
rect 12404 9280 12724 9924
rect 12404 9216 12412 9280
rect 12476 9216 12492 9280
rect 12556 9216 12572 9280
rect 12636 9216 12652 9280
rect 12716 9216 12724 9280
rect 12404 8192 12724 9216
rect 12404 8128 12412 8192
rect 12476 8128 12492 8192
rect 12556 8128 12572 8192
rect 12636 8128 12652 8192
rect 12716 8128 12724 8192
rect 12404 7104 12724 8128
rect 12404 7040 12412 7104
rect 12476 7040 12492 7104
rect 12556 7040 12572 7104
rect 12636 7040 12652 7104
rect 12716 7040 12724 7104
rect 12404 6780 12724 7040
rect 12404 6544 12446 6780
rect 12682 6544 12724 6780
rect 12404 6016 12724 6544
rect 12404 5952 12412 6016
rect 12476 5952 12492 6016
rect 12556 5952 12572 6016
rect 12636 5952 12652 6016
rect 12716 5952 12724 6016
rect 12404 4928 12724 5952
rect 12404 4864 12412 4928
rect 12476 4864 12492 4928
rect 12556 4864 12572 4928
rect 12636 4864 12652 4928
rect 12716 4864 12724 4928
rect 12404 3840 12724 4864
rect 12404 3776 12412 3840
rect 12476 3776 12492 3840
rect 12556 3776 12572 3840
rect 12636 3776 12652 3840
rect 12716 3776 12724 3840
rect 12404 3400 12724 3776
rect 12404 3164 12446 3400
rect 12682 3164 12724 3400
rect 12404 2752 12724 3164
rect 12404 2688 12412 2752
rect 12476 2688 12492 2752
rect 12556 2688 12572 2752
rect 12636 2688 12652 2752
rect 12716 2688 12724 2752
rect 12404 1664 12724 2688
rect 12404 1600 12412 1664
rect 12476 1600 12492 1664
rect 12556 1600 12572 1664
rect 12636 1600 12652 1664
rect 12716 1600 12724 1664
rect 12404 576 12724 1600
rect 12404 512 12412 576
rect 12476 512 12492 576
rect 12556 512 12572 576
rect 12636 512 12652 576
rect 12716 512 12724 576
rect 12404 -48 12724 512
rect 13954 10912 14274 10928
rect 13954 10848 13962 10912
rect 14026 10848 14042 10912
rect 14106 10848 14122 10912
rect 14186 10848 14202 10912
rect 14266 10848 14274 10912
rect 13954 9824 14274 10848
rect 13954 9760 13962 9824
rect 14026 9760 14042 9824
rect 14106 9760 14122 9824
rect 14186 9760 14202 9824
rect 14266 9760 14274 9824
rect 13954 8736 14274 9760
rect 13954 8672 13962 8736
rect 14026 8672 14042 8736
rect 14106 8672 14122 8736
rect 14186 8672 14202 8736
rect 14266 8672 14274 8736
rect 13954 8470 14274 8672
rect 13954 8234 13996 8470
rect 14232 8234 14274 8470
rect 13954 7648 14274 8234
rect 13954 7584 13962 7648
rect 14026 7584 14042 7648
rect 14106 7584 14122 7648
rect 14186 7584 14202 7648
rect 14266 7584 14274 7648
rect 13954 6560 14274 7584
rect 13954 6496 13962 6560
rect 14026 6496 14042 6560
rect 14106 6496 14122 6560
rect 14186 6496 14202 6560
rect 14266 6496 14274 6560
rect 13954 5472 14274 6496
rect 13954 5408 13962 5472
rect 14026 5408 14042 5472
rect 14106 5408 14122 5472
rect 14186 5408 14202 5472
rect 14266 5408 14274 5472
rect 13954 5090 14274 5408
rect 13954 4854 13996 5090
rect 14232 4854 14274 5090
rect 13954 4384 14274 4854
rect 13954 4320 13962 4384
rect 14026 4320 14042 4384
rect 14106 4320 14122 4384
rect 14186 4320 14202 4384
rect 14266 4320 14274 4384
rect 13954 3296 14274 4320
rect 13954 3232 13962 3296
rect 14026 3232 14042 3296
rect 14106 3232 14122 3296
rect 14186 3232 14202 3296
rect 14266 3232 14274 3296
rect 13954 2208 14274 3232
rect 13954 2144 13962 2208
rect 14026 2144 14042 2208
rect 14106 2144 14122 2208
rect 14186 2144 14202 2208
rect 14266 2144 14274 2208
rect 13954 1120 14274 2144
rect 13954 1056 13962 1120
rect 14026 1056 14042 1120
rect 14106 1056 14122 1120
rect 14186 1056 14202 1120
rect 14266 1056 14274 1120
rect 13954 32 14274 1056
rect 13954 -32 13962 32
rect 14026 -32 14042 32
rect 14106 -32 14122 32
rect 14186 -32 14202 32
rect 14266 -32 14274 32
rect 13954 -48 14274 -32
rect 15504 10368 15824 10928
rect 15504 10304 15512 10368
rect 15576 10304 15592 10368
rect 15656 10304 15672 10368
rect 15736 10304 15752 10368
rect 15816 10304 15824 10368
rect 15504 10160 15824 10304
rect 15504 9924 15546 10160
rect 15782 9924 15824 10160
rect 15504 9280 15824 9924
rect 15504 9216 15512 9280
rect 15576 9216 15592 9280
rect 15656 9216 15672 9280
rect 15736 9216 15752 9280
rect 15816 9216 15824 9280
rect 15504 8192 15824 9216
rect 15504 8128 15512 8192
rect 15576 8128 15592 8192
rect 15656 8128 15672 8192
rect 15736 8128 15752 8192
rect 15816 8128 15824 8192
rect 15504 7104 15824 8128
rect 15504 7040 15512 7104
rect 15576 7040 15592 7104
rect 15656 7040 15672 7104
rect 15736 7040 15752 7104
rect 15816 7040 15824 7104
rect 15504 6780 15824 7040
rect 15504 6544 15546 6780
rect 15782 6544 15824 6780
rect 15504 6016 15824 6544
rect 15504 5952 15512 6016
rect 15576 5952 15592 6016
rect 15656 5952 15672 6016
rect 15736 5952 15752 6016
rect 15816 5952 15824 6016
rect 15504 4928 15824 5952
rect 15504 4864 15512 4928
rect 15576 4864 15592 4928
rect 15656 4864 15672 4928
rect 15736 4864 15752 4928
rect 15816 4864 15824 4928
rect 15504 3840 15824 4864
rect 15504 3776 15512 3840
rect 15576 3776 15592 3840
rect 15656 3776 15672 3840
rect 15736 3776 15752 3840
rect 15816 3776 15824 3840
rect 15504 3400 15824 3776
rect 15504 3164 15546 3400
rect 15782 3164 15824 3400
rect 15504 2752 15824 3164
rect 15504 2688 15512 2752
rect 15576 2688 15592 2752
rect 15656 2688 15672 2752
rect 15736 2688 15752 2752
rect 15816 2688 15824 2752
rect 15504 1664 15824 2688
rect 15504 1600 15512 1664
rect 15576 1600 15592 1664
rect 15656 1600 15672 1664
rect 15736 1600 15752 1664
rect 15816 1600 15824 1664
rect 15504 576 15824 1600
rect 15504 512 15512 576
rect 15576 512 15592 576
rect 15656 512 15672 576
rect 15736 512 15752 576
rect 15816 512 15824 576
rect 15504 -48 15824 512
rect 17054 10912 17374 10928
rect 17054 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17222 10912
rect 17286 10848 17302 10912
rect 17366 10848 17374 10912
rect 17054 9824 17374 10848
rect 17054 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17222 9824
rect 17286 9760 17302 9824
rect 17366 9760 17374 9824
rect 17054 8736 17374 9760
rect 17054 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17222 8736
rect 17286 8672 17302 8736
rect 17366 8672 17374 8736
rect 17054 8470 17374 8672
rect 17054 8234 17096 8470
rect 17332 8234 17374 8470
rect 17054 7648 17374 8234
rect 17054 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17222 7648
rect 17286 7584 17302 7648
rect 17366 7584 17374 7648
rect 17054 6560 17374 7584
rect 17054 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17222 6560
rect 17286 6496 17302 6560
rect 17366 6496 17374 6560
rect 17054 5472 17374 6496
rect 17054 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17222 5472
rect 17286 5408 17302 5472
rect 17366 5408 17374 5472
rect 17054 5090 17374 5408
rect 17054 4854 17096 5090
rect 17332 4854 17374 5090
rect 17054 4384 17374 4854
rect 17054 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17222 4384
rect 17286 4320 17302 4384
rect 17366 4320 17374 4384
rect 17054 3296 17374 4320
rect 17054 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17222 3296
rect 17286 3232 17302 3296
rect 17366 3232 17374 3296
rect 17054 2208 17374 3232
rect 17054 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17222 2208
rect 17286 2144 17302 2208
rect 17366 2144 17374 2208
rect 17054 1120 17374 2144
rect 17054 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17222 1120
rect 17286 1056 17302 1120
rect 17366 1056 17374 1120
rect 17054 32 17374 1056
rect 17054 -32 17062 32
rect 17126 -32 17142 32
rect 17206 -32 17222 32
rect 17286 -32 17302 32
rect 17366 -32 17374 32
rect 17054 -48 17374 -32
<< via4 >>
rect 3146 9924 3382 10160
rect 3146 6544 3382 6780
rect 3146 3164 3382 3400
rect 4696 8234 4932 8470
rect 4696 4854 4932 5090
rect 6246 9924 6482 10160
rect 6246 6544 6482 6780
rect 6246 3164 6482 3400
rect 7796 8234 8032 8470
rect 7796 4854 8032 5090
rect 9346 9924 9582 10160
rect 9346 6544 9582 6780
rect 9346 3164 9582 3400
rect 10896 8234 11132 8470
rect 10896 4854 11132 5090
rect 12446 9924 12682 10160
rect 12446 6544 12682 6780
rect 12446 3164 12682 3400
rect 13996 8234 14232 8470
rect 13996 4854 14232 5090
rect 15546 9924 15782 10160
rect 15546 6544 15782 6780
rect 15546 3164 15782 3400
rect 17096 8234 17332 8470
rect 17096 4854 17332 5090
<< metal5 >>
rect 0 10160 18860 10202
rect 0 9924 3146 10160
rect 3382 9924 6246 10160
rect 6482 9924 9346 10160
rect 9582 9924 12446 10160
rect 12682 9924 15546 10160
rect 15782 9924 18860 10160
rect 0 9882 18860 9924
rect 0 8470 18860 8512
rect 0 8234 4696 8470
rect 4932 8234 7796 8470
rect 8032 8234 10896 8470
rect 11132 8234 13996 8470
rect 14232 8234 17096 8470
rect 17332 8234 18860 8470
rect 0 8192 18860 8234
rect 0 6780 18860 6822
rect 0 6544 3146 6780
rect 3382 6544 6246 6780
rect 6482 6544 9346 6780
rect 9582 6544 12446 6780
rect 12682 6544 15546 6780
rect 15782 6544 18860 6780
rect 0 6502 18860 6544
rect 0 5090 18860 5132
rect 0 4854 4696 5090
rect 4932 4854 7796 5090
rect 8032 4854 10896 5090
rect 11132 4854 13996 5090
rect 14232 4854 17096 5090
rect 17332 4854 18860 5090
rect 0 4812 18860 4854
rect 0 3400 18860 3442
rect 0 3164 3146 3400
rect 3382 3164 6246 3400
rect 6482 3164 9346 3400
rect 9582 3164 12446 3400
rect 12682 3164 15546 3400
rect 15782 3164 18860 3400
rect 0 3122 18860 3164
use sky130_fd_sc_hd__fill_2  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1012 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1564 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3
timestamp 1636915332
transform 1 0 276 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 276 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 0 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1636915332
transform 1 0 0 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1196 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _304_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 1564 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _473_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 368 0 -1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _410_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3312 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _359_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2944 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _303_
timestamp 1636915332
transform 1 0 2484 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1636915332
transform 1 0 2392 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1636915332
transform 1 0 2392 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_25
timestamp 1636915332
transform 1 0 2300 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp 1636915332
transform 1 0 2668 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25
timestamp 1636915332
transform 1 0 2300 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__SET_B $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 2668 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1636915332
transform 1 0 3588 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_49
timestamp 1636915332
transform 1 0 4508 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4140 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3680 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_1  _295_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 5612 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1636915332
transform 1 0 4784 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1636915332
transform 1 0 4784 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61
timestamp 1636915332
transform 1 0 5612 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__SET_B
timestamp 1636915332
transform 1 0 4600 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer10
timestamp 1636915332
transform 1 0 6808 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _421_
timestamp 1636915332
transform 1 0 6348 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1636915332
transform 1 0 5980 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66
timestamp 1636915332
transform 1 0 6072 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _476_
timestamp 1636915332
transform 1 0 4876 0 -1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__A1
timestamp 1636915332
transform 1 0 7268 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__RESET_B
timestamp 1636915332
transform -1 0 7636 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83
timestamp 1636915332
transform 1 0 7636 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_77
timestamp 1636915332
transform 1 0 7084 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1636915332
transform 1 0 7176 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1636915332
transform 1 0 8372 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1636915332
transform 1 0 7176 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _419_
timestamp 1636915332
transform 1 0 8464 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _475_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 9200 0 -1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__clkinv_2  _369_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9200 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1636915332
transform 1 0 9568 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1636915332
transform 1 0 9568 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_105
timestamp 1636915332
transform 1 0 9660 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101
timestamp 1636915332
transform 1 0 9292 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__RESET_B
timestamp 1636915332
transform 1 0 9660 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _332_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 10764 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _331_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 11224 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1636915332
transform 1 0 10764 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_122
timestamp 1636915332
transform 1 0 11224 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp 1636915332
transform 1 0 10396 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtn_1  _466_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9844 0 -1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__xor2_1  _368_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 12144 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 12328 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _309_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 12328 0 -1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1636915332
transform 1 0 11960 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1636915332
transform 1 0 11960 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_127
timestamp 1636915332
transform 1 0 11684 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131
timestamp 1636915332
transform 1 0 12052 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _367_
timestamp 1636915332
transform -1 0 13064 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _335_
timestamp 1636915332
transform -1 0 13616 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1636915332
transform 1 0 13156 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_148
timestamp 1636915332
transform 1 0 13616 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_142
timestamp 1636915332
transform 1 0 13064 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_144
timestamp 1636915332
transform 1 0 13248 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_1  _366_
timestamp 1636915332
transform 1 0 14536 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _336_
timestamp 1636915332
transform 1 0 13984 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1636915332
transform 1 0 14352 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1636915332
transform 1 0 14352 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_155
timestamp 1636915332
transform 1 0 14260 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_157
timestamp 1636915332
transform 1 0 14444 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__SET_B
timestamp 1636915332
transform 1 0 13800 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1636915332
transform 1 0 15548 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_165
timestamp 1636915332
transform 1 0 15180 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _465_
timestamp 1636915332
transform 1 0 14444 0 -1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_0_170
timestamp 1636915332
transform 1 0 15640 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _413_
timestamp 1636915332
transform 1 0 16836 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 16744 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _338_
timestamp 1636915332
transform -1 0 17112 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1636915332
transform 1 0 16744 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1636915332
transform 1 0 16744 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 18584 0 -1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _337_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 17388 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1636915332
transform 1 0 17940 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 17388 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_196
timestamp 1636915332
transform 1 0 18032 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1636915332
transform -1 0 18584 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1636915332
transform -1 0 18860 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1636915332
transform -1 0 18860 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_10
timestamp 1636915332
transform 1 0 920 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1636915332
transform 1 0 276 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1636915332
transform 1 0 0 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1636915332
transform 1 0 1196 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _300__4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 920 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtn_1  _472_
timestamp 1636915332
transform 1 0 1288 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__RESET_B
timestamp 1636915332
transform 1 0 3680 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_38
timestamp 1636915332
transform 1 0 3496 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_42
timestamp 1636915332
transform 1 0 3864 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1636915332
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _358_
timestamp 1636915332
transform 1 0 3128 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_50
timestamp 1636915332
transform 1 0 4600 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_60
timestamp 1636915332
transform 1 0 5520 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1636915332
transform 1 0 5980 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _371_
timestamp 1636915332
transform -1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _398_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4692 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _422_
timestamp 1636915332
transform 1 0 6072 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_82
timestamp 1636915332
transform 1 0 7544 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1636915332
transform 1 0 8372 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _297_
timestamp 1636915332
transform 1 0 7636 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _370_
timestamp 1636915332
transform -1 0 7544 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _420_
timestamp 1636915332
transform 1 0 8464 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_115
timestamp 1636915332
transform 1 0 10580 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1636915332
transform 1 0 10764 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10856 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _288_
timestamp 1636915332
transform -1 0 10304 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _329_
timestamp 1636915332
transform 1 0 10304 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _330_
timestamp 1636915332
transform -1 0 11500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 9936 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_2_125
timestamp 1636915332
transform 1 0 11500 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_131
timestamp 1636915332
transform 1 0 12052 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1636915332
transform 1 0 12972 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_147
timestamp 1636915332
transform 1 0 13524 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1636915332
transform 1 0 13156 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _312_
timestamp 1636915332
transform -1 0 13524 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _418_
timestamp 1636915332
transform 1 0 12144 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__RESET_B
timestamp 1636915332
transform 1 0 15916 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_151
timestamp 1636915332
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_170
timestamp 1636915332
transform 1 0 15640 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1636915332
transform 1 0 15548 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _333__6
timestamp 1636915332
transform 1 0 14260 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _334_
timestamp 1636915332
transform -1 0 14260 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _415_
timestamp 1636915332
transform 1 0 14720 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_2_196
timestamp 1636915332
transform 1 0 18032 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1636915332
transform 1 0 17940 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtn_1  _464_
timestamp 1636915332
transform 1 0 16100 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1636915332
transform -1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_12
timestamp 1636915332
transform 1 0 1104 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_20
timestamp 1636915332
transform 1 0 1840 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1636915332
transform 1 0 276 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1636915332
transform 1 0 0 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp 1636915332
transform 1 0 828 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _364_
timestamp 1636915332
transform -1 0 2392 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1636915332
transform 1 0 2392 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _301_
timestamp 1636915332
transform 1 0 2484 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _363_
timestamp 1636915332
transform 1 0 4140 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _411_
timestamp 1636915332
transform 1 0 3312 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer7
timestamp 1636915332
transform -1 0 4784 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1636915332
transform 1 0 4784 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o211ai_4  _313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4876 0 -1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__xor2_1  _372_
timestamp 1636915332
transform 1 0 6440 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A1
timestamp 1636915332
transform 1 0 7636 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_77
timestamp 1636915332
transform 1 0 7084 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_95
timestamp 1636915332
transform 1 0 8740 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_99
timestamp 1636915332
transform 1 0 9108 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1636915332
transform 1 0 7176 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _280_
timestamp 1636915332
transform -1 0 8464 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1636915332
transform -1 0 8740 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _294_
timestamp 1636915332
transform -1 0 7636 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _296_
timestamp 1636915332
transform -1 0 8188 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1636915332
transform 1 0 9568 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9660 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _287_
timestamp 1636915332
transform 1 0 9200 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10948 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 11408 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer13
timestamp 1636915332
transform -1 0 10948 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_3_131
timestamp 1636915332
transform 1 0 12052 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_137
timestamp 1636915332
transform 1 0 12604 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_147
timestamp 1636915332
transform 1 0 13524 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1636915332
transform 1 0 11960 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _417_
timestamp 1636915332
transform 1 0 12696 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_3_166
timestamp 1636915332
transform 1 0 15272 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_172
timestamp 1636915332
transform 1 0 15824 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1636915332
transform 1 0 14352 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _328_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 13800 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _414_
timestamp 1636915332
transform -1 0 16744 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _416_
timestamp 1636915332
transform 1 0 14444 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1636915332
transform 1 0 16744 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _438_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 16836 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_3_199
timestamp 1636915332
transform 1 0 18308 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1636915332
transform -1 0 18860 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_11
timestamp 1636915332
transform 1 0 1012 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_14
timestamp 1636915332
transform 1 0 1288 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1636915332
transform 1 0 276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1636915332
transform 1 0 644 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1636915332
transform 1 0 0 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1636915332
transform 1 0 1196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _299_
timestamp 1636915332
transform 1 0 736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _365_
timestamp 1636915332
transform 1 0 1840 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_4_34
timestamp 1636915332
transform 1 0 3128 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_47
timestamp 1636915332
transform 1 0 4324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1636915332
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 5244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _360_
timestamp 1636915332
transform 1 0 2484 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _361_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 3588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer12
timestamp 1636915332
transform -1 0 4324 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_4_57
timestamp 1636915332
transform 1 0 5244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1636915332
transform 1 0 5980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _293_
timestamp 1636915332
transform -1 0 6808 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _423_
timestamp 1636915332
transform 1 0 6808 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer6
timestamp 1636915332
transform -1 0 5980 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_4_83
timestamp 1636915332
transform 1 0 7636 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_92
timestamp 1636915332
transform 1 0 8464 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1636915332
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  _352_
timestamp 1636915332
transform 1 0 8556 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_4_100
timestamp 1636915332
transform 1 0 9200 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_107
timestamp 1636915332
transform 1 0 9844 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_115
timestamp 1636915332
transform 1 0 10580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_118
timestamp 1636915332
transform 1 0 10856 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1636915332
transform 1 0 10764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _310_
timestamp 1636915332
transform -1 0 11408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _315_
timestamp 1636915332
transform -1 0 11776 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer9
timestamp 1636915332
transform 1 0 9568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__RESET_B
timestamp 1636915332
transform 1 0 13248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_131
timestamp 1636915332
transform 1 0 12052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1636915332
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1636915332
transform -1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _467_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 13432 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1636915332
transform 1 0 15548 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _439_
timestamp 1636915332
transform 1 0 15640 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1636915332
transform 1 0 17940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _322_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 17112 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _324_
timestamp 1636915332
transform -1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1636915332
transform 1 0 17664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A
timestamp 1636915332
transform -1 0 18584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1636915332
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__RESET_B
timestamp 1636915332
transform 1 0 2116 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1636915332
transform 1 0 0 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _474_
timestamp 1636915332
transform 1 0 276 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_5_25
timestamp 1636915332
transform 1 0 2300 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1636915332
transform 1 0 2392 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _298_
timestamp 1636915332
transform 1 0 2484 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _362_
timestamp 1636915332
transform 1 0 4140 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1636915332
transform 1 0 3312 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_51
timestamp 1636915332
transform 1 0 4692 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1636915332
transform 1 0 4784 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _477_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5152 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer5
timestamp 1636915332
transform -1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_76
timestamp 1636915332
transform 1 0 6992 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_83
timestamp 1636915332
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_99
timestamp 1636915332
transform 1 0 9108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1636915332
transform 1 0 7176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 9108 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _289_
timestamp 1636915332
transform -1 0 8556 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _292_
timestamp 1636915332
transform -1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_103
timestamp 1636915332
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_108
timestamp 1636915332
transform 1 0 9936 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_120
timestamp 1636915332
transform 1 0 11040 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1636915332
transform 1 0 9568 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1636915332
transform -1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__SET_B
timestamp 1636915332
transform 1 0 11776 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1636915332
transform 1 0 11960 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _471_
timestamp 1636915332
transform 1 0 12052 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1636915332
transform 1 0 14352 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _326_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 14904 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _327_
timestamp 1636915332
transform 1 0 13984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _451_
timestamp 1636915332
transform 1 0 14904 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__B_N
timestamp 1636915332
transform 1 0 17572 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__D
timestamp 1636915332
transform 1 0 17756 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__RESET_B
timestamp 1636915332
transform 1 0 16836 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1636915332
transform -1 0 18124 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1636915332
transform 1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1636915332
transform 1 0 16744 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _323_
timestamp 1636915332
transform 1 0 17020 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_201
timestamp 1636915332
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1636915332
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1636915332
transform 1 0 1012 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_17
timestamp 1636915332
transform 1 0 1564 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1636915332
transform 1 0 276 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1636915332
transform 1 0 276 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1636915332
transform 1 0 0 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1636915332
transform 1 0 0 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1636915332
transform 1 0 1196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _321_
timestamp 1636915332
transform 1 0 1288 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_2  _468_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 460 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _318_
timestamp 1636915332
transform 1 0 2576 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _306_
timestamp 1636915332
transform -1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1636915332
transform 1 0 2392 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_27
timestamp 1636915332
transform 1 0 2484 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_28
timestamp 1636915332
transform 1 0 2576 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_25
timestamp 1636915332
transform 1 0 2300 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__SET_B
timestamp 1636915332
transform 1 0 2392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _425_
timestamp 1636915332
transform 1 0 3680 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _320_
timestamp 1636915332
transform 1 0 3404 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1636915332
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp 1636915332
transform 1 0 3404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_2  _373_
timestamp 1636915332
transform -1 0 4600 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__A1
timestamp 1636915332
transform 1 0 4508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer16
timestamp 1636915332
transform 1 0 5244 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer11
timestamp 1636915332
transform 1 0 4692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1636915332
transform 1 0 4784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_53
timestamp 1636915332
transform 1 0 4876 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_50
timestamp 1636915332
transform 1 0 4600 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_56
timestamp 1636915332
transform 1 0 5152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__477__RESET_B
timestamp 1636915332
transform 1 0 4968 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _424_
timestamp 1636915332
transform 1 0 6348 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _316_
timestamp 1636915332
transform 1 0 5612 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1636915332
transform 1 0 5980 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_67
timestamp 1636915332
transform 1 0 6164 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_66
timestamp 1636915332
transform 1 0 6072 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_64
timestamp 1636915332
transform 1 0 5888 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__RESET_B
timestamp 1636915332
transform 1 0 5980 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _340_
timestamp 1636915332
transform 1 0 7268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1636915332
transform 1 0 7176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_82
timestamp 1636915332
transform 1 0 7544 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_75
timestamp 1636915332
transform 1 0 6900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_84
timestamp 1636915332
transform 1 0 7728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_78
timestamp 1636915332
transform 1 0 7176 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__SET_B
timestamp 1636915332
transform 1 0 7820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_4  _341_
timestamp 1636915332
transform -1 0 9016 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _290_
timestamp 1636915332
transform 1 0 8004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1636915332
transform 1 0 8372 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_98
timestamp 1636915332
transform 1 0 9016 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_90
timestamp 1636915332
transform 1 0 8280 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _478_
timestamp 1636915332
transform 1 0 8464 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_6_113
timestamp 1636915332
transform 1 0 10396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_105
timestamp 1636915332
transform 1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1636915332
transform 1 0 9568 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1636915332
transform 1 0 10764 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _354_
timestamp 1636915332
transform 1 0 10856 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2ai_2  _355_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_4  _305__5
timestamp 1636915332
transform -1 0 12604 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1636915332
transform 1 0 11960 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_131
timestamp 1636915332
transform 1 0 12052 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_129
timestamp 1636915332
transform 1 0 11868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_125
timestamp 1636915332
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_131
timestamp 1636915332
transform 1 0 12052 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_125
timestamp 1636915332
transform 1 0 11500 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__RESET_B
timestamp 1636915332
transform 1 0 12236 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _325_
timestamp 1636915332
transform -1 0 13156 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1636915332
transform 1 0 13156 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp 1636915332
transform 1 0 12604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _453_
timestamp 1636915332
transform -1 0 14260 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _440_
timestamp 1636915332
transform 1 0 13248 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  split8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 14444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _283_
timestamp 1636915332
transform -1 0 15272 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1636915332
transform 1 0 14352 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_155
timestamp 1636915332
transform 1 0 14260 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1636915332
transform 1 0 15548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_168
timestamp 1636915332
transform 1 0 15456 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__RESET_B
timestamp 1636915332
transform 1 0 15640 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__A2
timestamp 1636915332
transform 1 0 15272 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _454_
timestamp 1636915332
transform 1 0 15824 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _452_
timestamp 1636915332
transform 1 0 14812 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__SET_B
timestamp 1636915332
transform 1 0 16836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__SET_B
timestamp 1636915332
transform 1 0 17020 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1636915332
transform -1 0 18308 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_196
timestamp 1636915332
transform 1 0 18032 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_187
timestamp 1636915332
transform 1 0 17204 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1636915332
transform 1 0 16744 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1636915332
transform 1 0 17940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  _392_
timestamp 1636915332
transform 1 0 17756 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_7_200
timestamp 1636915332
transform 1 0 18400 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1636915332
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1636915332
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1636915332
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_12
timestamp 1636915332
transform 1 0 1104 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1636915332
transform 1 0 276 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1636915332
transform 1 0 0 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1636915332
transform 1 0 1196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _319_
timestamp 1636915332
transform -1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _469_
timestamp 1636915332
transform 1 0 1288 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__RESET_B
timestamp 1636915332
transform 1 0 3220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_37
timestamp 1636915332
transform 1 0 3404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1636915332
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_1  _351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4508 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _426_
timestamp 1636915332
transform 1 0 3680 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_55
timestamp 1636915332
transform 1 0 5060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1636915332
transform 1 0 5980 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _317_
timestamp 1636915332
transform 1 0 5336 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _470_
timestamp 1636915332
transform 1 0 6072 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__463__SET_B
timestamp 1636915332
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_90
timestamp 1636915332
transform 1 0 8280 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_92
timestamp 1636915332
transform 1 0 8464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1636915332
transform 1 0 8372 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _342_
timestamp 1636915332
transform 1 0 7912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _463_
timestamp 1636915332
transform 1 0 8832 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1636915332
transform 1 0 10764 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _435_
timestamp 1636915332
transform 1 0 10856 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__RESET_B
timestamp 1636915332
transform 1 0 11868 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__456__RESET_B
timestamp 1636915332
transform 1 0 13248 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_127
timestamp 1636915332
transform 1 0 11684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_131
timestamp 1636915332
transform 1 0 12052 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1636915332
transform 1 0 13156 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _456_
timestamp 1636915332
transform 1 0 13432 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_8_170
timestamp 1636915332
transform 1 0 15640 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1636915332
transform 1 0 15548 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _455_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 15732 0 1 4352
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1636915332
transform 1 0 17940 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  split4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 18032 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1636915332
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_14
timestamp 1636915332
transform 1 0 1288 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_18
timestamp 1636915332
transform 1 0 1656 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1636915332
transform 1 0 276 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1636915332
transform 1 0 0 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp 1636915332
transform -1 0 1288 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _377_
timestamp 1636915332
transform 1 0 1748 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_9_43
timestamp 1636915332
transform 1 0 3956 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1636915332
transform 1 0 2392 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _248_
timestamp 1636915332
transform 1 0 2484 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _251_
timestamp 1636915332
transform 1 0 4508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _374_
timestamp 1636915332
transform 1 0 3312 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1636915332
transform 1 0 5704 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_68
timestamp 1636915332
transform 1 0 6256 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_72
timestamp 1636915332
transform 1 0 6624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1636915332
transform 1 0 4784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _250_
timestamp 1636915332
transform 1 0 4876 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  _375_
timestamp 1636915332
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_pll_clk
timestamp 1636915332
transform -1 0 7084 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_77
timestamp 1636915332
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_79
timestamp 1636915332
transform 1 0 7268 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_87
timestamp 1636915332
transform 1 0 8004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_97
timestamp 1636915332
transform 1 0 8924 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1636915332
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _222_
timestamp 1636915332
transform -1 0 9476 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _343_
timestamp 1636915332
transform 1 0 8280 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_9_103
timestamp 1636915332
transform 1 0 9476 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1636915332
transform 1 0 9568 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _441_
timestamp 1636915332
transform -1 0 11132 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_pll_clk
timestamp 1636915332
transform 1 0 11132 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__B
timestamp 1636915332
transform 1 0 11776 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1636915332
transform 1 0 11960 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _349_
timestamp 1636915332
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _448_
timestamp 1636915332
transform -1 0 13892 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__SET_B
timestamp 1636915332
transform 1 0 14168 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_151
timestamp 1636915332
transform 1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1636915332
transform 1 0 14352 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _492_
timestamp 1636915332
transform 1 0 14444 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_9_190
timestamp 1636915332
transform 1 0 17480 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1636915332
transform 1 0 16744 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _395_
timestamp 1636915332
transform -1 0 17480 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  split15
timestamp 1636915332
transform -1 0 16744 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1636915332
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1636915332
transform 1 0 276 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1636915332
transform 1 0 644 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1636915332
transform 1 0 0 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1636915332
transform 1 0 1196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _247__1
timestamp 1636915332
transform 1 0 736 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dfstp_1  _485_
timestamp 1636915332
transform 1 0 1288 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__RESET_B
timestamp 1636915332
transform 1 0 3956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__SET_B
timestamp 1636915332
transform 1 0 3220 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_37
timestamp 1636915332
transform 1 0 3404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_40
timestamp 1636915332
transform 1 0 3680 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1636915332
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtn_1  _484_
timestamp 1636915332
transform 1 0 4140 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_10_73
timestamp 1636915332
transform 1 0 6716 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1636915332
transform 1 0 5980 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _376_
timestamp 1636915332
transform 1 0 6072 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_10_92
timestamp 1636915332
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1636915332
transform 1 0 8372 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _442_
timestamp 1636915332
transform 1 0 6900 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 10488 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__RESET_B
timestamp 1636915332
transform 1 0 10948 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk_A
timestamp 1636915332
transform 1 0 10488 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_116
timestamp 1636915332
transform 1 0 10672 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_118
timestamp 1636915332
transform 1 0 10856 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1636915332
transform 1 0 10764 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _493_
timestamp 1636915332
transform 1 0 11132 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1636915332
transform 1 0 12972 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1636915332
transform 1 0 13156 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _391_
timestamp 1636915332
transform 1 0 13248 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__RESET_B
timestamp 1636915332
transform 1 0 15364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__RESET_B
timestamp 1636915332
transform 1 0 13984 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_151
timestamp 1636915332
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_166
timestamp 1636915332
transform 1 0 15272 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_170
timestamp 1636915332
transform 1 0 15640 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1636915332
transform 1 0 15548 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _218_
timestamp 1636915332
transform -1 0 14996 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 1636915332
transform 1 0 14996 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _394_
timestamp 1636915332
transform -1 0 16100 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1636915332
transform -1 0 18308 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_196
timestamp 1636915332
transform 1 0 18032 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1636915332
transform 1 0 17940 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _457_
timestamp 1636915332
transform -1 0 17940 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1636915332
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1636915332
transform 1 0 18308 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__RESET_B
timestamp 1636915332
transform 1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1636915332
transform 1 0 0 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _486_
timestamp 1636915332
transform 1 0 276 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_11_25
timestamp 1636915332
transform 1 0 2300 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_30
timestamp 1636915332
transform 1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_42
timestamp 1636915332
transform 1 0 3864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_49
timestamp 1636915332
transform 1 0 4508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1636915332
transform 1 0 2392 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _379_
timestamp 1636915332
transform 1 0 3956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _381_
timestamp 1636915332
transform -1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _428_
timestamp 1636915332
transform 1 0 3036 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_53
timestamp 1636915332
transform 1 0 4876 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1636915332
transform 1 0 4784 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _397_
timestamp 1636915332
transform 1 0 5244 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _427_
timestamp 1636915332
transform 1 0 6072 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__RESET_B
timestamp 1636915332
transform 1 0 9108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_75
timestamp 1636915332
transform 1 0 6900 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_79
timestamp 1636915332
transform 1 0 7268 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1636915332
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _220_
timestamp 1636915332
transform 1 0 8556 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _221_
timestamp 1636915332
transform 1 0 8004 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _230_
timestamp 1636915332
transform 1 0 7452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_101
timestamp 1636915332
transform 1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_105
timestamp 1636915332
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_117
timestamp 1636915332
transform 1 0 10764 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1636915332
transform 1 0 9568 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_125
timestamp 1636915332
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_131
timestamp 1636915332
transform 1 0 12052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_143
timestamp 1636915332
transform 1 0 13156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1636915332
transform 1 0 11960 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _216_
timestamp 1636915332
transform 1 0 12328 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1636915332
transform 1 0 11684 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _434_
timestamp 1636915332
transform 1 0 13432 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_155
timestamp 1636915332
transform 1 0 14260 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_157
timestamp 1636915332
transform 1 0 14444 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1636915332
transform 1 0 14352 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _390_
timestamp 1636915332
transform 1 0 14536 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp 1636915332
transform 1 0 14904 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_11_193
timestamp 1636915332
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1636915332
transform 1 0 16744 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_2  _274_
timestamp 1636915332
transform 1 0 16836 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_11_201
timestamp 1636915332
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1636915332
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1636915332
transform 1 0 1012 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_14
timestamp 1636915332
transform 1 0 1288 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1636915332
transform 1 0 276 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1636915332
transform 1 0 644 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1636915332
transform 1 0 0 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1636915332
transform 1 0 1196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _245_
timestamp 1636915332
transform 1 0 1564 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1636915332
transform 1 0 736 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_38
timestamp 1636915332
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_40
timestamp 1636915332
transform 1 0 3680 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1636915332
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _253_
timestamp 1636915332
transform -1 0 2668 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_4  _260_
timestamp 1636915332
transform -1 0 5428 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _429_
timestamp 1636915332
transform 1 0 2668 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__RESET_B
timestamp 1636915332
transform 1 0 5796 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_59
timestamp 1636915332
transform 1 0 5428 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1636915332
transform 1 0 5980 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _243_
timestamp 1636915332
transform 1 0 6072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _487_
timestamp 1636915332
transform -1 0 8372 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_12_92
timestamp 1636915332
transform 1 0 8464 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1636915332
transform 1 0 8372 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _491_
timestamp 1636915332
transform 1 0 8556 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_12_116
timestamp 1636915332
transform 1 0 10672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1636915332
transform 1 0 10764 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _443_
timestamp 1636915332
transform 1 0 10856 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_139
timestamp 1636915332
transform 1 0 12788 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_144
timestamp 1636915332
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1636915332
transform 1 0 13156 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _224_
timestamp 1636915332
transform -1 0 12788 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__RESET_B
timestamp 1636915332
transform 1 0 15640 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__SET_B
timestamp 1636915332
transform 1 0 14444 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1636915332
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_159
timestamp 1636915332
transform 1 0 14628 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1636915332
transform 1 0 15548 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _278_
timestamp 1636915332
transform -1 0 14444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _409_
timestamp 1636915332
transform 1 0 14720 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _460_
timestamp 1636915332
transform -1 0 17940 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1636915332
transform -1 0 18308 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_196
timestamp 1636915332
transform 1 0 18032 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1636915332
transform 1 0 17940 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1636915332
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1636915332
transform 1 0 18308 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1636915332
transform 1 0 0 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1636915332
transform 1 0 0 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1636915332
transform 1 0 276 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1636915332
transform 1 0 1012 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1636915332
transform -1 0 2484 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _273_
timestamp 1636915332
transform -1 0 1656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _272_
timestamp 1636915332
transform -1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1636915332
transform -1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1636915332
transform 1 0 1196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_19
timestamp 1636915332
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_15
timestamp 1636915332
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1636915332
transform 1 0 276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _401_
timestamp 1636915332
transform 1 0 2484 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _382_
timestamp 1636915332
transform 1 0 2484 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1636915332
transform 1 0 2392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_36
timestamp 1636915332
transform 1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_34
timestamp 1636915332
transform 1 0 3128 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _380_
timestamp 1636915332
transform 1 0 4232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _378_
timestamp 1636915332
transform -1 0 4232 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1636915332
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_49
timestamp 1636915332
transform 1 0 4508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_40
timestamp 1636915332
transform 1 0 3680 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__o211a_1  _254_
timestamp 1636915332
transform -1 0 5612 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_4  _228_
timestamp 1636915332
transform 1 0 5336 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1636915332
transform 1 0 4784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_52
timestamp 1636915332
transform 1 0 4784 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_61
timestamp 1636915332
transform 1 0 5612 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_1  _244_
timestamp 1636915332
transform 1 0 6440 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _229_
timestamp 1636915332
transform -1 0 6256 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1636915332
transform 1 0 5980 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_68
timestamp 1636915332
transform 1 0 6256 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__488__SET_B
timestamp 1636915332
transform 1 0 6072 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_1  _488_
timestamp 1636915332
transform 1 0 6256 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_14_89
timestamp 1636915332
transform 1 0 8188 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_92
timestamp 1636915332
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1636915332
transform 1 0 7176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1636915332
transform 1 0 8372 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _236_
timestamp 1636915332
transform 1 0 7268 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1636915332
transform 1 0 8464 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _433_
timestamp 1636915332
transform 1 0 7636 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk90
timestamp 1636915332
transform -1 0 10672 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_13_101
timestamp 1636915332
transform 1 0 9292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_105
timestamp 1636915332
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_116
timestamp 1636915332
transform 1 0 10672 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1636915332
transform 1 0 9568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1636915332
transform 1 0 10764 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _386_
timestamp 1636915332
transform -1 0 11224 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _405_
timestamp 1636915332
transform 1 0 10856 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _432_
timestamp 1636915332
transform 1 0 10028 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_pll_clk90
timestamp 1636915332
transform 1 0 11224 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _232_
timestamp 1636915332
transform 1 0 11684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _226_
timestamp 1636915332
transform -1 0 12420 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1636915332
transform 1 0 11960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_132
timestamp 1636915332
transform 1 0 12144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_126
timestamp 1636915332
transform 1 0 11592 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk90_A
timestamp 1636915332
transform 1 0 11960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_1  _225_
timestamp 1636915332
transform 1 0 12512 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _223_
timestamp 1636915332
transform 1 0 12420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_138
timestamp 1636915332
transform 1 0 12696 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _279_
timestamp 1636915332
transform 1 0 13524 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1636915332
transform 1 0 13156 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_146
timestamp 1636915332
transform 1 0 13432 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_142
timestamp 1636915332
transform 1 0 13064 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_146
timestamp 1636915332
transform 1 0 13432 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__SET_B
timestamp 1636915332
transform 1 0 13248 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_170
timestamp 1636915332
transform 1 0 15640 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1636915332
transform 1 0 14352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1636915332
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  _275_
timestamp 1636915332
transform -1 0 14444 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 13800 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2ai_2  _357_
timestamp 1636915332
transform -1 0 15548 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dfstp_4  _461_
timestamp 1636915332
transform -1 0 17940 0 1 7616
box -38 -48 2246 592
use sky130_fd_sc_hd__dfstp_1  _479_
timestamp 1636915332
transform 1 0 14444 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__SET_B
timestamp 1636915332
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_180
timestamp 1636915332
transform 1 0 16560 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_190
timestamp 1636915332
transform 1 0 17480 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_196
timestamp 1636915332
transform 1 0 18032 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1636915332
transform 1 0 16744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1636915332
transform 1 0 17940 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  _276_
timestamp 1636915332
transform 1 0 16836 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1636915332
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1636915332
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1636915332
transform 1 0 0 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _264_
timestamp 1636915332
transform -1 0 2392 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _480_
timestamp 1636915332
transform 1 0 276 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1636915332
transform 1 0 2392 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _383_
timestamp 1636915332
transform 1 0 2484 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _403_
timestamp 1636915332
transform 1 0 3956 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp 1636915332
transform 1 0 3128 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1636915332
transform 1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_59
timestamp 1636915332
transform 1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_70
timestamp 1636915332
transform 1 0 6440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1636915332
transform 1 0 4784 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _227_
timestamp 1636915332
transform 1 0 5704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _235_
timestamp 1636915332
transform -1 0 6440 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _263_
timestamp 1636915332
transform -1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _389_
timestamp 1636915332
transform 1 0 6532 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_15_79
timestamp 1636915332
transform 1 0 7268 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1636915332
transform 1 0 7176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _387_
timestamp 1636915332
transform 1 0 8924 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _444_
timestamp 1636915332
transform 1 0 7452 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1636915332
transform 1 0 10396 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1636915332
transform 1 0 9568 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  _353_
timestamp 1636915332
transform -1 0 11960 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _436_
timestamp 1636915332
transform -1 0 11316 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__SET_B
timestamp 1636915332
transform 1 0 13524 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_146
timestamp 1636915332
transform 1 0 13432 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1636915332
transform 1 0 11960 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _231_
timestamp 1636915332
transform 1 0 12052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _234_
timestamp 1636915332
transform 1 0 12328 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _237_
timestamp 1636915332
transform -1 0 13432 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _356_
timestamp 1636915332
transform 1 0 13708 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_15_160
timestamp 1636915332
transform 1 0 14720 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1636915332
transform 1 0 14352 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1636915332
transform -1 0 14720 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _458_
timestamp 1636915332
transform 1 0 14812 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1636915332
transform -1 0 18308 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_192
timestamp 1636915332
transform 1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_196
timestamp 1636915332
transform 1 0 18032 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1636915332
transform 1 0 16744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _437_
timestamp 1636915332
transform 1 0 16836 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1636915332
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1636915332
transform 1 0 18308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1636915332
transform -1 0 1472 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1636915332
transform 1 0 276 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_9
timestamp 1636915332
transform 1 0 828 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1636915332
transform 1 0 0 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1636915332
transform 1 0 1196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _268_
timestamp 1636915332
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1472 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__RESET_B
timestamp 1636915332
transform 1 0 2944 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_34
timestamp 1636915332
transform 1 0 3128 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_38
timestamp 1636915332
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_40
timestamp 1636915332
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1636915332
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _431_
timestamp 1636915332
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_50
timestamp 1636915332
transform 1 0 4600 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_62
timestamp 1636915332
transform 1 0 5704 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_66
timestamp 1636915332
transform 1 0 6072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1636915332
transform 1 0 5980 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _241_
timestamp 1636915332
transform -1 0 7176 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _257_
timestamp 1636915332
transform 1 0 5336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_pll_clk90
timestamp 1636915332
transform -1 0 6808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_78
timestamp 1636915332
transform 1 0 7176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_88
timestamp 1636915332
transform 1 0 8096 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1636915332
transform 1 0 8372 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _240_
timestamp 1636915332
transform -1 0 9200 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _242_
timestamp 1636915332
transform 1 0 7360 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_104
timestamp 1636915332
transform 1 0 9568 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1636915332
transform 1 0 10764 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _239_
timestamp 1636915332
transform -1 0 9568 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _388_
timestamp 1636915332
transform 1 0 10488 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _407_
timestamp 1636915332
transform 1 0 10856 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1636915332
transform 1 0 9660 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_127
timestamp 1636915332
transform 1 0 11684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_142
timestamp 1636915332
transform 1 0 13064 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1636915332
transform 1 0 13156 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _238_
timestamp 1636915332
transform -1 0 13064 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1636915332
transform 1 0 11868 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _490_
timestamp 1636915332
transform 1 0 13248 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__462__RESET_B
timestamp 1636915332
transform 1 0 15640 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_165
timestamp 1636915332
transform 1 0 15180 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1636915332
transform 1 0 15548 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _350_
timestamp 1636915332
transform -1 0 15548 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _462_
timestamp 1636915332
transform -1 0 17940 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_6  FILLER_16_196
timestamp 1636915332
transform 1 0 18032 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1636915332
transform 1 0 17940 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1636915332
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__481__SET_B
timestamp 1636915332
transform 1 0 2208 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1636915332
transform 1 0 0 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _481_
timestamp 1636915332
transform 1 0 276 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_17_47
timestamp 1636915332
transform 1 0 4324 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1636915332
transform 1 0 2392 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_2  _256_
timestamp 1636915332
transform -1 0 3772 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _258_
timestamp 1636915332
transform 1 0 3772 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _259_
timestamp 1636915332
transform 1 0 4048 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _265_
timestamp 1636915332
transform -1 0 2852 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_51
timestamp 1636915332
transform 1 0 4692 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1636915332
transform 1 0 4784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1636915332
transform -1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _261_
timestamp 1636915332
transform -1 0 6256 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _262_
timestamp 1636915332
transform -1 0 6624 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _430_
timestamp 1636915332
transform 1 0 4876 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__489__RESET_B
timestamp 1636915332
transform 1 0 7360 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_75
timestamp 1636915332
transform 1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_79
timestamp 1636915332
transform 1 0 7268 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1636915332
transform 1 0 7176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 1636915332
transform 1 0 7544 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_ext_clk_A
timestamp 1636915332
transform -1 0 9936 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_102
timestamp 1636915332
transform 1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_105
timestamp 1636915332
transform 1 0 9660 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1636915332
transform 1 0 9568 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ext_clk
timestamp 1636915332
transform 1 0 9936 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__459__RESET_B
timestamp 1636915332
transform 1 0 11776 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_135
timestamp 1636915332
transform 1 0 12420 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1636915332
transform 1 0 11960 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _459_
timestamp 1636915332
transform 1 0 12512 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_ext_clk
timestamp 1636915332
transform -1 0 12420 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__SET_B
timestamp 1636915332
transform 1 0 14536 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_157
timestamp 1636915332
transform 1 0 14444 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1636915332
transform 1 0 14352 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _446_
timestamp 1636915332
transform 1 0 14720 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_17_181
timestamp 1636915332
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_191
timestamp 1636915332
transform 1 0 17572 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1636915332
transform 1 0 16744 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1636915332
transform 1 0 16836 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_199
timestamp 1636915332
transform 1 0 18308 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1636915332
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1636915332
transform 1 0 276 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1636915332
transform 1 0 828 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1636915332
transform 1 0 0 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1636915332
transform 1 0 1196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _267__3
timestamp 1636915332
transform -1 0 828 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _269_
timestamp 1636915332
transform -1 0 1656 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _270_
timestamp 1636915332
transform -1 0 1196 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _482_
timestamp 1636915332
transform 1 0 1656 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__RESET_B
timestamp 1636915332
transform 1 0 3956 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_38
timestamp 1636915332
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_45
timestamp 1636915332
transform 1 0 4140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1636915332
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _384_
timestamp 1636915332
transform -1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__SET_B
timestamp 1636915332
transform 1 0 5796 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_57
timestamp 1636915332
transform 1 0 5244 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1636915332
transform 1 0 5980 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _483_
timestamp 1636915332
transform 1 0 6072 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__S
timestamp 1636915332
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__RESET_B
timestamp 1636915332
transform 1 0 8740 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1636915332
transform 1 0 8004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_94
timestamp 1636915332
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1636915332
transform 1 0 8372 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _450_
timestamp 1636915332
transform 1 0 8924 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1636915332
transform 1 0 10764 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _449_
timestamp 1636915332
transform 1 0 10856 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__SET_B
timestamp 1636915332
transform 1 0 12972 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_138
timestamp 1636915332
transform 1 0 12696 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1636915332
transform 1 0 13156 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _447_
timestamp 1636915332
transform 1 0 13248 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__SET_B
timestamp 1636915332
transform 1 0 15824 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_165
timestamp 1636915332
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_170
timestamp 1636915332
transform 1 0 15640 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1636915332
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1636915332
transform -1 0 18308 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_196
timestamp 1636915332
transform 1 0 18032 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1636915332
transform 1 0 17940 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _445_
timestamp 1636915332
transform 1 0 16008 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1636915332
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1636915332
transform 1 0 18308 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1636915332
transform 1 0 1012 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_14
timestamp 1636915332
transform 1 0 1288 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_20
timestamp 1636915332
transform 1 0 1840 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_24
timestamp 1636915332
transform 1 0 2208 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1636915332
transform 1 0 276 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1636915332
transform 1 0 0 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1636915332
transform 1 0 1196 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _266_
timestamp 1636915332
transform -1 0 2208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1636915332
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_47
timestamp 1636915332
transform 1 0 4324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1636915332
transform 1 0 2392 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1636915332
transform 1 0 3588 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _385_
timestamp 1636915332
transform 1 0 3680 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_19_51
timestamp 1636915332
transform 1 0 4692 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_53
timestamp 1636915332
transform 1 0 4876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_66
timestamp 1636915332
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_72
timestamp 1636915332
transform 1 0 6624 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1636915332
transform 1 0 4784 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1636915332
transform 1 0 5980 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _252__2
timestamp 1636915332
transform -1 0 6624 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_19_82
timestamp 1636915332
transform 1 0 7544 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1636915332
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1636915332
transform 1 0 8372 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _347_
timestamp 1636915332
transform 1 0 8464 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _348_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8004 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_ext_clk
timestamp 1636915332
transform 1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output10
timestamp 1636915332
transform 1 0 7268 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__RESET_B
timestamp 1636915332
transform 1 0 10856 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_101
timestamp 1636915332
transform 1 0 9292 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_105
timestamp 1636915332
transform 1 0 9660 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_112
timestamp 1636915332
transform 1 0 10304 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_116
timestamp 1636915332
transform 1 0 10672 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_120
timestamp 1636915332
transform 1 0 11040 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1636915332
transform 1 0 9568 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1636915332
transform 1 0 10764 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  output12
timestamp 1636915332
transform 1 0 10028 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1636915332
transform 1 0 11776 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_140
timestamp 1636915332
transform 1 0 12880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_144
timestamp 1636915332
transform 1 0 13248 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1636915332
transform 1 0 11960 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1636915332
transform 1 0 13156 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _344__9
timestamp 1636915332
transform -1 0 13800 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _399_
timestamp 1636915332
transform -1 0 12880 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_154
timestamp 1636915332
transform 1 0 14168 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_160
timestamp 1636915332
transform 1 0 14720 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_166
timestamp 1636915332
transform 1 0 15272 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1636915332
transform 1 0 14352 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1636915332
transform 1 0 15548 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _345__8
timestamp 1636915332
transform -1 0 15272 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  _396__13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 14720 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1636915332
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1636915332
transform -1 0 14168 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1636915332
transform -1 0 17940 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1636915332
transform 1 0 16376 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_188
timestamp 1636915332
transform 1 0 17296 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_192
timestamp 1636915332
transform 1 0 17664 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1636915332
transform 1 0 16744 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1636915332
transform 1 0 17940 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _346__7
timestamp 1636915332
transform -1 0 17296 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _393_
timestamp 1636915332
transform 1 0 18032 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1636915332
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1636915332
transform 1 0 18308 0 -1 10880
box -38 -48 314 592
<< labels >>
rlabel metal5 s 0 4812 18860 5132 6 VGND
port 0 nsew ground input
rlabel metal5 s 0 8192 18860 8512 6 VGND
port 0 nsew ground input
rlabel metal4 s 4654 -48 4974 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 7754 -48 8074 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 10854 -48 11174 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 13954 -48 14274 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 17054 -48 17374 10928 6 VGND
port 0 nsew ground input
rlabel metal5 s 0 3122 18860 3442 6 VPWR
port 1 nsew power input
rlabel metal5 s 0 6502 18860 6822 6 VPWR
port 1 nsew power input
rlabel metal5 s 0 9882 18860 10202 6 VPWR
port 1 nsew power input
rlabel metal4 s 3104 -48 3424 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 6204 -48 6524 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 9304 -48 9624 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 12404 -48 12724 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 15504 -48 15824 10928 6 VPWR
port 1 nsew power input
rlabel metal2 s 7102 11200 7158 12000 6 core_clk
port 2 nsew signal tristate
rlabel metal2 s 4250 11200 4306 12000 6 ext_clk
port 3 nsew signal input
rlabel metal3 s 19200 688 20000 808 6 ext_clk_sel
port 4 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 ext_reset
port 5 nsew signal input
rlabel metal2 s 15658 11200 15714 12000 6 pll_clk
port 6 nsew signal input
rlabel metal2 s 18510 11200 18566 12000 6 pll_clk90
port 7 nsew signal input
rlabel metal2 s 1398 11200 1454 12000 6 resetb
port 8 nsew signal input
rlabel metal2 s 12806 11200 12862 12000 6 resetb_sync
port 9 nsew signal tristate
rlabel metal3 s 19200 6672 20000 6792 6 sel2[0]
port 10 nsew signal input
rlabel metal3 s 19200 8168 20000 8288 6 sel2[1]
port 11 nsew signal input
rlabel metal3 s 19200 9664 20000 9784 6 sel2[2]
port 12 nsew signal input
rlabel metal3 s 19200 2184 20000 2304 6 sel[0]
port 13 nsew signal input
rlabel metal3 s 19200 3680 20000 3800 6 sel[1]
port 14 nsew signal input
rlabel metal3 s 19200 5176 20000 5296 6 sel[2]
port 15 nsew signal input
rlabel metal2 s 9954 11200 10010 12000 6 user_clk
port 16 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 12000
<< end >>
