module empty_macro ();
endmodule
