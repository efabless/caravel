* NGSPICE file created from mgmt_protect.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for mprj2_logic_high abstract view
.subckt mprj2_logic_high HI vccd2 vssd2
.ends

* Black-box entry subcircuit for mprj_logic_high abstract view
.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[287] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295]
+ HI[296] HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304]
+ HI[305] HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314]
+ HI[315] HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334]
+ HI[335] HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344]
+ HI[345] HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354]
+ HI[355] HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374]
+ HI[375] HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384]
+ HI[385] HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394]
+ HI[395] HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403]
+ HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413]
+ HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423]
+ HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[42] HI[430] HI[431] HI[432] HI[433]
+ HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443]
+ HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453]
+ HI[454] HI[455] HI[456] HI[457] HI[458] HI[459] HI[45] HI[460] HI[461] HI[462] HI[46]
+ HI[47] HI[48] HI[49] HI[4] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57]
+ HI[58] HI[59] HI[5] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68]
+ HI[69] HI[6] HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79]
+ HI[7] HI[80] HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8]
+ HI[90] HI[91] HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1
+ vssd1
.ends

* Black-box entry subcircuit for mgmt_protect_hv abstract view
.subckt mgmt_protect_hv mprj2_vdd_logic1 mprj_vdd_logic1 vccd vssd vdda1 vssa1 vdda2
+ vssa2
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102]
+ la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107]
+ la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[10] la_iena_mprj[110] la_iena_mprj[111]
+ la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116]
+ la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[11] la_iena_mprj[120]
+ la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125]
+ la_iena_mprj[126] la_iena_mprj[127] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14]
+ la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19]
+ la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23]
+ la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28]
+ la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32]
+ la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37]
+ la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3] la_iena_mprj[40] la_iena_mprj[41]
+ la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46]
+ la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[4] la_iena_mprj[50]
+ la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55]
+ la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[5]
+ la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64]
+ la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69]
+ la_iena_mprj[6] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73]
+ la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78]
+ la_iena_mprj[79] la_iena_mprj[7] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82]
+ la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87]
+ la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[8] la_iena_mprj[90] la_iena_mprj[91]
+ la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96]
+ la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[9] la_oenb_core[0]
+ la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104]
+ la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109]
+ la_oenb_core[10] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113]
+ la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118]
+ la_oenb_core[119] la_oenb_core[11] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122]
+ la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127]
+ la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16]
+ la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[1] la_oenb_core[20]
+ la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25]
+ la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[2]
+ la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34]
+ la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39]
+ la_oenb_core[3] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43]
+ la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48]
+ la_oenb_core[49] la_oenb_core[4] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52]
+ la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57]
+ la_oenb_core[58] la_oenb_core[59] la_oenb_core[5] la_oenb_core[60] la_oenb_core[61]
+ la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66]
+ la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[6] la_oenb_core[70]
+ la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75]
+ la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[7]
+ la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84]
+ la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89]
+ la_oenb_core[8] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93]
+ la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98]
+ la_oenb_core[99] la_oenb_core[9] la_oenb_mprj[0] la_oenb_mprj[100] la_oenb_mprj[101]
+ la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106]
+ la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[10] la_oenb_mprj[110]
+ la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115]
+ la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[11]
+ la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124]
+ la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] la_oenb_mprj[12] la_oenb_mprj[13]
+ la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18]
+ la_oenb_mprj[19] la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22]
+ la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27]
+ la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31]
+ la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36]
+ la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40]
+ la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45]
+ la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4]
+ la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54]
+ la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59]
+ la_oenb_mprj[5] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63]
+ la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68]
+ la_oenb_mprj[69] la_oenb_mprj[6] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72]
+ la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77]
+ la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[7] la_oenb_mprj[80] la_oenb_mprj[81]
+ la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86]
+ la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[8] la_oenb_mprj[90]
+ la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95]
+ la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[9]
+ mprj_ack_i_core mprj_ack_i_user mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11]
+ mprj_adr_o_core[12] mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15]
+ mprj_adr_o_core[16] mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19]
+ mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23]
+ mprj_adr_o_core[24] mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27]
+ mprj_adr_o_core[28] mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31]
+ mprj_adr_o_core[3] mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7]
+ mprj_adr_o_core[8] mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11]
+ mprj_adr_o_user[12] mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15]
+ mprj_adr_o_user[16] mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19]
+ mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23]
+ mprj_adr_o_user[24] mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27]
+ mprj_adr_o_user[28] mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31]
+ mprj_adr_o_user[3] mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7]
+ mprj_adr_o_user[8] mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0]
+ mprj_dat_i_core[10] mprj_dat_i_core[11] mprj_dat_i_core[12] mprj_dat_i_core[13]
+ mprj_dat_i_core[14] mprj_dat_i_core[15] mprj_dat_i_core[16] mprj_dat_i_core[17]
+ mprj_dat_i_core[18] mprj_dat_i_core[19] mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21]
+ mprj_dat_i_core[22] mprj_dat_i_core[23] mprj_dat_i_core[24] mprj_dat_i_core[25]
+ mprj_dat_i_core[26] mprj_dat_i_core[27] mprj_dat_i_core[28] mprj_dat_i_core[29]
+ mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31] mprj_dat_i_core[3] mprj_dat_i_core[4]
+ mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7] mprj_dat_i_core[8] mprj_dat_i_core[9]
+ mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11] mprj_dat_i_user[12] mprj_dat_i_user[13]
+ mprj_dat_i_user[14] mprj_dat_i_user[15] mprj_dat_i_user[16] mprj_dat_i_user[17]
+ mprj_dat_i_user[18] mprj_dat_i_user[19] mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21]
+ mprj_dat_i_user[22] mprj_dat_i_user[23] mprj_dat_i_user[24] mprj_dat_i_user[25]
+ mprj_dat_i_user[26] mprj_dat_i_user[27] mprj_dat_i_user[28] mprj_dat_i_user[29]
+ mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31] mprj_dat_i_user[3] mprj_dat_i_user[4]
+ mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7] mprj_dat_i_user[8] mprj_dat_i_user[9]
+ mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13]
+ mprj_dat_o_core[14] mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17]
+ mprj_dat_o_core[18] mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21]
+ mprj_dat_o_core[22] mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25]
+ mprj_dat_o_core[26] mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29]
+ mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4]
+ mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9]
+ mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13]
+ mprj_dat_o_user[14] mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17]
+ mprj_dat_o_user[18] mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21]
+ mprj_dat_o_user[22] mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25]
+ mprj_dat_o_user[26] mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29]
+ mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4]
+ mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9]
+ mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2] mprj_sel_o_core[3]
+ mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3] mprj_stb_o_core
+ mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood user1_vdd_powergood
+ user2_vcc_powergood user2_vdd_powergood user_clock user_clock2 user_irq[0] user_irq[1]
+ user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2] user_irq_ena[0] user_irq_ena[1]
+ user_irq_ena[2] user_reset vccd vccd1_uq1 vccd2_uq0 vdda1 vdda2 vssa1 vssa2 vssd
+ vssa2_uq0 vssa1_uq0 vdda2_uq0 vdda1_uq0 vssd2_uq0 vssd1_uq1
XFILLER_3_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1360 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1371 _343_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1382 _355_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1393 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1307 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_501_ _501_/A _501_/B vssd vssd vccd vccd _501_/X sky130_fd_sc_hd__and2_4
XANTENNA_202 _423_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_213 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_224 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 _434_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 _440_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1298 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_432_ _560_/A _432_/B _432_/C vssd vssd vccd vccd _432_/X sky130_fd_sc_hd__and3b_4
XFILLER_19_3677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_257 _441_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_268 _447_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_279 _449_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_363_ _363_/A _363_/B vssd vssd vccd vccd _363_/X sky130_fd_sc_hd__and2_4
XTAP_1888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_294_ _294_/A _294_/B vssd vssd vccd vccd _294_/X sky130_fd_sc_hd__and2_4
XFILLER_48_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[8\] mprj_dat_i_user[8] _294_/X vssd vssd vccd vccd _122_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_4327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_4051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4134 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_780 _603_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_791 _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[25\] la_data_out_core[25] _188_/X vssd vssd vccd vccd _008_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_36_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2402 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput467 _472_/X vssd vssd vccd vccd la_data_in_core[103] sky130_fd_sc_hd__buf_8
Xoutput478 _482_/X vssd vssd vccd vccd la_data_in_core[113] sky130_fd_sc_hd__buf_8
XFILLER_42_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput489 _492_/X vssd vssd vccd vccd la_data_in_core[123] sky130_fd_sc_hd__buf_8
XFILLER_47_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1190 _223_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_932 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_346 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4006 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_415_ _543_/A _415_/B _415_/C vssd vssd vccd vccd _415_/X sky130_fd_sc_hd__and3b_4
XTAP_2397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_346_ _346_/A _346_/B vssd vssd vccd vccd _346_/X sky130_fd_sc_hd__and2_4
XFILLER_35_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_277_ _277_/A _277_/B vssd vssd vccd vccd _277_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3854 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_200_ _200_/A _200_/B vssd vssd vccd vccd _200_/X sky130_fd_sc_hd__and2_2
XFILLER_19_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_131_ _131_/A vssd vssd vccd vccd _131_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_062_ _062_/A vssd vssd vccd vccd _062_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_4455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2605 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2616 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2627 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1904 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1915 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1926 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1937 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1948 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1959 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_329_ _329_/A _329_/B vssd vssd vccd vccd _329_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4522 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[92\] la_data_out_core[92] _255_/X vssd vssd vccd vccd _075_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_45_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_3680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1298 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_97 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3422 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_114_ _114_/A vssd vssd vccd vccd _114_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_045_ _045_/A vssd vssd vccd vccd _045_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_1630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2402 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2413 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2424 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2435 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2446 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1701 _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2457 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1712 _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1723 _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2468 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1734 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2479 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1745 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1756 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1767 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1778 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1789 _327_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[20\] mprj_dat_i_user[20] _294_/X vssd vssd vccd vccd _134_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_609 _511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_3910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1008 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1019 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput301 la_oenb_mprj[21] vssd vssd vccd vccd _518_/A sky130_fd_sc_hd__buf_6
Xinput312 la_oenb_mprj[31] vssd vssd vccd vccd _528_/A sky130_fd_sc_hd__buf_8
XFILLER_0_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput323 la_oenb_mprj[41] vssd vssd vccd vccd _538_/A sky130_fd_sc_hd__buf_4
XFILLER_44_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput334 la_oenb_mprj[51] vssd vssd vccd vccd _548_/A sky130_fd_sc_hd__buf_6
Xinput345 la_oenb_mprj[61] vssd vssd vccd vccd _558_/A sky130_fd_sc_hd__clkbuf_4
Xinput356 la_oenb_mprj[71] vssd vssd vccd vccd _568_/A sky130_fd_sc_hd__buf_8
Xinput367 la_oenb_mprj[81] vssd vssd vccd vccd _578_/A sky130_fd_sc_hd__buf_8
XFILLER_40_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput378 la_oenb_mprj[91] vssd vssd vccd vccd _588_/A sky130_fd_sc_hd__buf_6
Xinput389 mprj_adr_o_core[10] vssd vssd vccd vccd _315_/B sky130_fd_sc_hd__buf_8
XFILLER_2_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_594_ _594_/A _594_/B vssd vssd vccd vccd _594_/X sky130_fd_sc_hd__and2_4
XFILLER_35_4565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1774 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_5 la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput808 _562_/X vssd vssd vccd vccd la_oenb_core[65] sky130_fd_sc_hd__buf_8
XFILLER_29_3657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput819 _572_/X vssd vssd vccd vccd la_oenb_core[75] sky130_fd_sc_hd__buf_8
X_028_ _028_/A vssd vssd vccd vccd _028_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2210 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2221 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2232 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2243 _388_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2254 _555_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2265 _363_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1520 _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2276 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1531 _384_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2287 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1542 _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1553 _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2298 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1564 _392_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1575 _296_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1586 _492_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1597 _599_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[55\] la_data_out_core[55] _218_/X vssd vssd vccd vccd _038_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_48_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4516 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_406 _475_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_417 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_428 _479_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_439 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3751 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput120 la_data_out_mprj[8] vssd vssd vccd vccd _377_/C sky130_fd_sc_hd__clkbuf_4
Xinput131 la_data_out_mprj[9] vssd vssd vccd vccd _378_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput142 la_iena_mprj[109] vssd vssd vccd vccd _272_/B sky130_fd_sc_hd__clkbuf_4
Xinput153 la_iena_mprj[119] vssd vssd vccd vccd _282_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput164 la_iena_mprj[13] vssd vssd vccd vccd _176_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput175 la_iena_mprj[23] vssd vssd vccd vccd _186_/B sky130_fd_sc_hd__buf_4
XTAP_4652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput186 la_iena_mprj[33] vssd vssd vccd vccd _196_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput197 la_iena_mprj[43] vssd vssd vccd vccd _206_/B sky130_fd_sc_hd__buf_4
XFILLER_40_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_940 _621_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_951 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_962 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_577_ _577_/A _577_/B vssd vssd vccd vccd _577_/X sky130_fd_sc_hd__and2_4
XFILLER_32_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_973 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_984 _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_995 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput605 _095_/Y vssd vssd vccd vccd la_data_in_mprj[112] sky130_fd_sc_hd__buf_8
XFILLER_9_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput616 _105_/Y vssd vssd vccd vccd la_data_in_mprj[122] sky130_fd_sc_hd__buf_8
XFILLER_29_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput627 _000_/Y vssd vssd vccd vccd la_data_in_mprj[17] sky130_fd_sc_hd__buf_8
XFILLER_42_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput638 _010_/Y vssd vssd vccd vccd la_data_in_mprj[27] sky130_fd_sc_hd__buf_8
XFILLER_29_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput649 _020_/Y vssd vssd vccd vccd la_data_in_mprj[37] sky130_fd_sc_hd__buf_8
XFILLER_42_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2040 _318_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_2051 _353_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2062 output953/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2073 mprj_dat_i_user[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2084 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2095 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1350 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1361 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1372 _344_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1383 _356_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1394 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_602 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1076 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_500_ _500_/A _500_/B vssd vssd vccd vccd _500_/X sky130_fd_sc_hd__and2_4
XFILLER_22_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 _423_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_225 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_236 _435_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_602 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_431_ _559_/A _431_/B _431_/C vssd vssd vccd vccd _431_/X sky130_fd_sc_hd__and3b_4
XTAP_2557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 _440_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 _443_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 _447_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_362_ _362_/A _362_/B vssd vssd vccd vccd _362_/X sky130_fd_sc_hd__and2_4
XFILLER_14_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_293_ _293_/A _293_/B vssd vssd vccd vccd _293_/X sky130_fd_sc_hd__and2_1
XFILLER_42_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1891 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4146 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_770 _599_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_781 _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_792 _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[18\] la_data_out_core[18] _181_/X vssd vssd vccd vccd _001_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_9_4013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput468 _473_/X vssd vssd vccd vccd la_data_in_core[104] sky130_fd_sc_hd__buf_8
Xoutput479 _483_/X vssd vssd vccd vccd la_data_in_core[114] sky130_fd_sc_hd__buf_8
XFILLER_42_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1998 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1180 _216_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1191 _226_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_4107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_3597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3671 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_270 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_414_ _542_/A _414_/B _414_/C vssd vssd vccd vccd _414_/X sky130_fd_sc_hd__and3b_4
XTAP_2387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_345_ _345_/A _345_/B vssd vssd vccd vccd _345_/X sky130_fd_sc_hd__and2_4
XFILLER_50_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_276_ _276_/A _276_/B vssd vssd vccd vccd _276_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4147 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2723 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3866 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_130_ _130_/A vssd vssd vccd vccd _130_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_1071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_061_ _061_/A vssd vssd vccd vccd _061_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2606 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2617 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2628 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1905 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1916 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1927 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1938 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1949 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_328_ _328_/A _328_/B vssd vssd vccd vccd _328_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_259_ _259_/A _259_/B vssd vssd vccd vccd _259_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[85\] la_data_out_core[85] _248_/X vssd vssd vccd vccd _068_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_3971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_516 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_113_ _113_/A vssd vssd vccd vccd _113_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_044_ _044_/A vssd vssd vccd vccd _044_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_27_4231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2403 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2414 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2425 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2436 _357_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1702 _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2447 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2458 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1713 _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1724 _321_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2469 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1735 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1746 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1757 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1768 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1779 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[13\] mprj_dat_i_user[13] _294_/X vssd vssd vccd vccd _127_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[111\] la_data_out_core[111] _274_/X vssd vssd vccd vccd _094_/A
+ sky130_fd_sc_hd__nand2_8
XTAP_2909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_4379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1009 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput302 la_oenb_mprj[22] vssd vssd vccd vccd _519_/A sky130_fd_sc_hd__buf_4
XFILLER_22_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput313 la_oenb_mprj[32] vssd vssd vccd vccd _529_/A sky130_fd_sc_hd__buf_6
Xinput324 la_oenb_mprj[42] vssd vssd vccd vccd _539_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput335 la_oenb_mprj[52] vssd vssd vccd vccd _549_/A sky130_fd_sc_hd__buf_4
Xinput346 la_oenb_mprj[62] vssd vssd vccd vccd _559_/A sky130_fd_sc_hd__buf_6
Xinput357 la_oenb_mprj[72] vssd vssd vccd vccd _569_/A sky130_fd_sc_hd__buf_8
Xinput368 la_oenb_mprj[82] vssd vssd vccd vccd _579_/A sky130_fd_sc_hd__buf_8
XFILLER_5_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput379 la_oenb_mprj[92] vssd vssd vccd vccd _589_/A sky130_fd_sc_hd__buf_6
XFILLER_18_4208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_593_ _593_/A _593_/B vssd vssd vccd vccd _593_/X sky130_fd_sc_hd__and2_4
XFILLER_21_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_6 la_data_out_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput809 _563_/X vssd vssd vccd vccd la_oenb_core[66] sky130_fd_sc_hd__buf_8
XFILLER_42_4515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_027_ _027_/A vssd vssd vccd vccd _027_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_4526 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2200 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2211 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2222 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2233 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2244 _455_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1510 _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2255 _586_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1521 _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2266 _364_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2277 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1532 _384_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2288 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1543 _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2299 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1554 _387_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1565 _392_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1576 _296_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1587 _493_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1598 _599_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[48\] la_data_out_core[48] _211_/X vssd vssd vccd vccd _031_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_34_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_407 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_418 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_429 _479_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3475 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3763 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput110 la_data_out_mprj[80] vssd vssd vccd vccd _449_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_24_3588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput121 la_data_out_mprj[90] vssd vssd vccd vccd _459_/C sky130_fd_sc_hd__clkbuf_4
Xinput132 la_iena_mprj[0] vssd vssd vccd vccd _625_/B sky130_fd_sc_hd__clkbuf_4
Xinput143 la_iena_mprj[10] vssd vssd vccd vccd _173_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput154 la_iena_mprj[11] vssd vssd vccd vccd _174_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput165 la_iena_mprj[14] vssd vssd vccd vccd _177_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput176 la_iena_mprj[24] vssd vssd vccd vccd _187_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1050 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput187 la_iena_mprj[34] vssd vssd vccd vccd _197_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput198 la_iena_mprj[44] vssd vssd vccd vccd _207_/B sky130_fd_sc_hd__buf_4
XFILLER_36_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_930 _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_941 _621_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_576_ _576_/A _576_/B vssd vssd vccd vccd _576_/X sky130_fd_sc_hd__and2_4
XANTENNA_952 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_963 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_974 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_985 _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_996 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput606 _096_/Y vssd vssd vccd vccd la_data_in_mprj[113] sky130_fd_sc_hd__buf_8
Xoutput617 _106_/Y vssd vssd vccd vccd la_data_in_mprj[123] sky130_fd_sc_hd__buf_8
XFILLER_25_3308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput628 _001_/Y vssd vssd vccd vccd la_data_in_mprj[18] sky130_fd_sc_hd__buf_8
Xoutput639 _011_/Y vssd vssd vccd vccd la_data_in_mprj[28] sky130_fd_sc_hd__buf_8
XFILLER_29_2754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2030 _300_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2041 _319_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2052 _355_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2063 output953/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2074 _419_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1340 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2085 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2096 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1351 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1362 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1373 _299_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1384 _359_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1395 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2026 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3795 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_226 _425_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 _435_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_430_ _558_/A _430_/B _430_/C vssd vssd vccd vccd _430_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_4514 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_248 _440_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_614 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_259 _445_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_361_ _361_/A _361_/B vssd vssd vccd vccd _361_/X sky130_fd_sc_hd__and2_4
XFILLER_13_3212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_292_ _292_/A _292_/B vssd vssd vccd vccd _292_/X sky130_fd_sc_hd__and2_1
XFILLER_42_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4158 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_760 _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_771 _600_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_782 _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_559_ _559_/A _559_/B vssd vssd vccd vccd _559_/X sky130_fd_sc_hd__and2_4
XANTENNA_793 _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1954 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput469 _474_/X vssd vssd vccd vccd la_data_in_core[105] sky130_fd_sc_hd__buf_8
XFILLER_47_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1170 _211_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1181 _217_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1192 _226_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4271 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1242 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2198 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3514 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3683 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3476 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_413_ _541_/A _413_/B _413_/C vssd vssd vccd vccd _413_/X sky130_fd_sc_hd__and3b_4
XFILLER_26_282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_344_ _344_/A _344_/B vssd vssd vccd vccd _344_/X sky130_fd_sc_hd__and2_4
XFILLER_35_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_275_ _275_/A _275_/B vssd vssd vccd vccd _275_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2702 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2807 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2735 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4542 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[30\] la_data_out_core[30] _193_/X vssd vssd vccd vccd _013_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_33_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_590 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3878 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1083 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_060_ _060_/A vssd vssd vccd vccd _060_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2607 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2618 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2629 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1906 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1917 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_178 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1928 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1939 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_327_ _327_/A _327_/B vssd vssd vccd vccd _327_/X sky130_fd_sc_hd__and2_4
XFILLER_15_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_258_ _258_/A _258_/B vssd vssd vccd vccd _258_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_189_ _189_/A _189_/B vssd vssd vccd vccd _189_/X sky130_fd_sc_hd__and2_2
XFILLER_45_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[78\] la_data_out_core[78] _241_/X vssd vssd vccd vccd _061_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_4_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_112_ _112_/A vssd vssd vccd vccd _112_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_043_ _043_/A vssd vssd vccd vccd _043_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2404 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2415 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2426 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2437 _358_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2448 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1703 _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1714 _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2459 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2863 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1725 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1736 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1747 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1758 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1769 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_4280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[104\] la_data_out_core[104] _267_/X vssd vssd vccd vccd _087_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_52_100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput303 la_oenb_mprj[23] vssd vssd vccd vccd _520_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput314 la_oenb_mprj[33] vssd vssd vccd vccd _530_/A sky130_fd_sc_hd__buf_4
XFILLER_22_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput325 la_oenb_mprj[43] vssd vssd vccd vccd _540_/A sky130_fd_sc_hd__buf_8
Xinput336 la_oenb_mprj[53] vssd vssd vccd vccd _550_/A sky130_fd_sc_hd__buf_4
XFILLER_40_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput347 la_oenb_mprj[63] vssd vssd vccd vccd _560_/A sky130_fd_sc_hd__buf_6
Xinput358 la_oenb_mprj[73] vssd vssd vccd vccd _570_/A sky130_fd_sc_hd__buf_8
XFILLER_2_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput369 la_oenb_mprj[83] vssd vssd vccd vccd _580_/A sky130_fd_sc_hd__buf_8
XFILLER_28_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_592_ _592_/A _592_/B vssd vssd vccd vccd _592_/X sky130_fd_sc_hd__and2_4
XFILLER_38_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3298 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_7 la_data_out_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_026_ _026_/A vssd vssd vccd vccd _026_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_4538 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2201 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2212 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2223 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2234 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2245 _598_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1500 _379_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1511 _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2256 _595_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2267 _365_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1522 _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2278 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1533 _384_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1544 _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2289 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1555 _387_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3010 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1566 _392_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1577 _296_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1588 _495_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1599 _600_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1839 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_408 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_419 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4020 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput100 la_data_out_mprj[71] vssd vssd vccd vccd _440_/C sky130_fd_sc_hd__buf_6
XFILLER_24_2833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput111 la_data_out_mprj[81] vssd vssd vccd vccd _450_/C sky130_fd_sc_hd__buf_6
XFILLER_24_2844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput122 la_data_out_mprj[91] vssd vssd vccd vccd _460_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput133 la_iena_mprj[100] vssd vssd vccd vccd _263_/B sky130_fd_sc_hd__clkbuf_4
Xinput144 la_iena_mprj[110] vssd vssd vccd vccd _273_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput155 la_iena_mprj[120] vssd vssd vccd vccd _283_/B sky130_fd_sc_hd__buf_4
XTAP_4632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput166 la_iena_mprj[15] vssd vssd vccd vccd _178_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput177 la_iena_mprj[25] vssd vssd vccd vccd _188_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput188 la_iena_mprj[35] vssd vssd vccd vccd _198_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput199 la_iena_mprj[45] vssd vssd vccd vccd _208_/B sky130_fd_sc_hd__buf_4
XFILLER_29_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_920 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_931 _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_575_ _575_/A _575_/B vssd vssd vccd vccd _575_/X sky130_fd_sc_hd__and2_4
XANTENNA_942 _621_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_953 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_964 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_975 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_986 _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_997 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_354 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput607 _097_/Y vssd vssd vccd vccd la_data_in_mprj[114] sky130_fd_sc_hd__buf_8
XFILLER_9_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput618 _107_/Y vssd vssd vccd vccd la_data_in_mprj[124] sky130_fd_sc_hd__buf_8
Xoutput629 _002_/Y vssd vssd vccd vccd la_data_in_mprj[19] sky130_fd_sc_hd__buf_8
X_009_ _009_/A vssd vssd vccd vccd _009_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2020 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2031 _469_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2042 _322_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2053 _357_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2064 output953/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2075 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1330 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2086 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1341 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2097 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1352 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1363 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1374 _345_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[60\] la_data_out_core[60] _223_/X vssd vssd vccd vccd _043_/A
+ sky130_fd_sc_hd__nand2_2
XANTENNA_1385 _361_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1396 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_626 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4150 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_4408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1564 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1130 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_216 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_227 _425_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 _435_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 _440_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4526 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_626 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_360_ _360_/A _360_/B vssd vssd vccd vccd _360_/X sky130_fd_sc_hd__and2_4
XFILLER_17_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_291_ _291_/A _291_/B vssd vssd vccd vccd _291_/X sky130_fd_sc_hd__and2_1
XFILLER_52_3295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1052 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_750 _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_761 _598_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_772 _601_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_558_ _558_/A _558_/B vssd vssd vccd vccd _558_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_783 _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_794 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_489_ _617_/A _489_/B _489_/C vssd vssd vccd vccd _489_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3314 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1923 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_4452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1160 _199_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1171 _212_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3740 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1182 _217_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1193 _227_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3878 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1254 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1476 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput960 _295_/X vssd vssd vccd vccd user_reset sky130_fd_sc_hd__buf_8
XFILLER_5_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_412_ _540_/A _412_/B _412_/C vssd vssd vccd vccd _412_/X sky130_fd_sc_hd__and3b_4
XTAP_2367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_343_ _343_/A _343_/B vssd vssd vccd vccd _343_/X sky130_fd_sc_hd__and2_4
XTAP_1677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_274_ _274_/A _274_/B vssd vssd vccd vccd _274_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[6\] mprj_dat_i_user[6] _294_/X vssd vssd vccd vccd _120_/A sky130_fd_sc_hd__nand2_2
XFILLER_48_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_850 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2747 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_580 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_591 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[23\] la_data_out_core[23] _186_/X vssd vssd vccd vccd _006_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_36_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1858 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2608 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2619 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1907 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1918 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput790 _546_/X vssd vssd vccd vccd la_oenb_core[49] sky130_fd_sc_hd__buf_8
XANTENNA_1929 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_326_ _326_/A _326_/B vssd vssd vccd vccd _326_/X sky130_fd_sc_hd__and2_4
XFILLER_9_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_257_ _257_/A _257_/B vssd vssd vccd vccd _257_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_188_ _188_/A _188_/B vssd vssd vccd vccd _188_/X sky130_fd_sc_hd__and2_2
XFILLER_7_986 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_89 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_111_ _111_/A vssd vssd vccd vccd _111_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_042_ _042_/A vssd vssd vccd vccd _042_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2405 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2416 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2831 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2427 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_4051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2438 _360_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2449 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1704 _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1715 _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1726 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2875 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1737 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1748 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1759 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3236 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_309_ _309_/A _309_/B vssd vssd vccd vccd _309_/X sky130_fd_sc_hd__and2_2
XFILLER_30_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[90\] la_data_out_core[90] _253_/X vssd vssd vccd vccd _073_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_28_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1076 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput304 la_oenb_mprj[24] vssd vssd vccd vccd _521_/A sky130_fd_sc_hd__buf_4
XFILLER_40_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput315 la_oenb_mprj[34] vssd vssd vccd vccd _531_/A sky130_fd_sc_hd__buf_4
XFILLER_44_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput326 la_oenb_mprj[44] vssd vssd vccd vccd _541_/A sky130_fd_sc_hd__buf_4
XFILLER_22_4196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput337 la_oenb_mprj[54] vssd vssd vccd vccd _551_/A sky130_fd_sc_hd__buf_6
XFILLER_29_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput348 la_oenb_mprj[64] vssd vssd vccd vccd _561_/A sky130_fd_sc_hd__buf_6
XFILLER_40_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput359 la_oenb_mprj[74] vssd vssd vccd vccd _571_/A sky130_fd_sc_hd__buf_8
XFILLER_29_621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_654 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_591_ _591_/A _591_/B vssd vssd vccd vccd _591_/X sky130_fd_sc_hd__and2_4
XFILLER_35_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_025_ _025_/A vssd vssd vccd vccd _025_/Y sky130_fd_sc_hd__inv_2
XANTENNA_8 la_data_out_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4063 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2202 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2213 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2224 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2235 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2246 _600_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1501 _379_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1512 _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3478 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2257 _596_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2268 _366_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1523 _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2279 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1534 _384_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1545 _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1556 _387_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1567 _392_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1578 _296_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1589 _496_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_409 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_432 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3764 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput101 la_data_out_mprj[72] vssd vssd vccd vccd _441_/C sky130_fd_sc_hd__buf_4
XFILLER_7_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput112 la_data_out_mprj[82] vssd vssd vccd vccd _451_/C sky130_fd_sc_hd__buf_6
Xinput123 la_data_out_mprj[92] vssd vssd vccd vccd _461_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput134 la_iena_mprj[101] vssd vssd vccd vccd _264_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_4076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput145 la_iena_mprj[111] vssd vssd vccd vccd _274_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput156 la_iena_mprj[121] vssd vssd vccd vccd _284_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput167 la_iena_mprj[16] vssd vssd vccd vccd _179_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput178 la_iena_mprj[26] vssd vssd vccd vccd _189_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 la_iena_mprj[36] vssd vssd vccd vccd _199_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_4018 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_910 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_921 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_574_ _574_/A _574_/B vssd vssd vccd vccd _574_/X sky130_fd_sc_hd__and2_4
XANTENNA_932 _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_943 _621_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_954 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_965 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_976 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_987 _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_998 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput608 _098_/Y vssd vssd vccd vccd la_data_in_mprj[115] sky130_fd_sc_hd__buf_8
Xoutput619 _108_/Y vssd vssd vccd vccd la_data_in_mprj[125] sky130_fd_sc_hd__buf_8
X_008_ _008_/A vssd vssd vccd vccd _008_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2010 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2021 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2032 _414_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2043 _325_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2054 _362_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2065 output954/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1320 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1331 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2076 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2087 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1342 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2098 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1353 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1364 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1375 _346_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1386 _362_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1397 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[53\] la_data_out_core[53] _216_/X vssd vssd vccd vccd _036_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_48_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1068 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4280 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_228 _429_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_239 _435_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4538 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_290_ _290_/A _290_/B vssd vssd vccd vccd _290_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_740 _595_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_751 _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_762 _598_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_557_ _557_/A _557_/B vssd vssd vccd vccd _557_/X sky130_fd_sc_hd__and2_4
XANTENNA_773 _603_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_784 _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_795 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_488_ _616_/A _488_/B _488_/C vssd vssd vccd vccd _488_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3326 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1150 _197_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1161 _200_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1172 _332_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1183 _219_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1194 _227_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1266 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput950 _300_/X vssd vssd vccd vccd mprj_we_o_user sky130_fd_sc_hd__buf_8
XFILLER_25_4375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_411_ _539_/A _411_/B _411_/C vssd vssd vccd vccd _411_/X sky130_fd_sc_hd__and3b_4
XFILLER_14_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_342_ _342_/A _342_/B vssd vssd vccd vccd _342_/X sky130_fd_sc_hd__and2_4
XTAP_1678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_273_ _273_/A _273_/B vssd vssd vccd vccd _273_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_609_ _609_/A _609_/B vssd vssd vccd vccd _609_/X sky130_fd_sc_hd__and2_4
XFILLER_17_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_570 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_581 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_592 _507_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[16\] la_data_out_core[16] _179_/X vssd vssd vccd vccd _163_/A
+ sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_gates\[29\] mprj_dat_i_user[29] _294_/X vssd vssd vccd vccd _143_/A sky130_fd_sc_hd__nand2_2
XFILLER_31_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2422 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1743 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[127\] la_data_out_core[127] _290_/X vssd vssd vccd vccd _110_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_0_4355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2609 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1908 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput780 _500_/X vssd vssd vccd vccd la_oenb_core[3] sky130_fd_sc_hd__buf_8
XANTENNA_1919 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput791 _501_/X vssd vssd vccd vccd la_oenb_core[4] sky130_fd_sc_hd__buf_8
XFILLER_40_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_325_ _325_/A _325_/B vssd vssd vccd vccd _325_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_256_ _256_/A _256_/B vssd vssd vccd vccd _256_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_187_ _187_/A _187_/B vssd vssd vccd vccd _187_/X sky130_fd_sc_hd__and2_2
XFILLER_48_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_110_ _110_/A vssd vssd vccd vccd _110_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_041_ _041_/A vssd vssd vccd vccd _041_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2406 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2417 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2428 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2439 _366_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1705 _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1716 _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1727 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1738 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2887 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1749 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_308_ _308_/A _308_/B vssd vssd vccd vccd _308_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_239_ _239_/A _239_/B vssd vssd vccd vccd _239_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3126 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[83\] la_data_out_core[83] _246_/X vssd vssd vccd vccd _066_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_44_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_828 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3746 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_3914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1998 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput305 la_oenb_mprj[25] vssd vssd vccd vccd _522_/A sky130_fd_sc_hd__buf_4
XFILLER_2_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput316 la_oenb_mprj[35] vssd vssd vccd vccd _532_/A sky130_fd_sc_hd__buf_6
XFILLER_22_3441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput327 la_oenb_mprj[45] vssd vssd vccd vccd _542_/A sky130_fd_sc_hd__buf_4
XFILLER_22_3452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput338 la_oenb_mprj[55] vssd vssd vccd vccd _552_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput349 la_oenb_mprj[65] vssd vssd vccd vccd _562_/A sky130_fd_sc_hd__buf_6
XFILLER_29_600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_590_ _590_/A _590_/B vssd vssd vccd vccd _590_/X sky130_fd_sc_hd__and2_4
XFILLER_28_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_382 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_024_ _024_/A vssd vssd vccd vccd _024_/Y sky130_fd_sc_hd__inv_2
XANTENNA_9 la_data_out_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_2187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4075 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4158 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2203 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2214 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2225 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2236 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1502 _380_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2247 _602_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1513 _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2258 _362_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2269 _339_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1524 _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1535 _384_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1546 _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2695 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1557 _387_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1568 _394_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1579 _296_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[11\] mprj_dat_i_user[11] _294_/X vssd vssd vccd vccd _125_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_614 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_488 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput102 la_data_out_mprj[73] vssd vssd vccd vccd _442_/C sky130_fd_sc_hd__buf_4
XFILLER_24_2835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput113 la_data_out_mprj[83] vssd vssd vccd vccd _452_/C sky130_fd_sc_hd__buf_6
XFILLER_7_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput124 la_data_out_mprj[93] vssd vssd vccd vccd _462_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput135 la_iena_mprj[102] vssd vssd vccd vccd _265_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput146 la_iena_mprj[112] vssd vssd vccd vccd _275_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput157 la_iena_mprj[122] vssd vssd vccd vccd _285_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput168 la_iena_mprj[17] vssd vssd vccd vccd _180_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput179 la_iena_mprj[27] vssd vssd vccd vccd _190_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_29_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_900 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_911 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_573_ _573_/A _573_/B vssd vssd vccd vccd _573_/X sky130_fd_sc_hd__and2_4
XANTENNA_922 _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_933 _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_944 _621_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_955 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_966 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_977 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_988 _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_999 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput609 _099_/Y vssd vssd vccd vccd la_data_in_mprj[116] sky130_fd_sc_hd__buf_8
XFILLER_29_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_007_ _007_/A vssd vssd vccd vccd _007_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2000 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2011 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2022 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2033 _425_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2044 _311_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2055 _344_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1310 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2066 _069_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1321 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2077 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1332 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2088 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1343 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1354 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2099 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1365 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1376 _347_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1387 _363_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1398 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[46\] la_data_out_core[46] _209_/X vssd vssd vccd vccd _029_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[8\] la_data_out_core[8] _171_/X vssd vssd vccd vccd _155_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_25_3845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_4292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_207 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_229 _430_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_625_ _625_/A _625_/B vssd vssd vccd vccd _625_/X sky130_fd_sc_hd__and2_1
XTAP_3763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_730 _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_741 _595_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_752 _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_556_ _556_/A _556_/B vssd vssd vccd vccd _556_/X sky130_fd_sc_hd__and2_4
XFILLER_45_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_763 _598_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_774 _603_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_785 _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_796 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_487_ _615_/A _487_/B _487_/C vssd vssd vccd vccd _487_/X sky130_fd_sc_hd__and3b_4
XFILLER_38_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3338 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2604 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1080 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4410 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1140 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1151 _197_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1162 _201_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1173 _213_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1184 _219_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1195 _228_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_4361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4490 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput940 _342_/X vssd vssd vccd vccd mprj_dat_o_user[5] sky130_fd_sc_hd__buf_8
XFILLER_5_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput951 output951/A vssd vssd vccd vccd user1_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_25_4387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_410_ _538_/A _410_/B _410_/C vssd vssd vccd vccd _410_/X sky130_fd_sc_hd__and3b_4
XTAP_2347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_341_ _341_/A _341_/B vssd vssd vccd vccd _341_/X sky130_fd_sc_hd__and2_4
XFILLER_36_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_272_ _272_/A _272_/B vssd vssd vccd vccd _272_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_608_ _608_/A _608_/B vssd vssd vccd vccd _608_/X sky130_fd_sc_hd__and2_4
XTAP_3593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_560 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_571 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_582 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_539_ _539_/A _539_/B vssd vssd vccd vccd _539_/X sky130_fd_sc_hd__and2_4
XTAP_2892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_593 _510_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1711 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1766 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1909 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput770 _527_/X vssd vssd vccd vccd la_oenb_core[30] sky130_fd_sc_hd__buf_8
Xoutput781 _537_/X vssd vssd vccd vccd la_oenb_core[40] sky130_fd_sc_hd__buf_8
XFILLER_47_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput792 _547_/X vssd vssd vccd vccd la_oenb_core[50] sky130_fd_sc_hd__buf_8
XFILLER_21_3314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_324_ _324_/A _324_/B vssd vssd vccd vccd _324_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_255_ _255_/A _255_/B vssd vssd vccd vccd _255_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_186_ _186_/A _186_/B vssd vssd vccd vccd _186_/X sky130_fd_sc_hd__and2_1
XFILLER_7_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_682 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_390 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_040_ _040_/A vssd vssd vccd vccd _040_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2407 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2418 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2429 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1706 _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1717 _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1728 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1739 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_542 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_307_ _307_/A _307_/B vssd vssd vccd vccd _307_/X sky130_fd_sc_hd__and2_2
XFILLER_50_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_238_ _238_/A _238_/B vssd vssd vccd vccd _238_/X sky130_fd_sc_hd__and2_4
XFILLER_45_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_169_ _169_/A _169_/B vssd vssd vccd vccd _169_/X sky130_fd_sc_hd__and2_4
XFILLER_13_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[76\] la_data_out_core[76] _239_/X vssd vssd vccd vccd _059_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_23_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1170 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2072 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput306 la_oenb_mprj[26] vssd vssd vccd vccd _523_/A sky130_fd_sc_hd__buf_4
Xinput317 la_oenb_mprj[36] vssd vssd vccd vccd _533_/A sky130_fd_sc_hd__buf_8
XFILLER_2_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput328 la_oenb_mprj[46] vssd vssd vccd vccd _543_/A sky130_fd_sc_hd__buf_8
Xinput339 la_oenb_mprj[56] vssd vssd vccd vccd _553_/A sky130_fd_sc_hd__buf_4
XFILLER_22_3464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_023_ _023_/A vssd vssd vccd vccd _023_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2204 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2215 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2226 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2237 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1503 _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2248 _615_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1514 _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2259 _363_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1525 _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1536 _384_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1547 _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1558 _390_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1569 _394_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3068 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2334 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[102\] la_data_out_core[102] _265_/X vssd vssd vccd vccd _085_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_626 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput103 la_data_out_mprj[74] vssd vssd vccd vccd _443_/C sky130_fd_sc_hd__clkbuf_4
Xinput114 la_data_out_mprj[84] vssd vssd vccd vccd _453_/C sky130_fd_sc_hd__buf_8
XFILLER_49_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput125 la_data_out_mprj[94] vssd vssd vccd vccd _463_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput136 la_iena_mprj[103] vssd vssd vccd vccd _266_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput147 la_iena_mprj[113] vssd vssd vccd vccd _276_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput158 la_iena_mprj[123] vssd vssd vccd vccd _286_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput169 la_iena_mprj[18] vssd vssd vccd vccd _181_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_901 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_912 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_572_ _572_/A _572_/B vssd vssd vccd vccd _572_/X sky130_fd_sc_hd__and2_4
XFILLER_29_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_923 _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_934 _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_945 _621_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_956 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_967 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_978 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_989 _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_346 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_006_ _006_/A vssd vssd vccd vccd _006_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2001 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2758 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2012 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2023 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2034 _427_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2045 _314_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1300 _280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2056 _346_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1311 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1322 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2067 _070_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2078 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1333 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2089 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1344 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1355 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1366 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1377 _349_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1388 _364_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1399 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3711 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[39\] la_data_out_core[39] _202_/X vssd vssd vccd vccd _022_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_22_117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3728 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2590 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_219 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_624_ _624_/A _624_/B vssd vssd vccd vccd _624_/X sky130_fd_sc_hd__and2_4
XTAP_4498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_720 _594_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_731 _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_555_ _555_/A _555_/B vssd vssd vccd vccd _555_/X sky130_fd_sc_hd__and2_4
XANTENNA_742 _595_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_753 _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_764 _598_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_775 _603_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_786 _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_486_ _614_/A _486_/B _486_/C vssd vssd vccd vccd _486_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_797 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4018 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1130 _186_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1141 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2290 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1152 _197_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1163 _201_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1174 _214_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1185 _220_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1196 _228_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput930 _362_/X vssd vssd vccd vccd mprj_dat_o_user[25] sky130_fd_sc_hd__buf_8
XFILLER_25_4355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput941 _343_/X vssd vssd vccd vccd mprj_dat_o_user[6] sky130_fd_sc_hd__buf_8
XFILLER_9_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput952 output952/A vssd vssd vccd vccd user1_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_28_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2931 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_710 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_340_ _340_/A _340_/B vssd vssd vccd vccd _340_/X sky130_fd_sc_hd__and2_4
XFILLER_39_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_271_ _271_/A _271_/B vssd vssd vccd vccd _271_/X sky130_fd_sc_hd__and2_4
XFILLER_39_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4040 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_607_ _607_/A _607_/B vssd vssd vccd vccd _607_/X sky130_fd_sc_hd__and2_4
XFILLER_45_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_550 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_561 _499_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_572 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_538_ _538_/A _538_/B vssd vssd vccd vccd _538_/X sky130_fd_sc_hd__and2_4
XTAP_2893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_583 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_594 _510_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_469_ _597_/A _469_/B _469_/C vssd vssd vccd vccd _469_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_470 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1290 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_234 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3727 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput760 _518_/X vssd vssd vccd vccd la_oenb_core[21] sky130_fd_sc_hd__buf_8
XFILLER_5_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput771 _528_/X vssd vssd vccd vccd la_oenb_core[31] sky130_fd_sc_hd__buf_8
XFILLER_40_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput782 _538_/X vssd vssd vccd vccd la_oenb_core[41] sky130_fd_sc_hd__buf_8
XFILLER_8_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput793 _548_/X vssd vssd vccd vccd la_oenb_core[51] sky130_fd_sc_hd__buf_8
XFILLER_47_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_323_ _323_/A _323_/B vssd vssd vccd vccd _323_/X sky130_fd_sc_hd__and2_4
XFILLER_42_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_254_ _254_/A _254_/B vssd vssd vccd vccd _254_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_185_ _185_/A _185_/B vssd vssd vccd vccd _185_/X sky130_fd_sc_hd__and2_2
XFILLER_13_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[4\] mprj_dat_i_user[4] _294_/X vssd vssd vccd vccd _118_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_380 _469_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_391 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[21\] la_data_out_core[21] _184_/X vssd vssd vccd vccd _004_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_15_3664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3707 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2408 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2419 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1707 _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1718 _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput590 _378_/X vssd vssd vccd vccd la_data_in_core[9] sky130_fd_sc_hd__buf_8
XFILLER_44_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1729 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_306_ _306_/A _306_/B vssd vssd vccd vccd _306_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_237_ _237_/A _237_/B vssd vssd vccd vccd _237_/X sky130_fd_sc_hd__and2_4
XFILLER_45_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_168_ _168_/A _168_/B vssd vssd vccd vccd _168_/X sky130_fd_sc_hd__and2_4
XFILLER_45_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_099_ _099_/A vssd vssd vccd vccd _099_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_3034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[69\] la_data_out_core[69] _232_/X vssd vssd vccd vccd _052_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_39_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_104 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1182 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput307 la_oenb_mprj[27] vssd vssd vccd vccd _524_/A sky130_fd_sc_hd__buf_6
XFILLER_22_3432 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput318 la_oenb_mprj[37] vssd vssd vccd vccd _534_/A sky130_fd_sc_hd__buf_8
Xinput329 la_oenb_mprj[47] vssd vssd vccd vccd _544_/A sky130_fd_sc_hd__buf_8
XFILLER_25_1131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_022_ _022_/A vssd vssd vccd vccd _022_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2205 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2216 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2227 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2238 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2249 _619_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1504 _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1515 _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1526 _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1537 _384_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1548 _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1559 _390_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3792 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_4420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1716 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1764 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput104 la_data_out_mprj[75] vssd vssd vccd vccd _444_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput115 la_data_out_mprj[85] vssd vssd vccd vccd _454_/C sky130_fd_sc_hd__buf_8
Xinput126 la_data_out_mprj[95] vssd vssd vccd vccd _464_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput137 la_iena_mprj[104] vssd vssd vccd vccd _267_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput148 la_iena_mprj[114] vssd vssd vccd vccd _277_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput159 la_iena_mprj[124] vssd vssd vccd vccd _287_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_571_ _571_/A _571_/B vssd vssd vccd vccd _571_/X sky130_fd_sc_hd__and2_4
XANTENNA_902 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_913 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_924 _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_935 _621_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_946 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_957 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_968 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_979 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3970 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_005_ _005_/A vssd vssd vccd vccd _005_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2002 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2013 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2024 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2035 _465_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2046 _347_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1301 _280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2057 _304_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1312 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2068 _073_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1323 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2079 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1334 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1345 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1356 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1367 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1378 _350_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1389 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3707 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2580 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2591 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1890 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_623_ _623_/A _623_/B vssd vssd vccd vccd _623_/X sky130_fd_sc_hd__and2_4
XFILLER_29_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_710 _588_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_721 _594_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_554_ _554_/A _554_/B vssd vssd vccd vccd _554_/X sky130_fd_sc_hd__and2_4
XANTENNA_732 _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_743 _595_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_754 _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_765 _598_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_776 _603_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_485_ _613_/A _485_/B _485_/C vssd vssd vccd vccd _485_/X sky130_fd_sc_hd__and3b_4
XANTENNA_787 _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_798 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1120 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1131 _188_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1142 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1153 _197_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1164 _331_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1175 _214_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1186 _220_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1197 _229_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[51\] la_data_out_core[51] _214_/X vssd vssd vccd vccd _034_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_40_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput920 _353_/X vssd vssd vccd vccd mprj_dat_o_user[16] sky130_fd_sc_hd__buf_8
XFILLER_5_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput931 _363_/X vssd vssd vccd vccd mprj_dat_o_user[26] sky130_fd_sc_hd__buf_8
XFILLER_28_2033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput942 _344_/X vssd vssd vccd vccd mprj_dat_o_user[7] sky130_fd_sc_hd__buf_8
XFILLER_25_4367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput953 output953/A vssd vssd vccd vccd user2_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_45_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2943 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_298 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_270_ _270_/A _270_/B vssd vssd vccd vccd _270_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_606_ _606_/A _606_/B vssd vssd vccd vccd _606_/X sky130_fd_sc_hd__and2_4
XTAP_3573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_540 _496_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_551 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_562 _499_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_537_ _537_/A _537_/B vssd vssd vccd vccd _537_/X sky130_fd_sc_hd__and2_4
XTAP_2872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_573 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_584 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_595 _510_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_468_ _596_/A _468_/B _468_/C vssd vssd vccd vccd _468_/X sky130_fd_sc_hd__and3b_4
XFILLER_20_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_482 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_399_ _527_/A _399_/B _399_/C vssd vssd vccd vccd _399_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[99\] la_data_out_core[99] _262_/X vssd vssd vccd vccd _082_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_29_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3739 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4006 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput750 _509_/X vssd vssd vccd vccd la_oenb_core[12] sky130_fd_sc_hd__buf_8
Xoutput761 _519_/X vssd vssd vccd vccd la_oenb_core[22] sky130_fd_sc_hd__buf_8
Xoutput772 _529_/X vssd vssd vccd vccd la_oenb_core[32] sky130_fd_sc_hd__buf_8
XFILLER_5_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput783 _539_/X vssd vssd vccd vccd la_oenb_core[42] sky130_fd_sc_hd__buf_8
XFILLER_40_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput794 _549_/X vssd vssd vccd vccd la_oenb_core[52] sky130_fd_sc_hd__buf_8
XFILLER_5_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_322_ _322_/A _322_/B vssd vssd vccd vccd _322_/X sky130_fd_sc_hd__and2_4
XTAP_1478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_253_ _253_/A _253_/B vssd vssd vccd vccd _253_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_184_ _184_/A _184_/B vssd vssd vccd vccd _184_/X sky130_fd_sc_hd__and2_2
XFILLER_52_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1790 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_4480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_370 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_381 _470_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_392 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_gates\[27\] mprj_dat_i_user[27] _294_/X vssd vssd vccd vccd _141_/A sky130_fd_sc_hd__nand2_2
Xuser_to_mprj_in_gates\[14\] la_data_out_core[14] _177_/X vssd vssd vccd vccd _161_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_33_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3772 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[125\] la_data_out_core[125] _288_/X vssd vssd vccd vccd _108_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_9_1587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_842 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4488 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2409 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1708 _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1719 _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput580 _459_/X vssd vssd vccd vccd la_data_in_core[90] sky130_fd_sc_hd__buf_8
XFILLER_40_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput591 _147_/Y vssd vssd vccd vccd la_data_in_mprj[0] sky130_fd_sc_hd__buf_8
XFILLER_43_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_305_ _305_/A _305_/B vssd vssd vccd vccd _305_/X sky130_fd_sc_hd__and2_4
XFILLER_15_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_236_ _236_/A _236_/B vssd vssd vccd vccd _236_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_167_ _167_/A _167_/B vssd vssd vccd vccd _167_/X sky130_fd_sc_hd__and2_1
XFILLER_6_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_098_ _098_/A vssd vssd vccd vccd _098_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3440 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1058 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput308 la_oenb_mprj[28] vssd vssd vccd vccd _525_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_29_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput319 la_oenb_mprj[38] vssd vssd vccd vccd _535_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1018 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_021_ _021_/A vssd vssd vccd vccd _021_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2206 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2217 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2228 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2239 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1505 _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1516 _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1527 _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1538 _384_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1549 _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_219_ _219_/A _219_/B vssd vssd vccd vccd _219_/X sky130_fd_sc_hd__and2_2
XFILLER_32_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1990 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[81\] la_data_out_core[81] _244_/X vssd vssd vccd vccd _064_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_23_3720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4550 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2747 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput105 la_data_out_mprj[76] vssd vssd vccd vccd _445_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput116 la_data_out_mprj[86] vssd vssd vccd vccd _455_/C sky130_fd_sc_hd__buf_8
XFILLER_44_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput127 la_data_out_mprj[96] vssd vssd vccd vccd _465_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput138 la_iena_mprj[105] vssd vssd vccd vccd _268_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput149 la_iena_mprj[115] vssd vssd vccd vccd _278_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_570_ _570_/A _570_/B vssd vssd vccd vccd _570_/X sky130_fd_sc_hd__and2_4
XTAP_3958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_903 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_914 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_925 _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_936 _621_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_947 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_958 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_969 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_004_ _004_/A vssd vssd vccd vccd _004_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2003 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2014 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2025 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2036 _555_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2047 _348_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1302 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1313 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2058 _300_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2069 _074_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1324 _283_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1335 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1346 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2326 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1357 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1368 _294_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1379 _352_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2570 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2581 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2592 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1880 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1891 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_622_ _622_/A _622_/B vssd vssd vccd vccd _622_/X sky130_fd_sc_hd__and2_4
XTAP_4478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_700 _583_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_711 _591_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_553_ _553_/A _553_/B vssd vssd vccd vccd _553_/X sky130_fd_sc_hd__and2_4
XANTENNA_722 _594_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_733 _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_744 _595_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_755 _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_766 _598_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_484_ _612_/A _484_/B _484_/C vssd vssd vccd vccd _484_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_777 _603_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_788 _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_799 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1110 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1121 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1132 _189_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1143 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1154 _198_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1165 _205_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1176 _214_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1187 _221_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1198 _229_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[44\] la_data_out_core[44] _207_/X vssd vssd vccd vccd _027_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2572 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput910 _121_/Y vssd vssd vccd vccd mprj_dat_i_core[7] sky130_fd_sc_hd__buf_8
XFILLER_28_2012 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput921 _354_/X vssd vssd vccd vccd mprj_dat_o_user[17] sky130_fd_sc_hd__buf_8
Xoutput932 _364_/X vssd vssd vccd vccd mprj_dat_o_user[27] sky130_fd_sc_hd__buf_8
Xoutput943 _345_/X vssd vssd vccd vccd mprj_dat_o_user[8] sky130_fd_sc_hd__buf_8
XFILLER_47_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput954 output954/A vssd vssd vccd vccd user2_vdd_powergood sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[6\] la_data_out_core[6] _169_/X vssd vssd vccd vccd _153_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_25_3645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1960 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2250 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_605_ _605_/A _605_/B vssd vssd vccd vccd _605_/X sky130_fd_sc_hd__and2_4
XFILLER_45_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_530 _495_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_541 _496_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_536_ _536_/A _536_/B vssd vssd vccd vccd _536_/X sky130_fd_sc_hd__and2_4
XFILLER_19_3972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_552 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_563 _499_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_574 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_585 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_596 _510_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_467_ _595_/A _467_/B _467_/C vssd vssd vccd vccd _467_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_398_ _526_/A _398_/B _398_/C vssd vssd vccd vccd _398_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1270 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_4183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4036 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput740 _616_/X vssd vssd vccd vccd la_oenb_core[119] sky130_fd_sc_hd__buf_8
XFILLER_5_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput751 _510_/X vssd vssd vccd vccd la_oenb_core[13] sky130_fd_sc_hd__buf_8
XFILLER_47_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput762 _520_/X vssd vssd vccd vccd la_oenb_core[23] sky130_fd_sc_hd__buf_8
XFILLER_21_4018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput773 _530_/X vssd vssd vccd vccd la_oenb_core[33] sky130_fd_sc_hd__buf_8
XFILLER_9_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput784 _540_/X vssd vssd vccd vccd la_oenb_core[43] sky130_fd_sc_hd__buf_8
XFILLER_40_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput795 _550_/X vssd vssd vccd vccd la_oenb_core[53] sky130_fd_sc_hd__buf_8
XFILLER_5_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3271 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_321_ _321_/A _321_/B vssd vssd vccd vccd _321_/X sky130_fd_sc_hd__and2_4
XTAP_1457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_252_ _252_/A _252_/B vssd vssd vccd vccd _252_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_183_ _183_/A _183_/B vssd vssd vccd vccd _183_/X sky130_fd_sc_hd__and2_2
XFILLER_35_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_94 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_360 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_371 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_382 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_519_ _519_/A _519_/B vssd vssd vccd vccd _519_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_393 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[118\] la_data_out_core[118] _281_/X vssd vssd vccd vccd _101_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_3_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput570 _450_/X vssd vssd vccd vccd la_data_in_core[81] sky130_fd_sc_hd__buf_8
XFILLER_44_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1709 _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput581 _460_/X vssd vssd vccd vccd la_data_in_core[91] sky130_fd_sc_hd__buf_8
XFILLER_47_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput592 _083_/Y vssd vssd vccd vccd la_data_in_mprj[100] sky130_fd_sc_hd__buf_8
XFILLER_25_3283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_304_ _304_/A _304_/B vssd vssd vccd vccd _304_/X sky130_fd_sc_hd__and2_4
X_235_ _235_/A _235_/B vssd vssd vccd vccd _235_/X sky130_fd_sc_hd__and2_4
XFILLER_50_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_166_ _166_/A _166_/B vssd vssd vccd vccd _166_/X sky130_fd_sc_hd__and2_1
XFILLER_49_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1251 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_097_ _097_/A vssd vssd vccd vccd _097_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_190 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1020 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4271 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput309 la_oenb_mprj[29] vssd vssd vccd vccd _526_/A sky130_fd_sc_hd__buf_6
XFILLER_25_1100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_020_ _020_/A vssd vssd vccd vccd _020_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_4129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2207 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2218 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2229 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1506 _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1517 _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1528 _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1539 _384_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_218_ _218_/A _218_/B vssd vssd vccd vccd _218_/X sky130_fd_sc_hd__and2_2
XFILLER_45_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_149_ _149_/A vssd vssd vccd vccd _149_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_290 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[74\] la_data_out_core[74] _237_/X vssd vssd vccd vccd _057_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_3_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_4117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput106 la_data_out_mprj[77] vssd vssd vccd vccd _446_/C sky130_fd_sc_hd__buf_4
XFILLER_41_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput117 la_data_out_mprj[87] vssd vssd vccd vccd _456_/C sky130_fd_sc_hd__buf_8
XFILLER_48_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput128 la_data_out_mprj[97] vssd vssd vccd vccd _466_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput139 la_iena_mprj[106] vssd vssd vccd vccd _269_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2530 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_904 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_915 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_926 _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_937 _621_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_948 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_959 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_90 mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_003_ _003_/A vssd vssd vccd vccd _003_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2004 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2015 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2026 _304_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2037 _587_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2048 _349_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1303 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2059 output951/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1314 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1325 _283_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1336 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1347 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2338 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1358 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1369 _294_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1018 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2560 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2571 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2582 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2593 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1870 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1881 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1892 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[100\] la_data_out_core[100] _263_/X vssd vssd vccd vccd _083_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_39_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_621_ _621_/A _621_/B vssd vssd vccd vccd _621_/X sky130_fd_sc_hd__and2_4
XTAP_4468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_701 _583_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_712 _593_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_552_ _552_/A _552_/B vssd vssd vccd vccd _552_/X sky130_fd_sc_hd__and2_4
XTAP_3778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_723 _594_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_734 _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_745 _595_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_756 _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_767 _598_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_483_ _611_/A _483_/B _483_/C vssd vssd vccd vccd _483_/X sky130_fd_sc_hd__and3b_4
XFILLER_44_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_778 _603_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_789 _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_654 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1100 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1111 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1122 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1133 _190_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1144 _196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1155 _198_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1166 _206_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1177 _215_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1188 _221_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1199 _231_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_4201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[37\] la_data_out_core[37] _200_/X vssd vssd vccd vccd _020_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_53_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput900 _141_/Y vssd vssd vccd vccd mprj_dat_i_core[27] sky130_fd_sc_hd__buf_8
XFILLER_47_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput911 _122_/Y vssd vssd vccd vccd mprj_dat_i_core[8] sky130_fd_sc_hd__buf_8
XFILLER_28_2002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput922 _355_/X vssd vssd vccd vccd mprj_dat_o_user[18] sky130_fd_sc_hd__buf_8
Xoutput933 _365_/X vssd vssd vccd vccd mprj_dat_o_user[28] sky130_fd_sc_hd__buf_8
Xoutput944 _346_/X vssd vssd vccd vccd mprj_dat_o_user[9] sky130_fd_sc_hd__buf_8
XFILLER_8_2107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput955 _296_/X vssd vssd vccd vccd user_clock sky130_fd_sc_hd__buf_8
XFILLER_45_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4110 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2390 _335_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_4129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_604_ _604_/A _604_/B vssd vssd vccd vccd _604_/X sky130_fd_sc_hd__and2_4
XTAP_4298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1550 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_520 _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_531 _495_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_535_ _535_/A _535_/B vssd vssd vccd vccd _535_/X sky130_fd_sc_hd__and2_4
XFILLER_15_4549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_542 _497_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_553 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_564 _499_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_575 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_586 _315_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_597 _510_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_466_ _594_/A _466_/B _466_/C vssd vssd vccd vccd _466_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_4262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_397_ _525_/A _397_/B _397_/C vssd vssd vccd vccd _397_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1632 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4075 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput730 _507_/X vssd vssd vccd vccd la_oenb_core[10] sky130_fd_sc_hd__buf_8
XFILLER_25_3421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput741 _508_/X vssd vssd vccd vccd la_oenb_core[11] sky130_fd_sc_hd__buf_8
Xoutput752 _511_/X vssd vssd vccd vccd la_oenb_core[14] sky130_fd_sc_hd__buf_8
XFILLER_47_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput763 _521_/X vssd vssd vccd vccd la_oenb_core[24] sky130_fd_sc_hd__buf_8
Xoutput774 _531_/X vssd vssd vccd vccd la_oenb_core[34] sky130_fd_sc_hd__buf_8
XFILLER_25_4199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput785 _541_/X vssd vssd vccd vccd la_oenb_core[44] sky130_fd_sc_hd__buf_8
Xoutput796 _551_/X vssd vssd vccd vccd la_oenb_core[54] sky130_fd_sc_hd__buf_8
XFILLER_48_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_320_ _320_/A _320_/B vssd vssd vccd vccd _320_/X sky130_fd_sc_hd__and2_4
XFILLER_42_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_251_ _251_/A _251_/B vssd vssd vccd vccd _251_/X sky130_fd_sc_hd__and2_4
XFILLER_23_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2270 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_270 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_182_ _182_/A _182_/B vssd vssd vccd vccd _182_/X sky130_fd_sc_hd__and2_2
XFILLER_49_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_350 _310_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_361 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3634 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_518_ _518_/A _518_/B vssd vssd vccd vccd _518_/X sky130_fd_sc_hd__and2_4
XANTENNA_372 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_383 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_394 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_449_ _577_/A _449_/B _449_/C vssd vssd vccd vccd _449_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_4092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput560 _441_/X vssd vssd vccd vccd la_data_in_core[72] sky130_fd_sc_hd__buf_8
XFILLER_40_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput571 _451_/X vssd vssd vccd vccd la_data_in_core[82] sky130_fd_sc_hd__buf_8
XFILLER_43_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput582 _461_/X vssd vssd vccd vccd la_data_in_core[92] sky130_fd_sc_hd__buf_8
XFILLER_44_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput593 _084_/Y vssd vssd vccd vccd la_data_in_mprj[101] sky130_fd_sc_hd__buf_8
XFILLER_40_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_303_ _303_/A _303_/B vssd vssd vccd vccd _303_/X sky130_fd_sc_hd__and2_4
XTAP_1288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_590 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_94 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_234_ _234_/A _234_/B vssd vssd vccd vccd _234_/X sky130_fd_sc_hd__and2_4
XFILLER_7_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_165_ _165_/A _165_/B vssd vssd vccd vccd _165_/X sky130_fd_sc_hd__and2_1
XFILLER_6_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[2\] mprj_dat_i_user[2] _294_/X vssd vssd vccd vccd _116_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_096_ _096_/A vssd vssd vccd vccd _096_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3026 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3718 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_2908 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_180 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_191 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3464 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2054 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2076 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2208 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2219 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1507 _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1518 _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1529 _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3070 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_126 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3762 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_217_ _217_/A _217_/B vssd vssd vccd vccd _217_/X sky130_fd_sc_hd__and2_2
XFILLER_10_4095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_148_ _148_/A vssd vssd vccd vccd _148_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_13_1071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_079_ _079_/A vssd vssd vccd vccd _079_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[67\] la_data_out_core[67] _230_/X vssd vssd vccd vccd _050_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_22_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_847 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput107 la_data_out_mprj[78] vssd vssd vccd vccd _447_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput118 la_data_out_mprj[88] vssd vssd vccd vccd _457_/C sky130_fd_sc_hd__buf_8
XFILLER_41_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput129 la_data_out_mprj[98] vssd vssd vccd vccd _467_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2542 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2783 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_905 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_916 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_927 _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_938 _621_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_949 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_80 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_002_ _002_/A vssd vssd vccd vccd _002_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_91 mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2005 _302_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2016 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2027 _299_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2038 _588_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1304 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2049 _350_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1315 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1326 _284_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1337 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1348 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1359 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_4325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2550 _535_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2561 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2572 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2583 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2594 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1860 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1871 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1882 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1893 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_620_ _620_/A _620_/B vssd vssd vccd vccd _620_/X sky130_fd_sc_hd__and2_4
XTAP_4458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_702 _583_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_551_ _551_/A _551_/B vssd vssd vccd vccd _551_/X sky130_fd_sc_hd__and2_4
XTAP_3768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_713 _594_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_724 _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_735 _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_746 _595_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_482_ _610_/A _482_/B _482_/C vssd vssd vccd vccd _482_/X sky130_fd_sc_hd__and3b_4
XANTENNA_757 _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_768 _598_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_779 _603_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1101 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1112 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1123 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1134 _190_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1145 _196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1156 _198_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1167 _207_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_1178 _215_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1189 _333_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput460 user_irq_ena[0] vssd vssd vccd vccd _291_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput901 _142_/Y vssd vssd vccd vccd mprj_dat_i_core[28] sky130_fd_sc_hd__buf_8
Xoutput912 _123_/Y vssd vssd vccd vccd mprj_dat_i_core[9] sky130_fd_sc_hd__buf_8
Xoutput923 _356_/X vssd vssd vccd vccd mprj_dat_o_user[19] sky130_fd_sc_hd__buf_8
XFILLER_9_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput934 _366_/X vssd vssd vccd vccd mprj_dat_o_user[29] sky130_fd_sc_hd__buf_8
XFILLER_47_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput945 _301_/X vssd vssd vccd vccd mprj_sel_o_user[0] sky130_fd_sc_hd__buf_8
Xoutput956 _297_/X vssd vssd vccd vccd user_clock2 sky130_fd_sc_hd__buf_8
XFILLER_8_2119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2380 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2391 _271_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1690 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_603_ _603_/A _603_/B vssd vssd vccd vccd _603_/X sky130_fd_sc_hd__and2_4
XTAP_3532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_510 _490_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1562 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_521 _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_532 _495_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_534_ _534_/A _534_/B vssd vssd vccd vccd _534_/X sky130_fd_sc_hd__and2_4
XTAP_2842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_543 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_554 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_565 _499_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_576 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_465_ _593_/A _465_/B _465_/C vssd vssd vccd vccd _465_/X sky130_fd_sc_hd__and3b_4
XANTENNA_587 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_598 _510_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_396_ _524_/A _396_/B _396_/C vssd vssd vccd vccd _396_/X sky130_fd_sc_hd__and3b_4
XFILLER_43_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3923 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput290 la_oenb_mprj[127] vssd vssd vccd vccd _624_/A sky130_fd_sc_hd__buf_6
XFILLER_3_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput720 _597_/X vssd vssd vccd vccd la_oenb_core[100] sky130_fd_sc_hd__buf_8
XFILLER_47_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput731 _607_/X vssd vssd vccd vccd la_oenb_core[110] sky130_fd_sc_hd__buf_8
XFILLER_9_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput742 _617_/X vssd vssd vccd vccd la_oenb_core[120] sky130_fd_sc_hd__buf_8
Xoutput753 _512_/X vssd vssd vccd vccd la_oenb_core[15] sky130_fd_sc_hd__buf_8
XFILLER_43_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput764 _522_/X vssd vssd vccd vccd la_oenb_core[25] sky130_fd_sc_hd__buf_8
XFILLER_47_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput775 _532_/X vssd vssd vccd vccd la_oenb_core[35] sky130_fd_sc_hd__buf_8
XFILLER_5_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput786 _542_/X vssd vssd vccd vccd la_oenb_core[45] sky130_fd_sc_hd__buf_8
Xoutput797 _552_/X vssd vssd vccd vccd la_oenb_core[55] sky130_fd_sc_hd__buf_8
XFILLER_25_3477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_250_ _250_/A _250_/B vssd vssd vccd vccd _250_/X sky130_fd_sc_hd__and2_4
XFILLER_36_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2282 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_181_ _181_/A _181_/B vssd vssd vccd vccd _181_/X sky130_fd_sc_hd__and2_2
XFILLER_52_1450 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_irq_gates\[1\] user_irq_core[1] _292_/X vssd vssd vccd vccd _112_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_340 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_351 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_517_ _517_/A _517_/B vssd vssd vccd vccd _517_/X sky130_fd_sc_hd__and2_4
XTAP_2672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_362 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_373 _457_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_384 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_395 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1334 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_448_ _576_/A _448_/B _448_/C vssd vssd vccd vccd _448_/X sky130_fd_sc_hd__and3b_4
XTAP_1982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_379_ _507_/A _379_/B _379_/C vssd vssd vccd vccd _379_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[97\] la_data_out_core[97] _260_/X vssd vssd vccd vccd _080_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_6_3825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3352 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_4561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_856 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1618 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput550 _432_/X vssd vssd vccd vccd la_data_in_core[63] sky130_fd_sc_hd__buf_8
Xoutput561 _442_/X vssd vssd vccd vccd la_data_in_core[73] sky130_fd_sc_hd__buf_8
Xoutput572 _452_/X vssd vssd vccd vccd la_data_in_core[83] sky130_fd_sc_hd__buf_8
XFILLER_47_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput583 _462_/X vssd vssd vccd vccd la_data_in_core[93] sky130_fd_sc_hd__buf_8
Xoutput594 _085_/Y vssd vssd vccd vccd la_data_in_mprj[102] sky130_fd_sc_hd__buf_8
XFILLER_5_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_319 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1819 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_302_ _302_/A _302_/B vssd vssd vccd vccd _302_/X sky130_fd_sc_hd__and2_4
XFILLER_51_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3988 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_233_ _233_/A _233_/B vssd vssd vccd vccd _233_/X sky130_fd_sc_hd__and2_2
XFILLER_50_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_230 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_164_ _164_/A _164_/B vssd vssd vccd vccd _164_/X sky130_fd_sc_hd__and2_1
XFILLER_10_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_095_ _095_/A vssd vssd vccd vccd _095_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_4384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3672 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_170 mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_181 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_192 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[12\] la_data_out_core[12] _175_/X vssd vssd vccd vccd _159_/A
+ sky130_fd_sc_hd__nand2_4
Xuser_wb_dat_gates\[25\] mprj_dat_i_user[25] _294_/X vssd vssd vccd vccd _139_/A sky130_fd_sc_hd__nand2_2
XFILLER_50_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[123\] la_data_out_core[123] _286_/X vssd vssd vccd vccd _106_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_29_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2209 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1508 _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1519 _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3616 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_216_ _216_/A _216_/B vssd vssd vccd vccd _216_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4074 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_147_ _147_/A vssd vssd vccd vccd _147_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1083 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_078_ _078_/A vssd vssd vccd vccd _078_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3739 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput108 la_data_out_mprj[79] vssd vssd vccd vccd _448_/C sky130_fd_sc_hd__buf_4
XFILLER_44_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput119 la_data_out_mprj[89] vssd vssd vccd vccd _458_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1026 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2795 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_906 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_917 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_928 _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_939 _621_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_70 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_81 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_001_ _001_/A vssd vssd vccd vccd _001_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_92 mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2006 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2017 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2028 _300_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2039 _315_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1305 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1316 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1327 _284_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1338 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1349 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2540 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2551 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2562 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2573 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2584 _362_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1850 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2595 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1861 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1872 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_1883 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1894 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput90 la_data_out_mprj[62] vssd vssd vccd vccd _431_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2467 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_550_ _550_/A _550_/B vssd vssd vccd vccd _550_/X sky130_fd_sc_hd__and2_4
XTAP_3758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_703 _583_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_714 _594_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_725 _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_736 _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_481_ _609_/A _481_/B _481_/C vssd vssd vccd vccd _481_/X sky130_fd_sc_hd__and3b_4
XFILLER_16_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_747 _595_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_4461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_758 _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_769 _598_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1102 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1113 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1124 _185_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4438 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1135 _191_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1146 _196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1157 _198_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1168 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1179 _215_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput450 mprj_dat_o_core[7] vssd vssd vccd vccd _344_/B sky130_fd_sc_hd__buf_8
Xinput461 user_irq_ena[1] vssd vssd vccd vccd _292_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput902 _143_/Y vssd vssd vccd vccd mprj_dat_i_core[29] sky130_fd_sc_hd__buf_8
Xoutput913 _337_/X vssd vssd vccd vccd mprj_dat_o_user[0] sky130_fd_sc_hd__buf_8
Xoutput924 _338_/X vssd vssd vccd vccd mprj_dat_o_user[1] sky130_fd_sc_hd__buf_8
Xoutput935 _339_/X vssd vssd vccd vccd mprj_dat_o_user[2] sky130_fd_sc_hd__buf_8
XFILLER_9_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput946 _302_/X vssd vssd vccd vccd mprj_sel_o_user[1] sky130_fd_sc_hd__buf_8
Xoutput957 _111_/Y vssd vssd vccd vccd user_irq[0] sky130_fd_sc_hd__buf_8
XFILLER_3_4101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2370 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2381 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2392 _271_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1680 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1691 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_236 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_346 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_602_ _602_/A _602_/B vssd vssd vccd vccd _602_/X sky130_fd_sc_hd__and2_4
XTAP_4278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_500 _488_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_511 _490_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_533_ _533_/A _533_/B vssd vssd vccd vccd _533_/X sky130_fd_sc_hd__and2_4
XANTENNA_522 _492_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1574 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_533 _495_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_544 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_555 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_566 _499_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_464_ _592_/A _464_/B _464_/C vssd vssd vccd vccd _464_/X sky130_fd_sc_hd__and3b_4
XANTENNA_577 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_588 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_599 _510_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_395_ _523_/A _395_/B _395_/C vssd vssd vccd vccd _395_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput280 la_oenb_mprj[118] vssd vssd vccd vccd _615_/A sky130_fd_sc_hd__buf_6
XFILLER_0_2927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput291 la_oenb_mprj[12] vssd vssd vccd vccd _509_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[42\] la_data_out_core[42] _205_/X vssd vssd vccd vccd _025_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_3441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput710 _075_/Y vssd vssd vccd vccd la_data_in_mprj[92] sky130_fd_sc_hd__buf_8
Xoutput721 _598_/X vssd vssd vccd vccd la_oenb_core[101] sky130_fd_sc_hd__buf_8
Xoutput732 _608_/X vssd vssd vccd vccd la_oenb_core[111] sky130_fd_sc_hd__buf_8
XFILLER_47_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput743 _618_/X vssd vssd vccd vccd la_oenb_core[121] sky130_fd_sc_hd__buf_8
XFILLER_9_3664 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput754 _513_/X vssd vssd vccd vccd la_oenb_core[16] sky130_fd_sc_hd__buf_8
Xoutput765 _523_/X vssd vssd vccd vccd la_oenb_core[26] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[4\] la_data_out_core[4] _167_/X vssd vssd vccd vccd _151_/A
+ sky130_fd_sc_hd__nand2_1
Xoutput776 _533_/X vssd vssd vccd vccd la_oenb_core[36] sky130_fd_sc_hd__buf_8
XFILLER_28_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput787 _543_/X vssd vssd vccd vccd la_oenb_core[46] sky130_fd_sc_hd__buf_8
Xoutput798 _553_/X vssd vssd vccd vccd la_oenb_core[56] sky130_fd_sc_hd__buf_8
XFILLER_42_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_180_ _180_/A _180_/B vssd vssd vccd vccd _180_/X sky130_fd_sc_hd__and2_1
XFILLER_17_2294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_330 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_341 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_516_ _516_/A _516_/B vssd vssd vccd vccd _516_/X sky130_fd_sc_hd__and2_4
XANTENNA_352 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_363 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_374 _457_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_385 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_396 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_447_ _575_/A _447_/B _447_/C vssd vssd vccd vccd _447_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_250 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1346 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_378_ _506_/A _378_/B _378_/C vssd vssd vccd vccd _378_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3743 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1030 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput540 _423_/X vssd vssd vccd vccd la_data_in_core[54] sky130_fd_sc_hd__buf_8
XFILLER_47_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput551 _433_/X vssd vssd vccd vccd la_data_in_core[64] sky130_fd_sc_hd__buf_8
XFILLER_9_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput562 _443_/X vssd vssd vccd vccd la_data_in_core[74] sky130_fd_sc_hd__buf_8
XFILLER_5_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput573 _453_/X vssd vssd vccd vccd la_data_in_core[84] sky130_fd_sc_hd__buf_8
XFILLER_43_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput584 _463_/X vssd vssd vccd vccd la_data_in_core[94] sky130_fd_sc_hd__buf_8
Xoutput595 _086_/Y vssd vssd vccd vccd la_data_in_mprj[103] sky130_fd_sc_hd__buf_8
XFILLER_21_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_301_ _301_/A _301_/B vssd vssd vccd vccd _301_/X sky130_fd_sc_hd__and2_4
XTAP_1268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_232_ _232_/A _232_/B vssd vssd vccd vccd _232_/X sky130_fd_sc_hd__and2_2
XFILLER_24_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_163_ _163_/A vssd vssd vccd vccd _163_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_094_ _094_/A vssd vssd vccd vccd _094_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_4396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_171 mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_182 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_193 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[18\] mprj_dat_i_user[18] _294_/X vssd vssd vccd vccd _132_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3150 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[116\] la_data_out_core[116] _279_/X vssd vssd vccd vccd _099_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_42_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_879 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1509 _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3166 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_96 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_4020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_215_ _215_/A _215_/B vssd vssd vccd vccd _215_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_146_ _146_/A vssd vssd vccd vccd _146_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_077_ _077_/A vssd vssd vccd vccd _077_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput109 la_data_out_mprj[7] vssd vssd vccd vccd _376_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_6_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1038 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_907 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_918 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_929 _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_319 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_60 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_000_ _000_/A vssd vssd vccd vccd _000_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_71 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_82 mprj_dat_i_user[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_93 mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2007 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2018 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2029 _300_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1306 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1317 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1328 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1339 _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3739 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_129_ _129_/A vssd vssd vccd vccd _129_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2530 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2541 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3690 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2552 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2563 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2574 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1840 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[72\] la_data_out_core[72] _235_/X vssd vssd vccd vccd _055_/A
+ sky130_fd_sc_hd__nand2_4
XANTENNA_2585 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1851 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2596 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1862 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1873 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1884 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1895 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput80 la_data_out_mprj[53] vssd vssd vccd vccd _422_/C sky130_fd_sc_hd__buf_4
XFILLER_28_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput91 la_data_out_mprj[63] vssd vssd vccd vccd _432_/C sky130_fd_sc_hd__buf_4
XFILLER_43_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_704 _583_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_715 _594_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_726 _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_480_ _608_/A _480_/B _480_/C vssd vssd vccd vccd _480_/X sky130_fd_sc_hd__and3b_4
XANTENNA_737 _595_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_748 _596_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_759 _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1103 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1114 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1125 _185_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1136 _191_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1147 _196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1158 _199_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1169 _210_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput440 mprj_dat_o_core[27] vssd vssd vccd vccd _364_/B sky130_fd_sc_hd__buf_8
XFILLER_23_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput451 mprj_dat_o_core[8] vssd vssd vccd vccd _345_/B sky130_fd_sc_hd__buf_8
Xinput462 user_irq_ena[2] vssd vssd vccd vccd _293_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput903 _116_/Y vssd vssd vccd vccd mprj_dat_i_core[2] sky130_fd_sc_hd__buf_8
XFILLER_7_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput914 _347_/X vssd vssd vccd vccd mprj_dat_o_user[10] sky130_fd_sc_hd__buf_8
Xoutput925 _357_/X vssd vssd vccd vccd mprj_dat_o_user[20] sky130_fd_sc_hd__buf_8
XFILLER_47_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput936 _367_/X vssd vssd vccd vccd mprj_dat_o_user[30] sky130_fd_sc_hd__buf_8
XFILLER_25_3627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput947 _303_/X vssd vssd vccd vccd mprj_sel_o_user[2] sky130_fd_sc_hd__buf_8
Xoutput958 _112_/Y vssd vssd vccd vccd user_irq[1] sky130_fd_sc_hd__buf_8
XFILLER_23_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2360 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2371 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2382 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2393 _271_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1670 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1681 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1692 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2498 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1964 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_601_ _601_/A _601_/B vssd vssd vccd vccd _601_/X sky130_fd_sc_hd__and2_4
XTAP_3512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_501 _490_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_532_ _532_/A _532_/B vssd vssd vccd vccd _532_/X sky130_fd_sc_hd__and2_4
XANTENNA_512 _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_523 _493_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_534 _496_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_545 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_556 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_463_ _591_/A _463_/B _463_/C vssd vssd vccd vccd _463_/X sky130_fd_sc_hd__and3b_4
XANTENNA_567 _499_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_578 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_589 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_394_ _522_/A _394_/B _394_/C vssd vssd vccd vccd _394_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput270 la_oenb_mprj[109] vssd vssd vccd vccd _606_/A sky130_fd_sc_hd__buf_6
Xinput281 la_oenb_mprj[119] vssd vssd vccd vccd _616_/A sky130_fd_sc_hd__buf_6
XFILLER_7_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput292 la_oenb_mprj[13] vssd vssd vccd vccd _510_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[35\] la_data_out_core[35] _198_/X vssd vssd vccd vccd _018_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_17_1027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput700 _066_/Y vssd vssd vccd vccd la_data_in_mprj[83] sky130_fd_sc_hd__buf_8
XFILLER_9_4366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput711 _076_/Y vssd vssd vccd vccd la_data_in_mprj[93] sky130_fd_sc_hd__buf_8
XFILLER_9_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput722 _599_/X vssd vssd vccd vccd la_oenb_core[102] sky130_fd_sc_hd__buf_8
Xoutput733 _609_/X vssd vssd vccd vccd la_oenb_core[112] sky130_fd_sc_hd__buf_8
Xoutput744 _619_/X vssd vssd vccd vccd la_oenb_core[122] sky130_fd_sc_hd__buf_8
XFILLER_25_3435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput755 _514_/X vssd vssd vccd vccd la_oenb_core[17] sky130_fd_sc_hd__buf_8
XFILLER_47_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3676 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput766 _524_/X vssd vssd vccd vccd la_oenb_core[27] sky130_fd_sc_hd__buf_8
Xoutput777 _534_/X vssd vssd vccd vccd la_oenb_core[37] sky130_fd_sc_hd__buf_8
XFILLER_5_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput788 _544_/X vssd vssd vccd vccd la_oenb_core[47] sky130_fd_sc_hd__buf_8
XFILLER_25_2723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput799 _554_/X vssd vssd vccd vccd la_oenb_core[57] sky130_fd_sc_hd__buf_8
XFILLER_28_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2190 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_98 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_320 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_331 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_515_ _515_/A _515_/B vssd vssd vccd vccd _515_/X sky130_fd_sc_hd__and2_4
XANTENNA_342 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_353 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_364 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_375 _457_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_386 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_397 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_446_ _574_/A _446_/B _446_/C vssd vssd vccd vccd _446_/X sky130_fd_sc_hd__and3b_4
XTAP_1962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_377_ _505_/A _377_/B _377_/C vssd vssd vccd vccd _377_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_3372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3711 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1075 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2807 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput530 _414_/X vssd vssd vccd vccd la_data_in_core[45] sky130_fd_sc_hd__buf_8
XFILLER_9_3451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput541 _424_/X vssd vssd vccd vccd la_data_in_core[55] sky130_fd_sc_hd__buf_8
Xoutput552 _434_/X vssd vssd vccd vccd la_data_in_core[65] sky130_fd_sc_hd__buf_8
Xoutput563 _444_/X vssd vssd vccd vccd la_data_in_core[75] sky130_fd_sc_hd__buf_8
XFILLER_47_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput574 _454_/X vssd vssd vccd vccd la_data_in_core[85] sky130_fd_sc_hd__buf_8
Xoutput585 _464_/X vssd vssd vccd vccd la_data_in_core[95] sky130_fd_sc_hd__buf_8
Xoutput596 _087_/Y vssd vssd vccd vccd la_data_in_mprj[104] sky130_fd_sc_hd__buf_8
XFILLER_5_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_300_ _300_/A _300_/B vssd vssd vccd vccd _300_/X sky130_fd_sc_hd__and2_4
XFILLER_42_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_231_ _231_/A _231_/B vssd vssd vccd vccd _231_/X sky130_fd_sc_hd__and2_2
XFILLER_32_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_162_ _162_/A vssd vssd vccd vccd _162_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_093_ _093_/A vssd vssd vccd vccd _093_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3746 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_150 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_161 mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4168 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_172 mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_183 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_194 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_429_ _557_/A _429_/B _429_/C vssd vssd vccd vccd _429_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput1 caravel_clk vssd vssd vccd vccd _296_/B sky130_fd_sc_hd__buf_8
XFILLER_37_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[109\] la_data_out_core[109] _272_/X vssd vssd vccd vccd _092_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_0_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3178 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4319 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_214_ _214_/A _214_/B vssd vssd vccd vccd _214_/X sky130_fd_sc_hd__and2_2
XFILLER_7_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_145_ _145_/A vssd vssd vccd vccd _145_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[0\] mprj_dat_i_user[0] _294_/X vssd vssd vccd vccd _114_/A sky130_fd_sc_hd__nand2_1
XFILLER_49_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_076_ _076_/A vssd vssd vccd vccd _076_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[30\] mprj_dat_i_user[30] _294_/X vssd vssd vccd vccd _144_/A sky130_fd_sc_hd__nand2_2
XFILLER_21_327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_908 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_919 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_50 mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_61 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_72 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_83 mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_94 mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2008 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2019 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1307 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1318 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1329 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3830 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_128_ _128_/A vssd vssd vccd vccd _128_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_059_ _059_/A vssd vssd vccd vccd _059_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2520 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2531 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2542 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2553 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2564 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1830 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2575 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2586 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1841 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1852 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2597 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1863 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1874 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1885 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[65\] la_data_out_core[65] _228_/X vssd vssd vccd vccd _048_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_40_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1896 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput70 la_data_out_mprj[44] vssd vssd vccd vccd _413_/C sky130_fd_sc_hd__clkbuf_4
Xinput81 la_data_out_mprj[54] vssd vssd vccd vccd _423_/C sky130_fd_sc_hd__clkbuf_4
Xinput92 la_data_out_mprj[64] vssd vssd vccd vccd _433_/C sky130_fd_sc_hd__buf_4
XFILLER_45_4481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1746 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_705 _583_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_716 _594_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_727 _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_738 _595_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_749 _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_4474 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_146 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1104 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1115 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1126 _185_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1137 _192_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1148 _196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3728 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1159 _199_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput430 mprj_dat_o_core[18] vssd vssd vccd vccd _355_/B sky130_fd_sc_hd__buf_8
XFILLER_2_4372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput441 mprj_dat_o_core[28] vssd vssd vccd vccd _365_/B sky130_fd_sc_hd__buf_6
XFILLER_48_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput452 mprj_dat_o_core[9] vssd vssd vccd vccd _346_/B sky130_fd_sc_hd__buf_8
XFILLER_5_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4410 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput904 _144_/Y vssd vssd vccd vccd mprj_dat_i_core[30] sky130_fd_sc_hd__buf_8
XFILLER_28_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput915 _348_/X vssd vssd vccd vccd mprj_dat_o_user[11] sky130_fd_sc_hd__buf_8
XFILLER_28_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput926 _358_/X vssd vssd vccd vccd mprj_dat_o_user[21] sky130_fd_sc_hd__buf_8
Xoutput937 _368_/X vssd vssd vccd vccd mprj_dat_o_user[31] sky130_fd_sc_hd__buf_8
XFILLER_47_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput948 _304_/X vssd vssd vccd vccd mprj_sel_o_user[3] sky130_fd_sc_hd__buf_8
XFILLER_25_3639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput959 _113_/Y vssd vssd vccd vccd user_irq[2] sky130_fd_sc_hd__buf_8
XFILLER_7_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2350 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2361 _308_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2372 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2383 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2394 _271_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1660 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1671 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1682 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1693 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1988 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_600_ _600_/A _600_/B vssd vssd vccd vccd _600_/X sky130_fd_sc_hd__and2_4
XTAP_3513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_531_ _531_/A _531_/B vssd vssd vccd vccd _531_/X sky130_fd_sc_hd__and2_4
XTAP_2812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_502 _490_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_513 _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_524 _493_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_535 _496_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_546 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_462_ _590_/A _462_/B _462_/C vssd vssd vccd vccd _462_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_557 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4271 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_568 _500_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_579 _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_393_ _521_/A _393_/B _393_/C vssd vssd vccd vccd _393_/X sky130_fd_sc_hd__and3b_4
XFILLER_41_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput260 la_oenb_mprj[0] vssd vssd vccd vccd _497_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput271 la_oenb_mprj[10] vssd vssd vccd vccd _507_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput282 la_oenb_mprj[11] vssd vssd vccd vccd _508_/A sky130_fd_sc_hd__clkbuf_4
Xinput293 la_oenb_mprj[14] vssd vssd vccd vccd _511_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[28\] la_data_out_core[28] _191_/X vssd vssd vccd vccd _011_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput701 _067_/Y vssd vssd vccd vccd la_data_in_mprj[84] sky130_fd_sc_hd__buf_8
Xoutput712 _077_/Y vssd vssd vccd vccd la_data_in_mprj[94] sky130_fd_sc_hd__buf_8
XFILLER_25_3403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput723 _600_/X vssd vssd vccd vccd la_oenb_core[103] sky130_fd_sc_hd__buf_8
Xoutput734 _610_/X vssd vssd vccd vccd la_oenb_core[113] sky130_fd_sc_hd__buf_8
XFILLER_29_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput745 _620_/X vssd vssd vccd vccd la_oenb_core[123] sky130_fd_sc_hd__buf_8
Xoutput756 _515_/X vssd vssd vccd vccd la_oenb_core[18] sky130_fd_sc_hd__buf_8
XFILLER_42_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput767 _525_/X vssd vssd vccd vccd la_oenb_core[28] sky130_fd_sc_hd__buf_8
XFILLER_25_3447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput778 _535_/X vssd vssd vccd vccd la_oenb_core[38] sky130_fd_sc_hd__buf_8
XFILLER_29_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput789 _545_/X vssd vssd vccd vccd la_oenb_core[48] sky130_fd_sc_hd__buf_8
XFILLER_25_2735 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2180 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2191 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1490 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_310 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_321 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_514_ _514_/A _514_/B vssd vssd vccd vccd _514_/X sky130_fd_sc_hd__and2_4
XANTENNA_332 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_343 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_354 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_365 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_376 _465_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_445_ _573_/A _445_/B _445_/C vssd vssd vccd vccd _445_/X sky130_fd_sc_hd__and3b_4
XANTENNA_387 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_398 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_376_ _504_/A _376_/B _376_/C vssd vssd vccd vccd _376_/X sky130_fd_sc_hd__and3b_4
XFILLER_9_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1488 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3344 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1098 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput520 _405_/X vssd vssd vccd vccd la_data_in_core[36] sky130_fd_sc_hd__buf_8
Xoutput531 _415_/X vssd vssd vccd vccd la_data_in_core[46] sky130_fd_sc_hd__buf_8
XFILLER_44_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2819 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput542 _425_/X vssd vssd vccd vccd la_data_in_core[56] sky130_fd_sc_hd__buf_8
Xoutput553 _435_/X vssd vssd vccd vccd la_data_in_core[66] sky130_fd_sc_hd__buf_8
XFILLER_43_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput564 _445_/X vssd vssd vccd vccd la_data_in_core[76] sky130_fd_sc_hd__buf_8
Xoutput575 _455_/X vssd vssd vccd vccd la_data_in_core[86] sky130_fd_sc_hd__buf_8
XFILLER_47_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput586 _465_/X vssd vssd vccd vccd la_data_in_core[96] sky130_fd_sc_hd__buf_8
XFILLER_8_1004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput597 _088_/Y vssd vssd vccd vccd la_data_in_mprj[105] sky130_fd_sc_hd__buf_8
XFILLER_5_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_230_ _230_/A _230_/B vssd vssd vccd vccd _230_/X sky130_fd_sc_hd__and2_4
XFILLER_14_3660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_161_ _161_/A vssd vssd vccd vccd _161_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_3524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_98 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_092_ _092_/A vssd vssd vccd vccd _092_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_43_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_140 mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_173 mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_195 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_428_ _556_/A _428_/B _428_/C vssd vssd vccd vccd _428_/X sky130_fd_sc_hd__and3b_4
XFILLER_41_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_359_ _359_/A _359_/B vssd vssd vccd vccd _359_/X sky130_fd_sc_hd__and2_4
XFILLER_13_3192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[95\] la_data_out_core[95] _258_/X vssd vssd vccd vccd _078_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_44_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput2 caravel_clk2 vssd vssd vccd vccd _297_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_20_3185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_213_ _213_/A _213_/B vssd vssd vccd vccd _213_/X sky130_fd_sc_hd__and2_2
XFILLER_32_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4066 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_144_ _144_/A vssd vssd vccd vccd _144_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_075_ _075_/A vssd vssd vccd vccd _075_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_27_4541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[10\] la_data_out_core[10] _173_/X vssd vssd vccd vccd _157_/A
+ sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_gates\[23\] mprj_dat_i_user[23] _294_/X vssd vssd vccd vccd _137_/A sky130_fd_sc_hd__nand2_2
XFILLER_50_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4134 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[121\] la_data_out_core[121] _284_/X vssd vssd vccd vccd _104_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_39_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_909 _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_40 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_51 mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_62 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_73 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_84 mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_95 mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2009 _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1308 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1319 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_354 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_127_ _127_/A vssd vssd vccd vccd _127_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_058_ _058_/A vssd vssd vccd vccd _058_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2510 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2521 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2532 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2543 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2554 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2565 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1820 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1831 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2576 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2587 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1842 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1853 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2598 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1864 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1875 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1886 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1897 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[58\] la_data_out_core[58] _221_/X vssd vssd vccd vccd _041_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_19_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput60 la_data_out_mprj[35] vssd vssd vccd vccd _404_/C sky130_fd_sc_hd__clkbuf_4
Xinput71 la_data_out_mprj[45] vssd vssd vccd vccd _414_/C sky130_fd_sc_hd__clkbuf_4
Xinput82 la_data_out_mprj[55] vssd vssd vccd vccd _424_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput93 la_data_out_mprj[65] vssd vssd vccd vccd _434_/C sky130_fd_sc_hd__buf_6
XFILLER_41_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_706 _583_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_717 _594_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_728 _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_739 _595_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_4453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_4404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3714 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_4555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1105 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1116 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1127 _185_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1138 _194_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1149 _196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput420 mprj_cyc_o_core vssd vssd vccd vccd _298_/B sky130_fd_sc_hd__buf_8
Xinput431 mprj_dat_o_core[19] vssd vssd vccd vccd _356_/B sky130_fd_sc_hd__buf_8
XFILLER_40_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput442 mprj_dat_o_core[29] vssd vssd vccd vccd _366_/B sky130_fd_sc_hd__buf_6
XFILLER_0_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput453 mprj_iena_wb vssd vssd vccd vccd _294_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_48_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput905 _145_/Y vssd vssd vccd vccd mprj_dat_i_core[31] sky130_fd_sc_hd__buf_8
XFILLER_49_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput916 _349_/X vssd vssd vccd vccd mprj_dat_o_user[12] sky130_fd_sc_hd__buf_8
XFILLER_29_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput927 _359_/X vssd vssd vccd vccd mprj_dat_o_user[22] sky130_fd_sc_hd__buf_8
XFILLER_28_2029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput938 _340_/X vssd vssd vccd vccd mprj_dat_o_user[3] sky130_fd_sc_hd__buf_8
Xoutput949 _299_/X vssd vssd vccd vccd mprj_stb_o_user sky130_fd_sc_hd__buf_8
XFILLER_45_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2340 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2351 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2362 _309_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2373 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2384 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1650 _588_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2395 _271_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1661 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1672 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1683 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1694 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_530_ _530_/A _530_/B vssd vssd vccd vccd _530_/X sky130_fd_sc_hd__and2_4
XTAP_3558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_503 _490_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_514 _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_525 _494_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_536 _496_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_461_ _589_/A _461_/B _461_/C vssd vssd vccd vccd _461_/X sky130_fd_sc_hd__and3b_4
XANTENNA_547 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_558 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_569 _501_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_392_ _520_/A _392_/B _392_/C vssd vssd vccd vccd _392_/X sky130_fd_sc_hd__and3b_4
XFILLER_52_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1298 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput250 la_iena_mprj[91] vssd vssd vccd vccd _254_/B sky130_fd_sc_hd__clkbuf_4
Xinput261 la_oenb_mprj[100] vssd vssd vccd vccd _597_/A sky130_fd_sc_hd__buf_6
Xinput272 la_oenb_mprj[110] vssd vssd vccd vccd _607_/A sky130_fd_sc_hd__buf_6
Xinput283 la_oenb_mprj[120] vssd vssd vccd vccd _617_/A sky130_fd_sc_hd__buf_6
XFILLER_23_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput294 la_oenb_mprj[15] vssd vssd vccd vccd _512_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3488 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput702 _068_/Y vssd vssd vccd vccd la_data_in_mprj[85] sky130_fd_sc_hd__buf_8
XFILLER_9_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput713 _078_/Y vssd vssd vccd vccd la_data_in_mprj[95] sky130_fd_sc_hd__buf_8
Xoutput724 _601_/X vssd vssd vccd vccd la_oenb_core[104] sky130_fd_sc_hd__buf_8
XFILLER_25_4149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput735 _611_/X vssd vssd vccd vccd la_oenb_core[114] sky130_fd_sc_hd__buf_8
XFILLER_25_3415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput746 _621_/X vssd vssd vccd vccd la_oenb_core[124] sky130_fd_sc_hd__buf_8
Xoutput757 _516_/X vssd vssd vccd vccd la_oenb_core[19] sky130_fd_sc_hd__buf_8
XFILLER_47_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput768 _526_/X vssd vssd vccd vccd la_oenb_core[29] sky130_fd_sc_hd__buf_8
Xoutput779 _536_/X vssd vssd vccd vccd la_oenb_core[39] sky130_fd_sc_hd__buf_8
XFILLER_25_3459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2170 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2181 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2192 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1480 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1491 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3880 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3706 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_300 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_311 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_513_ _513_/A _513_/B vssd vssd vccd vccd _513_/X sky130_fd_sc_hd__and2_4
XANTENNA_322 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_333 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_344 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_355 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_366 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_444_ _572_/A _444_/B _444_/C vssd vssd vccd vccd _444_/X sky130_fd_sc_hd__and3b_4
XANTENNA_377 _466_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_388 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_399 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_375_ _503_/A _375_/B _375_/C vssd vssd vccd vccd _375_/X sky130_fd_sc_hd__and3b_4
XTAP_1997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1467 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2644 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[40\] la_data_out_core[40] _203_/X vssd vssd vccd vccd _023_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_24_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput510 _396_/X vssd vssd vccd vccd la_data_in_core[27] sky130_fd_sc_hd__buf_8
XFILLER_9_4176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput521 _406_/X vssd vssd vccd vccd la_data_in_core[37] sky130_fd_sc_hd__buf_8
Xoutput532 _416_/X vssd vssd vccd vccd la_data_in_core[47] sky130_fd_sc_hd__buf_8
XFILLER_44_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput543 _426_/X vssd vssd vccd vccd la_data_in_core[57] sky130_fd_sc_hd__buf_8
XFILLER_25_3223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput554 _436_/X vssd vssd vccd vccd la_data_in_core[67] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[2\] la_data_out_core[2] _165_/X vssd vssd vccd vccd _149_/A
+ sky130_fd_sc_hd__nand2_2
Xoutput565 _446_/X vssd vssd vccd vccd la_data_in_core[77] sky130_fd_sc_hd__buf_8
XFILLER_5_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput576 _456_/X vssd vssd vccd vccd la_data_in_core[87] sky130_fd_sc_hd__buf_8
Xoutput587 _466_/X vssd vssd vccd vccd la_data_in_core[97] sky130_fd_sc_hd__buf_8
XFILLER_47_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput598 _089_/Y vssd vssd vccd vccd la_data_in_mprj[106] sky130_fd_sc_hd__buf_8
XFILLER_8_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_160_ _160_/A vssd vssd vccd vccd _160_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_3683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_091_ _091_/A vssd vssd vccd vccd _091_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_130 mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 mprj_dat_i_user[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_152 mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_163 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_185 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_196 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_427_ _555_/A _427_/B _427_/C vssd vssd vccd vccd _427_/X sky130_fd_sc_hd__and3b_4
XFILLER_18_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_358_ _358_/A _358_/B vssd vssd vccd vccd _358_/X sky130_fd_sc_hd__and2_4
XFILLER_50_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_289_ _289_/A _289_/B vssd vssd vccd vccd _289_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[88\] la_data_out_core[88] _251_/X vssd vssd vccd vccd _071_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_3587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput3 caravel_rstn vssd vssd vccd vccd input3/X sky130_fd_sc_hd__buf_8
XFILLER_20_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_598 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_4019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2352 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_212_ _212_/A _212_/B vssd vssd vccd vccd _212_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_143_ _143_/A vssd vssd vccd vccd _143_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_52_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2080 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_074_ _074_/A vssd vssd vccd vccd _074_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[16\] mprj_dat_i_user[16] _294_/X vssd vssd vccd vccd _130_/A sky130_fd_sc_hd__nand2_2
XFILLER_31_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_4124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_4146 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[114\] la_data_out_core[114] _277_/X vssd vssd vccd vccd _097_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_39_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_30 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_41 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_52 mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_63 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_74 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_85 mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_96 mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1309 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3876 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_126_ _126_/A vssd vssd vccd vccd _126_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_057_ _057_/A vssd vssd vccd vccd _057_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2500 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2511 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2522 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2533 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2544 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_1810 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2555 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3546 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2566 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1821 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1832 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2577 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2588 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1843 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1854 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2599 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1865 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1876 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1887 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1898 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1514 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput50 la_data_out_mprj[26] vssd vssd vccd vccd _395_/C sky130_fd_sc_hd__clkbuf_4
Xinput61 la_data_out_mprj[36] vssd vssd vccd vccd _405_/C sky130_fd_sc_hd__clkbuf_4
Xinput72 la_data_out_mprj[46] vssd vssd vccd vccd _415_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput83 la_data_out_mprj[56] vssd vssd vccd vccd _425_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput94 la_data_out_mprj[66] vssd vssd vccd vccd _435_/C sky130_fd_sc_hd__buf_6
XFILLER_28_3457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_707 _584_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_718 _594_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_4432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_729 _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3726 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1106 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1117 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1128 _186_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1139 _194_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput410 mprj_adr_o_core[2] vssd vssd vccd vccd _307_/B sky130_fd_sc_hd__buf_8
XFILLER_20_3719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput421 mprj_dat_o_core[0] vssd vssd vccd vccd _337_/B sky130_fd_sc_hd__buf_8
XFILLER_7_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput432 mprj_dat_o_core[1] vssd vssd vccd vccd _338_/B sky130_fd_sc_hd__buf_8
XFILLER_0_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput443 mprj_dat_o_core[2] vssd vssd vccd vccd _339_/B sky130_fd_sc_hd__buf_8
XFILLER_40_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput454 mprj_sel_o_core[0] vssd vssd vccd vccd _301_/B sky130_fd_sc_hd__buf_8
XFILLER_5_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3695 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3236 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_109_ _109_/A vssd vssd vccd vccd _109_/Y sky130_fd_sc_hd__clkinv_2
Xoutput906 _117_/Y vssd vssd vccd vccd mprj_dat_i_core[3] sky130_fd_sc_hd__buf_8
Xoutput917 _350_/X vssd vssd vccd vccd mprj_dat_o_user[13] sky130_fd_sc_hd__buf_8
XFILLER_45_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput928 _360_/X vssd vssd vccd vccd mprj_dat_o_user[23] sky130_fd_sc_hd__buf_8
XFILLER_7_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput939 _341_/X vssd vssd vccd vccd mprj_dat_o_user[4] sky130_fd_sc_hd__buf_8
XFILLER_7_4263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2330 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2341 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2352 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2363 _309_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2374 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2385 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1640 _571_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[70\] la_data_out_core[70] _233_/X vssd vssd vccd vccd _053_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1651 _594_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2396 _271_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1662 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1673 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1684 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1695 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_504 _490_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_515 _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_526 _495_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_460_ _588_/A _460_/B _460_/C vssd vssd vccd vccd _460_/X sky130_fd_sc_hd__and3b_4
XANTENNA_537 _496_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_548 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_559 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_391_ _519_/A _391_/B _391_/C vssd vssd vccd vccd _391_/X sky130_fd_sc_hd__and3b_4
XFILLER_17_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput240 la_iena_mprj[82] vssd vssd vccd vccd _245_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_20_3549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput251 la_iena_mprj[92] vssd vssd vccd vccd _255_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput262 la_oenb_mprj[101] vssd vssd vccd vccd _598_/A sky130_fd_sc_hd__clkbuf_8
Xinput273 la_oenb_mprj[111] vssd vssd vccd vccd _608_/A sky130_fd_sc_hd__buf_6
XFILLER_0_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput284 la_oenb_mprj[121] vssd vssd vccd vccd _618_/A sky130_fd_sc_hd__buf_6
Xinput295 la_oenb_mprj[16] vssd vssd vccd vccd _513_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_3401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_589_ _589_/A _589_/B vssd vssd vccd vccd _589_/X sky130_fd_sc_hd__and2_4
XFILLER_38_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_4336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput703 _069_/Y vssd vssd vccd vccd la_data_in_mprj[86] sky130_fd_sc_hd__buf_8
Xoutput714 _079_/Y vssd vssd vccd vccd la_data_in_mprj[96] sky130_fd_sc_hd__buf_8
Xoutput725 _602_/X vssd vssd vccd vccd la_oenb_core[105] sky130_fd_sc_hd__buf_8
XFILLER_47_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput736 _612_/X vssd vssd vccd vccd la_oenb_core[115] sky130_fd_sc_hd__buf_8
XFILLER_29_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput747 _622_/X vssd vssd vccd vccd la_oenb_core[125] sky130_fd_sc_hd__buf_8
Xoutput758 _498_/X vssd vssd vccd vccd la_oenb_core[1] sky130_fd_sc_hd__buf_8
XFILLER_42_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput769 _499_/X vssd vssd vccd vccd la_oenb_core[2] sky130_fd_sc_hd__buf_8
XFILLER_47_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2160 _280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2171 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2182 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2193 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1470 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1481 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1492 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_626 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_301 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_512_ _512_/A _512_/B vssd vssd vccd vccd _512_/X sky130_fd_sc_hd__and2_4
XFILLER_19_3732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_312 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_323 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_334 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_345 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_356 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_443_ _571_/A _443_/B _443_/C vssd vssd vccd vccd _443_/X sky130_fd_sc_hd__and3b_4
XTAP_2677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_367 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_378 _466_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_389 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_374_ _502_/A _374_/B _374_/C vssd vssd vccd vccd _374_/X sky130_fd_sc_hd__and3b_4
XTAP_1987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[33\] la_data_out_core[33] _196_/X vssd vssd vccd vccd _016_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_51_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_890 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput500 _387_/X vssd vssd vccd vccd la_data_in_core[18] sky130_fd_sc_hd__buf_8
Xoutput511 _397_/X vssd vssd vccd vccd la_data_in_core[28] sky130_fd_sc_hd__buf_8
Xoutput522 _407_/X vssd vssd vccd vccd la_data_in_core[38] sky130_fd_sc_hd__buf_8
XFILLER_9_4188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput533 _417_/X vssd vssd vccd vccd la_data_in_core[48] sky130_fd_sc_hd__buf_8
XFILLER_47_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput544 _427_/X vssd vssd vccd vccd la_data_in_core[58] sky130_fd_sc_hd__buf_8
Xoutput555 _437_/X vssd vssd vccd vccd la_data_in_core[68] sky130_fd_sc_hd__buf_8
XFILLER_25_3235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput566 _447_/X vssd vssd vccd vccd la_data_in_core[78] sky130_fd_sc_hd__buf_8
Xoutput577 _457_/X vssd vssd vccd vccd la_data_in_core[88] sky130_fd_sc_hd__buf_8
XFILLER_5_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput588 _467_/X vssd vssd vccd vccd la_data_in_core[98] sky130_fd_sc_hd__buf_8
Xoutput599 _090_/Y vssd vssd vccd vccd la_data_in_mprj[107] sky130_fd_sc_hd__buf_8
XFILLER_25_2556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4352 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_090_ _090_/A vssd vssd vccd vccd _090_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3830 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_4334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3738 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_858 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_120 mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_142 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_153 mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_164 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_175 mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_186 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_426_ _554_/A _426_/B _426_/C vssd vssd vccd vccd _426_/X sky130_fd_sc_hd__and3b_4
XFILLER_37_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_197 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_357_ _357_/A _357_/B vssd vssd vccd vccd _357_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_288_ _288_/A _288_/B vssd vssd vccd vccd _288_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2898 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput4 la_data_out_mprj[0] vssd vssd vccd vccd _369_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_20_2464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_89 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_211_ _211_/A _211_/B vssd vssd vccd vccd _211_/X sky130_fd_sc_hd__and2_1
XFILLER_49_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_142_ _142_/A vssd vssd vccd vccd _142_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_073_ _073_/A vssd vssd vccd vccd _073_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_2655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_4543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1998 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_409_ _537_/A _409_/B _409_/C vssd vssd vccd vccd _409_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4158 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[107\] la_data_out_core[107] _270_/X vssd vssd vccd vccd _090_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_53_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_20 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_31 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_42 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_53 mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_64 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_75 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_86 mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_97 mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3822 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1139 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_125_ _125_/A vssd vssd vccd vccd _125_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_056_ _056_/A vssd vssd vccd vccd _056_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_2485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2501 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2512 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2523 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2534 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2545 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1800 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1811 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2556 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1822 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2567 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1833 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3558 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2578 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2589 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1844 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1855 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1866 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1877 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1888 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1899 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput40 la_data_out_mprj[17] vssd vssd vccd vccd _386_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput51 la_data_out_mprj[27] vssd vssd vccd vccd _396_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput62 la_data_out_mprj[37] vssd vssd vccd vccd _406_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput73 la_data_out_mprj[47] vssd vssd vccd vccd _416_/C sky130_fd_sc_hd__buf_4
Xinput84 la_data_out_mprj[57] vssd vssd vccd vccd _426_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput95 la_data_out_mprj[67] vssd vssd vccd vccd _436_/C sky130_fd_sc_hd__buf_6
XFILLER_45_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1738 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_708 _323_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_719 _594_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3738 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1107 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1118 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1129 _186_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput400 mprj_adr_o_core[20] vssd vssd vccd vccd _325_/B sky130_fd_sc_hd__buf_8
Xinput411 mprj_adr_o_core[30] vssd vssd vccd vccd _335_/B sky130_fd_sc_hd__buf_8
XFILLER_40_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput422 mprj_dat_o_core[10] vssd vssd vccd vccd _347_/B sky130_fd_sc_hd__buf_8
Xinput433 mprj_dat_o_core[20] vssd vssd vccd vccd _357_/B sky130_fd_sc_hd__buf_8
XFILLER_7_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput444 mprj_dat_o_core[30] vssd vssd vccd vccd _367_/B sky130_fd_sc_hd__buf_6
Xinput455 mprj_sel_o_core[1] vssd vssd vccd vccd _302_/B sky130_fd_sc_hd__buf_8
XFILLER_22_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_488 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_108_ _108_/A vssd vssd vccd vccd _108_/Y sky130_fd_sc_hd__clkinv_2
Xoutput907 _118_/Y vssd vssd vccd vccd mprj_dat_i_core[4] sky130_fd_sc_hd__buf_8
XFILLER_49_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput918 _351_/X vssd vssd vccd vccd mprj_dat_o_user[14] sky130_fd_sc_hd__buf_8
Xoutput929 _361_/X vssd vssd vccd vccd mprj_dat_o_user[24] sky130_fd_sc_hd__buf_8
XFILLER_7_4253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_039_ _039_/A vssd vssd vccd vccd _039_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_2320 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2331 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2919 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2342 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2353 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2364 _309_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2375 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1630 _551_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1641 _571_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2386 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2397 _271_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1652 _595_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1663 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1674 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1685 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1696 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[63\] la_data_out_core[63] _226_/X vssd vssd vccd vccd _046_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_23_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_505 _490_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_516 _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_527 _495_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_538 _496_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_549 _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_390_ _518_/A _390_/B _390_/C vssd vssd vccd vccd _390_/X sky130_fd_sc_hd__and3b_4
XFILLER_52_4285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_296 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_992 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_4387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput230 la_iena_mprj[73] vssd vssd vccd vccd _236_/B sky130_fd_sc_hd__clkbuf_4
Xinput241 la_iena_mprj[83] vssd vssd vccd vccd _246_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput252 la_iena_mprj[93] vssd vssd vccd vccd _256_/B sky130_fd_sc_hd__clkbuf_4
Xinput263 la_oenb_mprj[102] vssd vssd vccd vccd _599_/A sky130_fd_sc_hd__buf_6
Xinput274 la_oenb_mprj[112] vssd vssd vccd vccd _609_/A sky130_fd_sc_hd__buf_6
XFILLER_49_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput285 la_oenb_mprj[122] vssd vssd vccd vccd _619_/A sky130_fd_sc_hd__buf_6
XFILLER_40_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput296 la_oenb_mprj[17] vssd vssd vccd vccd _514_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_588_ _588_/A _588_/B vssd vssd vccd vccd _588_/X sky130_fd_sc_hd__and2_4
XFILLER_34_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput704 _070_/Y vssd vssd vccd vccd la_data_in_mprj[87] sky130_fd_sc_hd__buf_8
XFILLER_29_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput715 _080_/Y vssd vssd vccd vccd la_data_in_mprj[97] sky130_fd_sc_hd__buf_8
Xoutput726 _603_/X vssd vssd vccd vccd la_oenb_core[106] sky130_fd_sc_hd__buf_8
XFILLER_42_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput737 _613_/X vssd vssd vccd vccd la_oenb_core[116] sky130_fd_sc_hd__buf_8
XFILLER_47_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput748 _623_/X vssd vssd vccd vccd la_oenb_core[126] sky130_fd_sc_hd__buf_8
XFILLER_7_4061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput759 _517_/X vssd vssd vccd vccd la_oenb_core[20] sky130_fd_sc_hd__buf_8
XFILLER_42_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2150 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2161 _280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2172 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2183 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2194 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1460 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1471 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1482 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1493 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1766 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_511_ _511_/A _511_/B vssd vssd vccd vccd _511_/X sky130_fd_sc_hd__and2_4
XANTENNA_302 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1354 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_313 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_324 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_4489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_335 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_346 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_442_ _570_/A _442_/B _442_/C vssd vssd vccd vccd _442_/X sky130_fd_sc_hd__and3b_4
XANTENNA_357 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_368 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_379 _468_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_373_ _501_/A _373_/B _373_/C vssd vssd vccd vccd _373_/X sky130_fd_sc_hd__and3b_4
XTAP_1988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[9\] mprj_dat_i_user[9] _294_/X vssd vssd vccd vccd _123_/A sky130_fd_sc_hd__nand2_2
XFILLER_26_4427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_880 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_891 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[26\] la_data_out_core[26] _189_/X vssd vssd vccd vccd _009_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_36_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput501 _388_/X vssd vssd vccd vccd la_data_in_core[19] sky130_fd_sc_hd__buf_8
Xoutput512 _398_/X vssd vssd vccd vccd la_data_in_core[29] sky130_fd_sc_hd__buf_8
XFILLER_29_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput523 _408_/X vssd vssd vccd vccd la_data_in_core[39] sky130_fd_sc_hd__buf_8
Xoutput534 _418_/X vssd vssd vccd vccd la_data_in_core[49] sky130_fd_sc_hd__buf_8
XFILLER_44_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput545 _428_/X vssd vssd vccd vccd la_data_in_core[59] sky130_fd_sc_hd__buf_8
XFILLER_47_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput556 _438_/X vssd vssd vccd vccd la_data_in_core[69] sky130_fd_sc_hd__buf_8
XFILLER_25_3247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput567 _448_/X vssd vssd vccd vccd la_data_in_core[79] sky130_fd_sc_hd__buf_8
XFILLER_5_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput578 _458_/X vssd vssd vccd vccd la_data_in_core[89] sky130_fd_sc_hd__buf_8
Xoutput589 _468_/X vssd vssd vccd vccd la_data_in_core[99] sky130_fd_sc_hd__buf_8
XFILLER_47_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1290 _279_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_402 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4346 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_4357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_110 mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_870 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_132 mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_165 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_187 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_425_ _553_/A _425_/B _425_/C vssd vssd vccd vccd _425_/X sky130_fd_sc_hd__and3b_4
XTAP_2497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 _396_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_356_ _356_/A _356_/B vssd vssd vccd vccd _356_/X sky130_fd_sc_hd__and2_4
XFILLER_35_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_287_ _287_/A _287_/B vssd vssd vccd vccd _287_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput5 la_data_out_mprj[100] vssd vssd vccd vccd _469_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_20_3177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3994 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3296 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3758 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_210_ _210_/A _210_/B vssd vssd vccd vccd _210_/X sky130_fd_sc_hd__and2_1
XFILLER_51_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_141_ _141_/A vssd vssd vccd vccd _141_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_13_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_072_ _072_/A vssd vssd vccd vccd _072_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_4515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4526 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_408_ _536_/A _408_/B _408_/C vssd vssd vccd vccd _408_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_339_ _339_/A _339_/B vssd vssd vccd vccd _339_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1708 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[93\] la_data_out_core[93] _256_/X vssd vssd vccd vccd _076_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_41_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_10 la_data_out_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_21 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_32 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_43 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_54 mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_65 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_76 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_87 mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_98 mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_124_ _124_/A vssd vssd vccd vccd _124_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_055_ _055_/A vssd vssd vccd vccd _055_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_49_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2502 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2513 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2524 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2535 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1801 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2546 _362_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2557 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1812 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2568 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1823 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1834 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2579 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1845 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1856 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1867 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1878 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1889 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3319 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3098 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[21\] mprj_dat_i_user[21] _294_/X vssd vssd vccd vccd _135_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput30 la_data_out_mprj[123] vssd vssd vccd vccd _492_/C sky130_fd_sc_hd__buf_4
XFILLER_50_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput41 la_data_out_mprj[18] vssd vssd vccd vccd _387_/C sky130_fd_sc_hd__clkbuf_4
Xinput52 la_data_out_mprj[28] vssd vssd vccd vccd _397_/C sky130_fd_sc_hd__clkbuf_4
Xinput63 la_data_out_mprj[38] vssd vssd vccd vccd _407_/C sky130_fd_sc_hd__clkbuf_4
Xinput74 la_data_out_mprj[48] vssd vssd vccd vccd _417_/C sky130_fd_sc_hd__clkbuf_4
Xinput85 la_data_out_mprj[58] vssd vssd vccd vccd _427_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_41_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput96 la_data_out_mprj[68] vssd vssd vccd vccd _437_/C sky130_fd_sc_hd__buf_6
XFILLER_45_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_709 _585_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3820 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3842 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1108 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1119 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput401 mprj_adr_o_core[21] vssd vssd vccd vccd _326_/B sky130_fd_sc_hd__buf_8
XFILLER_24_3879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput412 mprj_adr_o_core[31] vssd vssd vccd vccd _336_/B sky130_fd_sc_hd__buf_8
XFILLER_22_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput423 mprj_dat_o_core[11] vssd vssd vccd vccd _348_/B sky130_fd_sc_hd__buf_8
XFILLER_40_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput434 mprj_dat_o_core[21] vssd vssd vccd vccd _358_/B sky130_fd_sc_hd__buf_8
Xinput445 mprj_dat_o_core[31] vssd vssd vccd vccd _368_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput456 mprj_sel_o_core[2] vssd vssd vccd vccd _303_/B sky130_fd_sc_hd__buf_8
XFILLER_22_3592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_107_ _107_/A vssd vssd vccd vccd _107_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput908 _119_/Y vssd vssd vccd vccd mprj_dat_i_core[5] sky130_fd_sc_hd__buf_8
Xoutput919 _352_/X vssd vssd vccd vccd mprj_dat_o_user[15] sky130_fd_sc_hd__buf_8
XFILLER_45_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_038_ _038_/A vssd vssd vccd vccd _038_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_2310 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2321 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2332 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2343 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4068 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2354 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1620 _525_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2365 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2376 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1631 _554_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2387 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1642 _572_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1653 _596_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2398 _271_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1664 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1675 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1686 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1697 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[56\] la_data_out_core[56] _219_/X vssd vssd vccd vccd _039_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_35_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_506 _490_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_517 _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_528 _495_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_539 _496_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1880 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2931 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput220 la_iena_mprj[64] vssd vssd vccd vccd _227_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_1_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput231 la_iena_mprj[74] vssd vssd vccd vccd _237_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput242 la_iena_mprj[84] vssd vssd vccd vccd _247_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput253 la_iena_mprj[94] vssd vssd vccd vccd _257_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput264 la_oenb_mprj[103] vssd vssd vccd vccd _600_/A sky130_fd_sc_hd__buf_6
Xinput275 la_oenb_mprj[113] vssd vssd vccd vccd _610_/A sky130_fd_sc_hd__buf_6
Xinput286 la_oenb_mprj[123] vssd vssd vccd vccd _620_/A sky130_fd_sc_hd__buf_6
Xinput297 la_oenb_mprj[18] vssd vssd vccd vccd _515_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_587_ _587_/A _587_/B vssd vssd vccd vccd _587_/X sky130_fd_sc_hd__and2_4
XFILLER_32_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_463 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput705 _071_/Y vssd vssd vccd vccd la_data_in_mprj[88] sky130_fd_sc_hd__buf_8
Xoutput716 _081_/Y vssd vssd vccd vccd la_data_in_mprj[98] sky130_fd_sc_hd__buf_8
XFILLER_29_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput727 _604_/X vssd vssd vccd vccd la_oenb_core[107] sky130_fd_sc_hd__buf_8
Xoutput738 _614_/X vssd vssd vccd vccd la_oenb_core[117] sky130_fd_sc_hd__buf_8
XFILLER_42_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput749 _624_/X vssd vssd vccd vccd la_oenb_core[127] sky130_fd_sc_hd__buf_8
XFILLER_47_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2140 _260_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2151 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2162 _280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2173 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2184 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1450 _372_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2195 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1461 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1472 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1483 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1494 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4270 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1778 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_510_ _510_/A _510_/B vssd vssd vccd vccd _510_/X sky130_fd_sc_hd__and2_4
XFILLER_22_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_303 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_314 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_325 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_336 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_441_ _569_/A _441_/B _441_/C vssd vssd vccd vccd _441_/X sky130_fd_sc_hd__and3b_4
XTAP_1912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_347 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_358 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_369 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_372_ _500_/A _372_/B _372_/C vssd vssd vccd vccd _372_/X sky130_fd_sc_hd__and3b_4
XTAP_1967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_870 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_881 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_892 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[19\] la_data_out_core[19] _182_/X vssd vssd vccd vccd _002_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_32_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput502 _370_/X vssd vssd vccd vccd la_data_in_core[1] sky130_fd_sc_hd__buf_8
XFILLER_44_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput513 _371_/X vssd vssd vccd vccd la_data_in_core[2] sky130_fd_sc_hd__buf_8
XFILLER_48_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput524 _372_/X vssd vssd vccd vccd la_data_in_core[3] sky130_fd_sc_hd__buf_8
XFILLER_9_3445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput535 _373_/X vssd vssd vccd vccd la_data_in_core[4] sky130_fd_sc_hd__buf_8
Xoutput546 _374_/X vssd vssd vccd vccd la_data_in_core[5] sky130_fd_sc_hd__buf_8
XFILLER_44_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput557 _375_/X vssd vssd vccd vccd la_data_in_core[6] sky130_fd_sc_hd__buf_8
Xoutput568 _376_/X vssd vssd vccd vccd la_data_in_core[7] sky130_fd_sc_hd__buf_8
XFILLER_47_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput579 _377_/X vssd vssd vccd vccd la_data_in_core[8] sky130_fd_sc_hd__buf_8
XFILLER_5_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1280 _276_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1291 _279_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_2318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_598 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_458 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3602 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1130 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_122 mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_882 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_144 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_166 mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_424_ _552_/A _424_/B _424_/C vssd vssd vccd vccd _424_/X sky130_fd_sc_hd__and3b_4
XTAP_1742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 _398_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_355_ _355_/A _355_/B vssd vssd vccd vccd _355_/X sky130_fd_sc_hd__and2_4
XFILLER_50_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_598 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_286_ _286_/A _286_/B vssd vssd vccd vccd _286_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput6 la_data_out_mprj[101] vssd vssd vccd vccd _470_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[0\] la_data_out_core[0] _625_/X vssd vssd vccd vccd _147_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_9_2563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2344 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1862 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_134 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_140_ _140_/A vssd vssd vccd vccd _140_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_11_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_071_ _071_/A vssd vssd vccd vccd _071_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4538 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_407_ _535_/A _407_/B _407_/C vssd vssd vccd vccd _407_/X sky130_fd_sc_hd__and3b_4
XTAP_1572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_338_ _338_/A _338_/B vssd vssd vccd vccd _338_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_269_ _269_/A _269_/B vssd vssd vccd vccd _269_/X sky130_fd_sc_hd__and2_4
XFILLER_28_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[86\] la_data_out_core[86] _249_/X vssd vssd vccd vccd _069_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_39_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_11 la_data_out_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_22 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_33 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_44 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_55 mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_66 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_77 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_88 mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_99 mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4271 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_123_ _123_/A vssd vssd vccd vccd _123_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_054_ _054_/A vssd vssd vccd vccd _054_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_7_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2503 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2514 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2525 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2536 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1802 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2547 _309_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1813 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2558 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1824 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2569 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1835 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1846 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1857 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1868 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1879 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[14\] mprj_dat_i_user[14] _294_/X vssd vssd vccd vccd _128_/A sky130_fd_sc_hd__nand2_1
Xinput20 la_data_out_mprj[114] vssd vssd vccd vccd _483_/C sky130_fd_sc_hd__buf_6
XFILLER_28_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput31 la_data_out_mprj[124] vssd vssd vccd vccd _493_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_50_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput42 la_data_out_mprj[19] vssd vssd vccd vccd _388_/C sky130_fd_sc_hd__clkbuf_4
Xinput53 la_data_out_mprj[29] vssd vssd vccd vccd _398_/C sky130_fd_sc_hd__clkbuf_4
Xinput64 la_data_out_mprj[39] vssd vssd vccd vccd _408_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput75 la_data_out_mprj[49] vssd vssd vccd vccd _418_/C sky130_fd_sc_hd__buf_4
XFILLER_7_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput86 la_data_out_mprj[59] vssd vssd vccd vccd _428_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput97 la_data_out_mprj[69] vssd vssd vccd vccd _438_/C sky130_fd_sc_hd__buf_6
XFILLER_45_4486 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[112\] la_data_out_core[112] _275_/X vssd vssd vccd vccd _095_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_2_1718 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_402 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1464 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_630 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1109 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput402 mprj_adr_o_core[22] vssd vssd vccd vccd _327_/B sky130_fd_sc_hd__buf_8
Xinput413 mprj_adr_o_core[3] vssd vssd vccd vccd _308_/B sky130_fd_sc_hd__buf_8
Xinput424 mprj_dat_o_core[12] vssd vssd vccd vccd _349_/B sky130_fd_sc_hd__buf_8
Xinput435 mprj_dat_o_core[22] vssd vssd vccd vccd _359_/B sky130_fd_sc_hd__buf_8
Xinput446 mprj_dat_o_core[3] vssd vssd vccd vccd _340_/B sky130_fd_sc_hd__buf_8
XFILLER_0_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput457 mprj_sel_o_core[3] vssd vssd vccd vccd _304_/B sky130_fd_sc_hd__buf_8
XFILLER_21_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_106_ _106_/A vssd vssd vccd vccd _106_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput909 _120_/Y vssd vssd vccd vccd mprj_dat_i_core[6] sky130_fd_sc_hd__buf_8
X_037_ _037_/A vssd vssd vccd vccd _037_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2300 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2311 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2322 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2333 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2344 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1610 _614_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2355 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1621 _527_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2366 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1632 _555_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2377 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2388 _535_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1643 _574_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1654 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2399 _271_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1665 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1676 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1687 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1698 _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[49\] la_data_out_core[49] _212_/X vssd vssd vccd vccd _032_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_34_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_507 _490_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_518 _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_529 _495_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput210 la_iena_mprj[55] vssd vssd vccd vccd _218_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput221 la_iena_mprj[65] vssd vssd vccd vccd _228_/B sky130_fd_sc_hd__buf_4
XFILLER_24_3699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput232 la_iena_mprj[75] vssd vssd vccd vccd _238_/B sky130_fd_sc_hd__clkbuf_4
Xinput243 la_iena_mprj[85] vssd vssd vccd vccd _248_/B sky130_fd_sc_hd__clkbuf_4
Xinput254 la_iena_mprj[95] vssd vssd vccd vccd _258_/B sky130_fd_sc_hd__clkbuf_4
Xinput265 la_oenb_mprj[104] vssd vssd vccd vccd _601_/A sky130_fd_sc_hd__buf_6
XFILLER_48_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput276 la_oenb_mprj[114] vssd vssd vccd vccd _611_/A sky130_fd_sc_hd__buf_6
Xinput287 la_oenb_mprj[124] vssd vssd vccd vccd _621_/A sky130_fd_sc_hd__buf_6
XFILLER_18_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput298 la_oenb_mprj[19] vssd vssd vccd vccd _516_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_586_ _586_/A _586_/B vssd vssd vccd vccd _586_/X sky130_fd_sc_hd__and2_4
XFILLER_16_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput706 _072_/Y vssd vssd vccd vccd la_data_in_mprj[89] sky130_fd_sc_hd__buf_8
XFILLER_10_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput717 _082_/Y vssd vssd vccd vccd la_data_in_mprj[99] sky130_fd_sc_hd__buf_8
XFILLER_9_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput728 _605_/X vssd vssd vccd vccd la_oenb_core[108] sky130_fd_sc_hd__buf_8
Xoutput739 _615_/X vssd vssd vccd vccd la_oenb_core[118] sky130_fd_sc_hd__buf_8
XFILLER_42_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2707 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2130 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2141 _260_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2152 _278_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2163 _280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2174 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1440 _370_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2185 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1451 _372_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2196 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1462 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1473 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1484 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1495 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4458 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_304 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_315 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_326 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_337 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_440_ _568_/A _440_/B _440_/C vssd vssd vccd vccd _440_/X sky130_fd_sc_hd__and3b_4
XTAP_2658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_348 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_359 _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_371_ _499_/A _371_/B _371_/C vssd vssd vccd vccd _371_/X sky130_fd_sc_hd__and3b_4
XFILLER_18_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_4057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_860 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_871 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_569_ _569_/A _569_/B vssd vssd vccd vccd _569_/X sky130_fd_sc_hd__and2_4
XANTENNA_882 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_893 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput503 _389_/X vssd vssd vccd vccd la_data_in_core[20] sky130_fd_sc_hd__buf_8
Xoutput514 _399_/X vssd vssd vccd vccd la_data_in_core[30] sky130_fd_sc_hd__buf_8
XFILLER_44_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput525 _409_/X vssd vssd vccd vccd la_data_in_core[40] sky130_fd_sc_hd__buf_8
XFILLER_48_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput536 _419_/X vssd vssd vccd vccd la_data_in_core[50] sky130_fd_sc_hd__buf_8
XFILLER_47_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput547 _429_/X vssd vssd vccd vccd la_data_in_core[60] sky130_fd_sc_hd__buf_8
XFILLER_42_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput558 _439_/X vssd vssd vccd vccd la_data_in_core[70] sky130_fd_sc_hd__buf_8
Xoutput569 _449_/X vssd vssd vccd vccd la_data_in_core[80] sky130_fd_sc_hd__buf_8
XFILLER_47_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1270 _275_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1281 _276_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1292 _279_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3614 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3783 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_101 mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_123 mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1186 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_145 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_167 mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_423_ _551_/A _423_/B _423_/C vssd vssd vccd vccd _423_/X sky130_fd_sc_hd__and3b_4
XFILLER_14_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_178 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_189 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_354_ _354_/A _354_/B vssd vssd vccd vccd _354_/X sky130_fd_sc_hd__and2_4
XFILLER_35_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_285_ _285_/A _285_/B vssd vssd vccd vccd _285_/X sky130_fd_sc_hd__and2_4
XFILLER_26_4215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1307 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput7 la_data_out_mprj[102] vssd vssd vccd vccd _471_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[31\] la_data_out_core[31] _194_/X vssd vssd vccd vccd _014_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_690 _581_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_514 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1874 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_146 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4016 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_374 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_070_ _070_/A vssd vssd vccd vccd _070_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_49_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_234 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2063 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3516 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_406_ _534_/A _406_/B _406_/C vssd vssd vccd vccd _406_/X sky130_fd_sc_hd__and3b_4
XPHY_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_337_ _337_/A _337_/B vssd vssd vccd vccd _337_/X sky130_fd_sc_hd__and2_4
XFILLER_30_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_268_ _268_/A _268_/B vssd vssd vccd vccd _268_/X sky130_fd_sc_hd__and2_4
XFILLER_45_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_199_ _199_/A _199_/B vssd vssd vccd vccd _199_/X sky130_fd_sc_hd__and2_2
XFILLER_6_4117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2654 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2518 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[79\] la_data_out_core[79] _242_/X vssd vssd vccd vccd _062_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_12 la_data_out_core[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_23 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_34 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_45 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_56 mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_67 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_78 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_89 mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4236 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_122_ _122_/A vssd vssd vccd vccd _122_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1710 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_053_ _053_/A vssd vssd vccd vccd _053_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_27_4343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2504 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2515 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2526 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2537 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1803 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2548 _309_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2559 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1814 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1825 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1836 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1847 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1858 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1869 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput10 la_data_out_mprj[105] vssd vssd vccd vccd _474_/C sky130_fd_sc_hd__clkbuf_4
Xinput21 la_data_out_mprj[115] vssd vssd vccd vccd _484_/C sky130_fd_sc_hd__buf_4
XFILLER_28_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput32 la_data_out_mprj[125] vssd vssd vccd vccd _494_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_11_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput43 la_data_out_mprj[1] vssd vssd vccd vccd _370_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput54 la_data_out_mprj[2] vssd vssd vccd vccd _371_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput65 la_data_out_mprj[3] vssd vssd vccd vccd _372_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput76 la_data_out_mprj[4] vssd vssd vccd vccd _373_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput87 la_data_out_mprj[5] vssd vssd vccd vccd _374_/C sky130_fd_sc_hd__clkbuf_4
Xinput98 la_data_out_mprj[6] vssd vssd vccd vccd _375_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_45_4498 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[105\] la_data_out_core[105] _268_/X vssd vssd vccd vccd _088_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_53_712 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_414 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_4447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj2_logic_high_inst output953/A vccd2_uq0 vssd2_uq0 mprj2_logic_high
XFILLER_11_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput403 mprj_adr_o_core[23] vssd vssd vccd vccd _328_/B sky130_fd_sc_hd__buf_8
XFILLER_44_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput414 mprj_adr_o_core[4] vssd vssd vccd vccd _309_/B sky130_fd_sc_hd__buf_8
XFILLER_0_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput425 mprj_dat_o_core[13] vssd vssd vccd vccd _350_/B sky130_fd_sc_hd__buf_8
Xinput436 mprj_dat_o_core[23] vssd vssd vccd vccd _360_/B sky130_fd_sc_hd__buf_8
XFILLER_40_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput447 mprj_dat_o_core[4] vssd vssd vccd vccd _341_/B sky130_fd_sc_hd__buf_8
Xinput458 mprj_stb_o_core vssd vssd vccd vccd _299_/B sky130_fd_sc_hd__buf_8
XFILLER_2_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4022 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3310 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3398 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_105_ _105_/A vssd vssd vccd vccd _105_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_036_ _036_/A vssd vssd vccd vccd _036_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2301 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2312 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2323 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2334 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1600 _602_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2345 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2356 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1611 _615_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2367 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1622 _528_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2378 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1633 _560_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1644 _575_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2389 _330_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1655 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1666 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1677 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1688 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1699 _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_296 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_4560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high_inst _295_/B _395_/B _396_/B _397_/B _398_/B _399_/B _400_/B _401_/B
+ _402_/B _403_/B _404_/B _305_/A _405_/B _406_/B _407_/B _408_/B _409_/B _410_/B
+ _411_/B _412_/B _413_/B _414_/B _306_/A _415_/B _416_/B _417_/B _418_/B _419_/B
+ _420_/B _421_/B _422_/B _423_/B _424_/B _307_/A _425_/B _426_/B _427_/B _428_/B
+ _429_/B _430_/B _431_/B _432_/B _433_/B _434_/B _308_/A _435_/B _436_/B _437_/B
+ _438_/B _439_/B _440_/B _441_/B _442_/B _443_/B _444_/B _309_/A _445_/B _446_/B
+ _447_/B _448_/B _449_/B _450_/B _451_/B _452_/B _453_/B _454_/B _310_/A _455_/B
+ _456_/B _457_/B _458_/B _459_/B _460_/B _461_/B _462_/B _463_/B _464_/B _311_/A
+ _465_/B _466_/B _467_/B _468_/B _469_/B _470_/B _471_/B _472_/B _473_/B _474_/B
+ _312_/A _475_/B _476_/B _477_/B _478_/B _479_/B _480_/B _481_/B _482_/B _483_/B
+ _484_/B _313_/A _485_/B _486_/B _487_/B _488_/B _489_/B _490_/B _491_/B _492_/B
+ _493_/B _494_/B _314_/A _296_/A _495_/B _496_/B _497_/B _498_/B _499_/B _500_/B
+ _501_/B _502_/B _503_/B _504_/B _315_/A _505_/B _506_/B _507_/B _508_/B _509_/B
+ _510_/B _511_/B _512_/B _513_/B _514_/B _316_/A _515_/B _516_/B _517_/B _518_/B
+ _519_/B _520_/B _521_/B _522_/B _523_/B _524_/B _317_/A _525_/B _526_/B _527_/B
+ _528_/B _529_/B _530_/B _531_/B _532_/B _533_/B _534_/B _318_/A _535_/B _536_/B
+ _537_/B _538_/B _539_/B _540_/B _541_/B _542_/B _543_/B _544_/B _319_/A _545_/B
+ _546_/B _547_/B _548_/B _549_/B _550_/B _551_/B _552_/B _553_/B _554_/B _320_/A
+ _555_/B _556_/B _557_/B _558_/B _559_/B _560_/B _561_/B _562_/B _563_/B _564_/B
+ _321_/A _565_/B _566_/B _567_/B _568_/B _569_/B _570_/B _571_/B _572_/B _573_/B
+ _574_/B _322_/A _575_/B _576_/B _577_/B _578_/B _579_/B _580_/B _581_/B _582_/B
+ _583_/B _584_/B _323_/A _585_/B _586_/B _587_/B _588_/B _589_/B _590_/B _591_/B
+ _592_/B _593_/B _594_/B _324_/A _297_/A _595_/B _596_/B _597_/B _598_/B _599_/B
+ _600_/B _601_/B _602_/B _603_/B _604_/B _325_/A _605_/B _606_/B _607_/B _608_/B
+ _609_/B _610_/B _611_/B _612_/B _613_/B _614_/B _326_/A _615_/B _616_/B _617_/B
+ _618_/B _619_/B _620_/B _621_/B _622_/B _623_/B _624_/B _327_/A _625_/A _164_/A
+ _165_/A _166_/A _167_/A _168_/A _169_/A _170_/A _171_/A _172_/A _328_/A _173_/A
+ _174_/A _175_/A _176_/A _177_/A _178_/A _179_/A _180_/A _181_/A _182_/A _329_/A
+ _183_/A _184_/A _185_/A _186_/A _187_/A _188_/A _189_/A _190_/A _191_/A _192_/A
+ _330_/A _193_/A _194_/A _195_/A _196_/A _197_/A _198_/A _199_/A _200_/A _201_/A
+ _202_/A _331_/A _203_/A _204_/A _205_/A _206_/A _207_/A _208_/A _209_/A _210_/A
+ _211_/A _212_/A _332_/A _213_/A _214_/A _215_/A _216_/A _217_/A _218_/A _219_/A
+ _220_/A _221_/A _222_/A _333_/A _223_/A _224_/A _225_/A _226_/A _227_/A _228_/A
+ _229_/A _230_/A _231_/A _232_/A _334_/A _298_/A _233_/A _234_/A _235_/A _236_/A
+ _237_/A _238_/A _239_/A _240_/A _241_/A _242_/A _335_/A _243_/A _244_/A _245_/A
+ _246_/A _247_/A _248_/A _249_/A _250_/A _251_/A _252_/A _336_/A _253_/A _254_/A
+ _255_/A _256_/A _257_/A _258_/A _259_/A _260_/A _261_/A _262_/A _337_/A _263_/A
+ _264_/A _265_/A _266_/A _267_/A _268_/A _269_/A _270_/A _271_/A _272_/A _338_/A
+ _273_/A _274_/A _275_/A _276_/A _277_/A _278_/A _279_/A _280_/A _281_/A _282_/A
+ _339_/A _283_/A _284_/A _285_/A _286_/A _287_/A _288_/A _289_/A _290_/A _291_/A
+ _292_/A _340_/A _293_/A output951/A _294_/A _341_/A _342_/A _343_/A _344_/A _299_/A
+ _345_/A _346_/A _347_/A _348_/A _349_/A _350_/A _351_/A _352_/A _353_/A _354_/A
+ _300_/A _355_/A _356_/A _357_/A _358_/A _359_/A _360_/A _361_/A _362_/A _363_/A
+ _364_/A _301_/A _365_/A _366_/A _367_/A _368_/A _369_/B _370_/B _371_/B _372_/B
+ _373_/B _374_/B _302_/A _375_/B _376_/B _377_/B _378_/B _379_/B _380_/B _381_/B
+ _382_/B _383_/B _384_/B _303_/A _385_/B _386_/B _387_/B _388_/B _389_/B _390_/B
+ _391_/B _392_/B _393_/B _394_/B _304_/A vccd1_uq1 vssd1_uq1 mprj_logic_high
XTAP_3508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_508 _490_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_519 _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput200 la_iena_mprj[46] vssd vssd vccd vccd _209_/B sky130_fd_sc_hd__buf_4
XFILLER_20_3509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput211 la_iena_mprj[56] vssd vssd vccd vccd _219_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput222 la_iena_mprj[66] vssd vssd vccd vccd _229_/B sky130_fd_sc_hd__buf_4
XFILLER_0_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput233 la_iena_mprj[76] vssd vssd vccd vccd _239_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput244 la_iena_mprj[86] vssd vssd vccd vccd _249_/B sky130_fd_sc_hd__clkbuf_4
Xinput255 la_iena_mprj[96] vssd vssd vccd vccd _259_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput266 la_oenb_mprj[105] vssd vssd vccd vccd _602_/A sky130_fd_sc_hd__buf_6
XFILLER_40_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput277 la_oenb_mprj[115] vssd vssd vccd vccd _612_/A sky130_fd_sc_hd__buf_6
Xinput288 la_oenb_mprj[125] vssd vssd vccd vccd _622_/A sky130_fd_sc_hd__buf_6
XFILLER_40_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput299 la_oenb_mprj[1] vssd vssd vccd vccd _498_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_4019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_585_ _585_/A _585_/B vssd vssd vccd vccd _585_/X sky130_fd_sc_hd__and2_4
XFILLER_17_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput707 _155_/Y vssd vssd vccd vccd la_data_in_mprj[8] sky130_fd_sc_hd__buf_8
Xoutput718 _156_/Y vssd vssd vccd vccd la_data_in_mprj[9] sky130_fd_sc_hd__buf_8
XFILLER_10_2082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput729 _606_/X vssd vssd vccd vccd la_oenb_core[109] sky130_fd_sc_hd__buf_8
X_019_ _019_/A vssd vssd vccd vccd _019_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2120 _167_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2131 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2142 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2153 _278_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2164 _280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1430 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2175 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1441 _371_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2186 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2197 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1452 _373_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1463 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1474 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1485 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[61\] la_data_out_core[61] _224_/X vssd vssd vccd vccd _044_/A
+ sky130_fd_sc_hd__nand2_2
XANTENNA_1496 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3794 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_305 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_316 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_327 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_338 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_349 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_370_ _498_/A _370_/B _370_/C vssd vssd vccd vccd _370_/X sky130_fd_sc_hd__and3b_4
XTAP_1947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3460 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_850 _613_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_861 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_872 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_568_ _568_/A _568_/B vssd vssd vccd vccd _568_/X sky130_fd_sc_hd__and2_4
XANTENNA_883 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_894 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_499_ _499_/A _499_/B vssd vssd vccd vccd _499_/X sky130_fd_sc_hd__and2_4
XFILLER_31_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput504 _390_/X vssd vssd vccd vccd la_data_in_core[21] sky130_fd_sc_hd__buf_8
XFILLER_29_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput515 _400_/X vssd vssd vccd vccd la_data_in_core[31] sky130_fd_sc_hd__buf_8
XFILLER_44_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput526 _410_/X vssd vssd vccd vccd la_data_in_core[41] sky130_fd_sc_hd__buf_8
Xoutput537 _420_/X vssd vssd vccd vccd la_data_in_core[51] sky130_fd_sc_hd__buf_8
Xoutput548 _430_/X vssd vssd vccd vccd la_data_in_core[61] sky130_fd_sc_hd__buf_8
XFILLER_5_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput559 _440_/X vssd vssd vccd vccd la_data_in_core[71] sky130_fd_sc_hd__buf_8
XFILLER_5_991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1260 _273_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1271 _275_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1282 _276_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1293 _279_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_534 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_578 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3834 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_113 mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_146 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_422_ _550_/A _422_/B _422_/C vssd vssd vccd vccd _422_/X sky130_fd_sc_hd__and3b_4
XTAP_1722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3588 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_179 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3110 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_353_ _353_/A _353_/B vssd vssd vccd vccd _353_/X sky130_fd_sc_hd__and2_4
XTAP_1788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_284_ _284_/A _284_/B vssd vssd vccd vccd _284_/X sky130_fd_sc_hd__and2_4
XFILLER_52_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[7\] mprj_dat_i_user[7] _294_/X vssd vssd vccd vccd _121_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput8 la_data_out_mprj[103] vssd vssd vccd vccd _472_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_139 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_680 _576_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_691 _582_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[24\] la_data_out_core[24] _187_/X vssd vssd vccd vccd _007_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_36_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1886 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3731 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1090 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput890 _132_/Y vssd vssd vccd vccd mprj_dat_i_core[18] sky130_fd_sc_hd__buf_8
XFILLER_43_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2075 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4168 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_4518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3352 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_405_ _533_/A _405_/B _405_/C vssd vssd vccd vccd _405_/X sky130_fd_sc_hd__and3b_4
XTAP_1552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_336_ _336_/A _336_/B vssd vssd vccd vccd _336_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_267_ _267_/A _267_/B vssd vssd vccd vccd _267_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_198_ _198_/A _198_/B vssd vssd vccd vccd _198_/X sky130_fd_sc_hd__and2_2
XFILLER_45_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_13 la_data_out_core[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_24 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_35 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_46 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_57 mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_68 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_79 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_121_ _121_/A vssd vssd vccd vccd _121_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_4311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_052_ _052_/A vssd vssd vccd vccd _052_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1766 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2505 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2516 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2527 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_2538 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1804 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2549 _362_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1815 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1826 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1837 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1848 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1859 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xpowergood_check output954/A output952/A powergood_check/vccd powergood_check/vssd
+ powergood_check/vdda1 powergood_check/vssa1 powergood_check/vdda2 powergood_check/vssa2
+ mgmt_protect_hv
XFILLER_19_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_319_ _319_/A _319_/B vssd vssd vccd vccd _319_/X sky130_fd_sc_hd__and2_4
XFILLER_50_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput11 la_data_out_mprj[106] vssd vssd vccd vccd _475_/C sky130_fd_sc_hd__clkbuf_4
Xinput22 la_data_out_mprj[116] vssd vssd vccd vccd _485_/C sky130_fd_sc_hd__clkbuf_4
Xinput33 la_data_out_mprj[126] vssd vssd vccd vccd _495_/C sky130_fd_sc_hd__clkbuf_8
Xinput44 la_data_out_mprj[20] vssd vssd vccd vccd _389_/C sky130_fd_sc_hd__clkbuf_4
Xinput55 la_data_out_mprj[30] vssd vssd vccd vccd _399_/C sky130_fd_sc_hd__clkbuf_4
Xinput66 la_data_out_mprj[40] vssd vssd vccd vccd _409_/C sky130_fd_sc_hd__clkbuf_4
Xinput77 la_data_out_mprj[50] vssd vssd vccd vccd _419_/C sky130_fd_sc_hd__buf_4
XFILLER_45_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput88 la_data_out_mprj[60] vssd vssd vccd vccd _429_/C sky130_fd_sc_hd__clkbuf_4
Xinput99 la_data_out_mprj[70] vssd vssd vccd vccd _439_/C sky130_fd_sc_hd__buf_6
XFILLER_28_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[91\] la_data_out_core[91] _254_/X vssd vssd vccd vccd _074_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_48_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_426 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput404 mprj_adr_o_core[24] vssd vssd vccd vccd _329_/B sky130_fd_sc_hd__buf_8
XFILLER_40_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput415 mprj_adr_o_core[5] vssd vssd vccd vccd _310_/B sky130_fd_sc_hd__buf_8
XFILLER_44_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput426 mprj_dat_o_core[14] vssd vssd vccd vccd _351_/B sky130_fd_sc_hd__buf_8
XFILLER_22_4296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput437 mprj_dat_o_core[24] vssd vssd vccd vccd _361_/B sky130_fd_sc_hd__buf_8
XFILLER_40_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput448 mprj_dat_o_core[5] vssd vssd vccd vccd _342_/B sky130_fd_sc_hd__buf_8
Xinput459 mprj_we_o_core vssd vssd vccd vccd _300_/B sky130_fd_sc_hd__buf_8
XFILLER_2_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4034 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_104_ _104_/A vssd vssd vccd vccd _104_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_8_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_035_ _035_/A vssd vssd vccd vccd _035_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2302 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2313 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_2324 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2335 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2346 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1601 _603_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2357 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1612 _616_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1623 _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2368 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2379 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1634 _564_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1645 _576_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1656 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1667 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1678 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1689 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_509 _490_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3898 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput201 la_iena_mprj[47] vssd vssd vccd vccd _210_/B sky130_fd_sc_hd__buf_4
XFILLER_27_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput212 la_iena_mprj[57] vssd vssd vccd vccd _220_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput223 la_iena_mprj[67] vssd vssd vccd vccd _230_/B sky130_fd_sc_hd__buf_4
XTAP_4700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput234 la_iena_mprj[77] vssd vssd vccd vccd _240_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput245 la_iena_mprj[87] vssd vssd vccd vccd _250_/B sky130_fd_sc_hd__clkbuf_4
Xinput256 la_iena_mprj[97] vssd vssd vccd vccd _260_/B sky130_fd_sc_hd__clkbuf_4
Xinput267 la_oenb_mprj[106] vssd vssd vccd vccd _603_/A sky130_fd_sc_hd__buf_6
XFILLER_22_3392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput278 la_oenb_mprj[116] vssd vssd vccd vccd _613_/A sky130_fd_sc_hd__buf_6
Xinput289 la_oenb_mprj[126] vssd vssd vccd vccd _623_/A sky130_fd_sc_hd__buf_6
XFILLER_2_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_584_ _584_/A _584_/B vssd vssd vccd vccd _584_/X sky130_fd_sc_hd__and2_4
XFILLER_16_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput708 _073_/Y vssd vssd vccd vccd la_data_in_mprj[90] sky130_fd_sc_hd__buf_8
Xoutput719 _497_/X vssd vssd vccd vccd la_oenb_core[0] sky130_fd_sc_hd__buf_8
X_018_ _018_/A vssd vssd vccd vccd _018_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_2110 _165_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2121 _167_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2132 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2143 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2154 _278_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2165 _280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1420 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1431 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2176 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1442 _371_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2187 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2198 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1453 _373_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1464 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1475 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1486 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1497 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[54\] la_data_out_core[54] _217_/X vssd vssd vccd vccd _037_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_48_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_306 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_317 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_328 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_339 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_840 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_851 _614_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_567_ _567_/A _567_/B vssd vssd vccd vccd _567_/X sky130_fd_sc_hd__and2_4
XFILLER_32_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_862 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_873 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_884 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_895 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_498_ _498_/A _498_/B vssd vssd vccd vccd _498_/X sky130_fd_sc_hd__and2_4
XFILLER_18_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput505 _391_/X vssd vssd vccd vccd la_data_in_core[22] sky130_fd_sc_hd__buf_8
Xoutput516 _401_/X vssd vssd vccd vccd la_data_in_core[32] sky130_fd_sc_hd__buf_8
Xoutput527 _411_/X vssd vssd vccd vccd la_data_in_core[42] sky130_fd_sc_hd__buf_8
XFILLER_29_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput538 _421_/X vssd vssd vccd vccd la_data_in_core[52] sky130_fd_sc_hd__buf_8
Xoutput549 _431_/X vssd vssd vccd vccd la_data_in_core[62] sky130_fd_sc_hd__buf_8
XFILLER_42_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1250 _272_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1261 _273_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1272 _275_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1283 _276_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1294 _279_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3683 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3846 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_103 mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_125 mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_421_ _549_/A _421_/B _421_/C vssd vssd vccd vccd _421_/X sky130_fd_sc_hd__and3b_4
XTAP_1712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_136 mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_169 mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_352_ _352_/A _352_/B vssd vssd vccd vccd _352_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3122 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ _283_/A _283_/B vssd vssd vccd vccd _283_/X sky130_fd_sc_hd__and2_4
XFILLER_52_2470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput9 la_data_out_mprj[104] vssd vssd vccd vccd _473_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_619_ _619_/A _619_/B vssd vssd vccd vccd _619_/X sky130_fd_sc_hd__and2_4
XFILLER_35_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_670 _574_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_681 _576_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_692 _582_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[17\] la_data_out_core[17] _180_/X vssd vssd vccd vccd _000_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_31_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1832 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1080 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1091 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1054 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput880 _298_/X vssd vssd vccd vccd mprj_cyc_o_user sky130_fd_sc_hd__buf_8
XFILLER_21_4136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput891 _133_/Y vssd vssd vccd vccd mprj_dat_i_core[19] sky130_fd_sc_hd__buf_8
XFILLER_25_3571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_4032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_126 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_404_ _532_/A _404_/B _404_/C vssd vssd vccd vccd _404_/X sky130_fd_sc_hd__and3b_4
XPHY_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_335_ _335_/A _335_/B vssd vssd vccd vccd _335_/X sky130_fd_sc_hd__and2_2
XFILLER_30_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_266_ _266_/A _266_/B vssd vssd vccd vccd _266_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_197_ _197_/A _197_/B vssd vssd vccd vccd _197_/X sky130_fd_sc_hd__and2_1
XFILLER_10_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1139 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_14 la_data_out_core[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_25 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_36 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_47 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_58 mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_69 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_120_ _120_/A vssd vssd vccd vccd _120_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_051_ _051_/A vssd vssd vccd vccd _051_/Y sky130_fd_sc_hd__inv_4
XFILLER_49_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1723 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2506 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2517 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3666 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2528 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2539 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1805 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1816 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1827 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_1838 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1849 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_630 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_318_ _318_/A _318_/B vssd vssd vccd vccd _318_/X sky130_fd_sc_hd__and2_4
Xinput12 la_data_out_mprj[107] vssd vssd vccd vccd _476_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_30_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput23 la_data_out_mprj[117] vssd vssd vccd vccd _486_/C sky130_fd_sc_hd__clkbuf_4
Xinput34 la_data_out_mprj[127] vssd vssd vccd vccd _496_/C sky130_fd_sc_hd__clkbuf_8
Xinput45 la_data_out_mprj[21] vssd vssd vccd vccd _390_/C sky130_fd_sc_hd__clkbuf_4
X_249_ _249_/A _249_/B vssd vssd vccd vccd _249_/X sky130_fd_sc_hd__and2_4
XFILLER_45_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput56 la_data_out_mprj[31] vssd vssd vccd vccd _400_/C sky130_fd_sc_hd__clkbuf_4
Xinput67 la_data_out_mprj[41] vssd vssd vccd vccd _410_/C sky130_fd_sc_hd__clkbuf_4
Xinput78 la_data_out_mprj[51] vssd vssd vccd vccd _420_/C sky130_fd_sc_hd__buf_4
Xinput89 la_data_out_mprj[61] vssd vssd vccd vccd _430_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_45_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[84\] la_data_out_core[84] _247_/X vssd vssd vccd vccd _067_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_44_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3824 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput405 mprj_adr_o_core[25] vssd vssd vccd vccd _330_/B sky130_fd_sc_hd__buf_8
XFILLER_40_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput416 mprj_adr_o_core[6] vssd vssd vccd vccd _311_/B sky130_fd_sc_hd__buf_8
XFILLER_2_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput427 mprj_dat_o_core[15] vssd vssd vccd vccd _352_/B sky130_fd_sc_hd__buf_8
XFILLER_44_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput438 mprj_dat_o_core[25] vssd vssd vccd vccd _362_/B sky130_fd_sc_hd__buf_8
XFILLER_5_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput449 mprj_dat_o_core[6] vssd vssd vccd vccd _343_/B sky130_fd_sc_hd__buf_8
XFILLER_9_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4046 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_4418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_103_ _103_/A vssd vssd vccd vccd _103_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_034_ _034_/A vssd vssd vccd vccd _034_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_4225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2303 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2314 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2325 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2336 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2347 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1602 _604_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2751 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2358 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1613 _617_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1624 _532_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2369 _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1635 _564_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1646 _577_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1657 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1668 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1679 _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[12\] mprj_dat_i_user[12] _294_/X vssd vssd vccd vccd _126_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[110\] la_data_out_core[110] _273_/X vssd vssd vccd vccd _093_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_27_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4462 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput202 la_iena_mprj[48] vssd vssd vccd vccd _211_/B sky130_fd_sc_hd__buf_4
Xinput213 la_iena_mprj[58] vssd vssd vccd vccd _221_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4083 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput224 la_iena_mprj[68] vssd vssd vccd vccd _231_/B sky130_fd_sc_hd__buf_4
XTAP_4701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput235 la_iena_mprj[78] vssd vssd vccd vccd _241_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_4188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput246 la_iena_mprj[88] vssd vssd vccd vccd _251_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput257 la_iena_mprj[98] vssd vssd vccd vccd _261_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput268 la_oenb_mprj[107] vssd vssd vccd vccd _604_/A sky130_fd_sc_hd__buf_6
XFILLER_40_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput279 la_oenb_mprj[117] vssd vssd vccd vccd _614_/A sky130_fd_sc_hd__buf_6
XFILLER_2_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_583_ _583_/A _583_/B vssd vssd vccd vccd _583_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_3608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput709 _074_/Y vssd vssd vccd vccd la_data_in_mprj[91] sky130_fd_sc_hd__buf_8
XFILLER_29_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_017_ _017_/A vssd vssd vccd vccd _017_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_46_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2100 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_2111 _165_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2122 _167_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2133 _204_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2144 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1410 _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2155 _278_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2166 _280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1421 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1432 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2177 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1443 _371_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2188 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2199 _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1454 _373_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1465 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1476 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1487 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1498 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[47\] la_data_out_core[47] _210_/X vssd vssd vccd vccd _030_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_14_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[9\] la_data_out_core[9] _172_/X vssd vssd vccd vccd _156_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_41_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1727 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_307 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4130 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_318 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_329 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_830 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_841 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_852 _614_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_566_ _566_/A _566_/B vssd vssd vccd vccd _566_/X sky130_fd_sc_hd__and2_4
XANTENNA_863 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_874 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_885 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_896 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_497_ _497_/A _497_/B vssd vssd vccd vccd _497_/X sky130_fd_sc_hd__and2_4
XFILLER_38_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput506 _392_/X vssd vssd vccd vccd la_data_in_core[23] sky130_fd_sc_hd__buf_8
Xoutput517 _402_/X vssd vssd vccd vccd la_data_in_core[33] sky130_fd_sc_hd__buf_8
Xoutput528 _412_/X vssd vssd vccd vccd la_data_in_core[43] sky130_fd_sc_hd__buf_8
XFILLER_9_2704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput539 _422_/X vssd vssd vccd vccd la_data_in_core[53] sky130_fd_sc_hd__buf_8
XFILLER_29_1920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1240 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1251 _272_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1262 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1273 _275_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1284 _276_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1295 _279_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_104 mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_420_ _548_/A _420_/B _420_/C vssd vssd vccd vccd _420_/X sky130_fd_sc_hd__and3b_4
XANTENNA_137 mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_351_ _351_/A _351_/B vssd vssd vccd vccd _351_/X sky130_fd_sc_hd__and2_4
XFILLER_42_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_282_ _282_/A _282_/B vssd vssd vccd vccd _282_/X sky130_fd_sc_hd__and2_2
XFILLER_30_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3296 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_618_ _618_/A _618_/B vssd vssd vccd vccd _618_/X sky130_fd_sc_hd__and2_4
XTAP_3693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_660 _569_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_671 _574_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_549_ _549_/A _549_/B vssd vssd vccd vccd _549_/X sky130_fd_sc_hd__and2_4
XFILLER_18_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_682 _576_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_693 _582_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1070 _182_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1081 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_606 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1092 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput870 _307_/X vssd vssd vccd vccd mprj_adr_o_user[2] sky130_fd_sc_hd__buf_8
XFILLER_5_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput881 _114_/Y vssd vssd vccd vccd mprj_dat_i_core[0] sky130_fd_sc_hd__buf_8
XFILLER_5_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput892 _115_/Y vssd vssd vccd vccd mprj_dat_i_core[1] sky130_fd_sc_hd__buf_8
XFILLER_21_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_4066 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_403_ _531_/A _403_/B _403_/C vssd vssd vccd vccd _403_/X sky130_fd_sc_hd__and3b_4
XTAP_2277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_50 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_334_ _334_/A _334_/B vssd vssd vccd vccd _334_/X sky130_fd_sc_hd__and2_4
XTAP_1598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_265_ _265_/A _265_/B vssd vssd vccd vccd _265_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_196_ _196_/A _196_/B vssd vssd vccd vccd _196_/X sky130_fd_sc_hd__and2_2
XFILLER_41_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_406 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_490 _488_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_15 la_data_out_core[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_26 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_37 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_48 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_59 mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_318 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_050_ _050_/A vssd vssd vccd vccd _050_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_20_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2507 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2518 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2529 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3678 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1806 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1817 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1828 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1839 _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_642 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_317_ _317_/A _317_/B vssd vssd vccd vccd _317_/X sky130_fd_sc_hd__and2_4
XFILLER_50_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput13 la_data_out_mprj[108] vssd vssd vccd vccd _477_/C sky130_fd_sc_hd__clkbuf_4
Xinput24 la_data_out_mprj[118] vssd vssd vccd vccd _487_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_248_ _248_/A _248_/B vssd vssd vccd vccd _248_/X sky130_fd_sc_hd__and2_4
XFILLER_7_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput35 la_data_out_mprj[12] vssd vssd vccd vccd _381_/C sky130_fd_sc_hd__clkbuf_4
Xinput46 la_data_out_mprj[22] vssd vssd vccd vccd _391_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput57 la_data_out_mprj[32] vssd vssd vccd vccd _401_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_32_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput68 la_data_out_mprj[42] vssd vssd vccd vccd _411_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_32_1993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput79 la_data_out_mprj[52] vssd vssd vccd vccd _421_/C sky130_fd_sc_hd__buf_4
X_179_ _179_/A _179_/B vssd vssd vccd vccd _179_/X sky130_fd_sc_hd__and2_2
XFILLER_13_1392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[77\] la_data_out_core[77] _240_/X vssd vssd vccd vccd _060_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_22_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput406 mprj_adr_o_core[26] vssd vssd vccd vccd _331_/B sky130_fd_sc_hd__buf_8
XFILLER_22_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput417 mprj_adr_o_core[7] vssd vssd vccd vccd _312_/B sky130_fd_sc_hd__buf_8
Xinput428 mprj_dat_o_core[16] vssd vssd vccd vccd _353_/B sky130_fd_sc_hd__buf_8
XFILLER_22_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput439 mprj_dat_o_core[26] vssd vssd vccd vccd _363_/B sky130_fd_sc_hd__buf_8
XFILLER_29_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_102_ _102_/A vssd vssd vccd vccd _102_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_33_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_033_ _033_/A vssd vssd vccd vccd _033_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_4_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2304 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2315 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2326 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2337 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2348 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1603 _605_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1614 _617_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2763 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2359 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1625 _533_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1636 _568_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1647 _585_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1658 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_1669 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[103\] la_data_out_core[103] _266_/X vssd vssd vccd vccd _086_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_26_715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput203 la_iena_mprj[49] vssd vssd vccd vccd _212_/B sky130_fd_sc_hd__buf_4
XFILLER_44_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput214 la_iena_mprj[59] vssd vssd vccd vccd _222_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2947 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput225 la_iena_mprj[69] vssd vssd vccd vccd _232_/B sky130_fd_sc_hd__buf_4
XFILLER_22_4095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput236 la_iena_mprj[79] vssd vssd vccd vccd _242_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput247 la_iena_mprj[89] vssd vssd vccd vccd _252_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput258 la_iena_mprj[99] vssd vssd vccd vccd _262_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput269 la_oenb_mprj[108] vssd vssd vccd vccd _605_/A sky130_fd_sc_hd__buf_6
XFILLER_18_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_542 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_582_ _582_/A _582_/B vssd vssd vccd vccd _582_/X sky130_fd_sc_hd__and2_4
XFILLER_17_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_016_ _016_/A vssd vssd vccd vccd _016_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2074 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2101 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2112 _165_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2123 _167_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2134 _218_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2145 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1400 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2156 _278_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1411 _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2167 _280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1422 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1433 _369_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2178 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1444 _371_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2189 _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1455 _374_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1466 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1477 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1488 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1499 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_980 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1739 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_308 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_319 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1850 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_820 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_831 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_842 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_565_ _565_/A _565_/B vssd vssd vccd vccd _565_/X sky130_fd_sc_hd__and2_4
XFILLER_18_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_853 _614_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_864 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_875 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_886 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_496_ _624_/A _496_/B _496_/C vssd vssd vccd vccd _496_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_897 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput507 _393_/X vssd vssd vccd vccd la_data_in_core[24] sky130_fd_sc_hd__buf_8
XFILLER_9_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput518 _403_/X vssd vssd vccd vccd la_data_in_core[34] sky130_fd_sc_hd__buf_8
XFILLER_29_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput529 _413_/X vssd vssd vccd vccd la_data_in_core[44] sky130_fd_sc_hd__buf_8
XFILLER_42_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1932 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1230 _262_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1241 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1252 _272_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1263 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1274 _275_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1285 _276_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1296 _279_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1102 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_105 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_116 mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_149 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ _350_/A _350_/B vssd vssd vccd vccd _350_/X sky130_fd_sc_hd__and2_4
XTAP_1758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_281_ _281_/A _281_/B vssd vssd vccd vccd _281_/X sky130_fd_sc_hd__and2_4
XFILLER_39_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_617_ _617_/A _617_/B vssd vssd vccd vccd _617_/X sky130_fd_sc_hd__and2_4
XFILLER_45_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_650 _568_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_661 _569_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_548_ _548_/A _548_/B vssd vssd vccd vccd _548_/X sky130_fd_sc_hd__and2_4
XFILLER_53_2225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_672 _574_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_683 _576_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_694 _582_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_479_ _607_/A _479_/B _479_/C vssd vssd vccd vccd _479_/X sky130_fd_sc_hd__and3b_4
XFILLER_20_518 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2502 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4352 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1060 _176_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1071 _182_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1082 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1093 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1906 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput860 _325_/X vssd vssd vccd vccd mprj_adr_o_user[20] sky130_fd_sc_hd__buf_8
Xoutput871 _335_/X vssd vssd vccd vccd mprj_adr_o_user[30] sky130_fd_sc_hd__buf_8
Xoutput882 _124_/Y vssd vssd vccd vccd mprj_dat_i_core[10] sky130_fd_sc_hd__buf_8
XFILLER_8_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput893 _134_/Y vssd vssd vccd vccd mprj_dat_i_core[20] sky130_fd_sc_hd__buf_8
XFILLER_5_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4070 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3344 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_402_ _530_/A _402_/B _402_/C vssd vssd vccd vccd _402_/X sky130_fd_sc_hd__and3b_4
XTAP_1522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_333_ _333_/A _333_/B vssd vssd vccd vccd _333_/X sky130_fd_sc_hd__and2_4
XTAP_1588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_264_ _264_/A _264_/B vssd vssd vccd vccd _264_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_195_ _195_/A _195_/B vssd vssd vccd vccd _195_/X sky130_fd_sc_hd__and2_2
XFILLER_6_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[5\] mprj_dat_i_user[5] _294_/X vssd vssd vccd vccd _119_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_794 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_480 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[22\] la_data_out_core[22] _185_/X vssd vssd vccd vccd _005_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_36_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_491 _488_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3764 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_16 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_27 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_38 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_49 mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3954 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2508 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4514 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2519 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1807 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1818 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1829 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput690 _057_/Y vssd vssd vccd vccd la_data_in_mprj[74] sky130_fd_sc_hd__buf_8
XFILLER_40_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_654 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_316_ _316_/A _316_/B vssd vssd vccd vccd _316_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput14 la_data_out_mprj[109] vssd vssd vccd vccd _478_/C sky130_fd_sc_hd__clkbuf_4
X_247_ _247_/A _247_/B vssd vssd vccd vccd _247_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput25 la_data_out_mprj[119] vssd vssd vccd vccd _488_/C sky130_fd_sc_hd__clkbuf_4
Xinput36 la_data_out_mprj[13] vssd vssd vccd vccd _382_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_45_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput47 la_data_out_mprj[23] vssd vssd vccd vccd _392_/C sky130_fd_sc_hd__clkbuf_4
Xinput58 la_data_out_mprj[33] vssd vssd vccd vccd _402_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_48_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput69 la_data_out_mprj[43] vssd vssd vccd vccd _412_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3694 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_178_ _178_/A _178_/B vssd vssd vccd vccd _178_/X sky130_fd_sc_hd__and2_2
XFILLER_7_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput407 mprj_adr_o_core[27] vssd vssd vccd vccd _332_/B sky130_fd_sc_hd__buf_8
XFILLER_5_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput418 mprj_adr_o_core[8] vssd vssd vccd vccd _313_/B sky130_fd_sc_hd__buf_8
Xinput429 mprj_dat_o_core[17] vssd vssd vccd vccd _354_/B sky130_fd_sc_hd__buf_8
XFILLER_2_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_101_ _101_/A vssd vssd vccd vccd _101_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_032_ _032_/A vssd vssd vccd vccd _032_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_3719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2305 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2316 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2327 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2338 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1604 _607_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2349 mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1615 _619_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1626 _534_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2775 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1637 _568_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1648 _586_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1659 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_727 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_988 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput204 la_iena_mprj[4] vssd vssd vccd vccd _167_/B sky130_fd_sc_hd__clkbuf_4
Xinput215 la_iena_mprj[5] vssd vssd vccd vccd _168_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput226 la_iena_mprj[6] vssd vssd vccd vccd _169_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2959 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput237 la_iena_mprj[7] vssd vssd vccd vccd _170_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput248 la_iena_mprj[8] vssd vssd vccd vccd _171_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput259 la_iena_mprj[9] vssd vssd vccd vccd _172_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1072 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_581_ _581_/A _581_/B vssd vssd vccd vccd _581_/X sky130_fd_sc_hd__and2_4
XFILLER_38_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_015_ _015_/A vssd vssd vccd vccd _015_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2102 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2113 _165_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2124 _167_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2135 _218_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1401 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2146 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2157 _278_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1412 _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2168 _280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1423 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1434 _369_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2179 _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1445 _371_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1456 _374_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1467 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1478 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1489 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_992 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3903 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3682 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1990 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_309 _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4078 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_810 _608_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_821 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_832 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_564_ _564_/A _564_/B vssd vssd vccd vccd _564_/X sky130_fd_sc_hd__and2_2
XTAP_3898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_843 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_854 _614_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_865 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_876 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_495_ _623_/A _495_/B _495_/C vssd vssd vccd vccd _495_/X sky130_fd_sc_hd__and3b_4
XANTENNA_887 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_898 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput508 _394_/X vssd vssd vccd vccd la_data_in_core[25] sky130_fd_sc_hd__buf_8
XFILLER_5_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput519 _404_/X vssd vssd vccd vccd la_data_in_core[35] sky130_fd_sc_hd__buf_8
XFILLER_49_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1220 _256_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_ack_gate mprj_ack_i_user _294_/X vssd vssd vccd vccd _146_/A sky130_fd_sc_hd__nand2_1
XANTENNA_1231 _262_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1242 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1253 _272_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1264 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1275 _275_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1286 _276_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1297 _279_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[52\] la_data_out_core[52] _215_/X vssd vssd vccd vccd _035_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_48_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_106 mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_128 mprj_dat_i_user[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_280_ _280_/A _280_/B vssd vssd vccd vccd _280_/X sky130_fd_sc_hd__and2_4
XFILLER_13_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1783 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2807 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_616_ _616_/A _616_/B vssd vssd vccd vccd _616_/X sky130_fd_sc_hd__and2_4
XTAP_3673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_640 _566_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_651 _568_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_547_ _547_/A _547_/B vssd vssd vccd vccd _547_/X sky130_fd_sc_hd__and2_4
XANTENNA_662 _569_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_673 _574_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_684 _577_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_695 _582_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_478_ _606_/A _478_/B _478_/C vssd vssd vccd vccd _478_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1050 _167_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1061 _176_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1072 _182_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1083 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1094 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3746 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_4231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3839 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput850 _316_/X vssd vssd vccd vccd mprj_adr_o_user[11] sky130_fd_sc_hd__buf_8
XFILLER_25_4275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput861 _326_/X vssd vssd vccd vccd mprj_adr_o_user[21] sky130_fd_sc_hd__buf_8
XFILLER_47_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput872 _336_/X vssd vssd vccd vccd mprj_adr_o_user[31] sky130_fd_sc_hd__buf_8
XFILLER_5_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput883 _125_/Y vssd vssd vccd vccd mprj_dat_i_core[11] sky130_fd_sc_hd__buf_8
Xoutput894 _135_/Y vssd vssd vccd vccd mprj_dat_i_core[21] sky130_fd_sc_hd__buf_8
XFILLER_43_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_401_ _529_/A _401_/B _401_/C vssd vssd vccd vccd _401_/X sky130_fd_sc_hd__and3b_4
XTAP_2257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_332_ _332_/A _332_/B vssd vssd vccd vccd _332_/X sky130_fd_sc_hd__and2_4
XTAP_1578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_263_ _263_/A _263_/B vssd vssd vccd vccd _263_/X sky130_fd_sc_hd__and2_4
XFILLER_6_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_194_ _194_/A _194_/B vssd vssd vccd vccd _194_/X sky130_fd_sc_hd__and2_1
XFILLER_6_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3994 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_470 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_481 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_492 _488_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_17 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_28 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_338 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[28\] mprj_dat_i_user[28] _294_/X vssd vssd vccd vccd _142_/A sky130_fd_sc_hd__nand2_2
Xuser_to_mprj_in_gates\[15\] la_data_out_core[15] _178_/X vssd vssd vccd vccd _162_/A
+ sky130_fd_sc_hd__nand2_2
XANTENNA_39 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[126\] la_data_out_core[126] _289_/X vssd vssd vccd vccd _109_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_20_4172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_964 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_2509 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_4526 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1808 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1819 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput680 _048_/Y vssd vssd vccd vccd la_data_in_mprj[65] sky130_fd_sc_hd__buf_8
XFILLER_27_2979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput691 _058_/Y vssd vssd vccd vccd la_data_in_mprj[75] sky130_fd_sc_hd__buf_8
XFILLER_43_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_315_ _315_/A _315_/B vssd vssd vccd vccd _315_/X sky130_fd_sc_hd__and2_4
XTAP_1397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_246_ _246_/A _246_/B vssd vssd vccd vccd _246_/X sky130_fd_sc_hd__and2_4
Xinput15 la_data_out_mprj[10] vssd vssd vccd vccd _379_/C sky130_fd_sc_hd__clkbuf_4
Xinput26 la_data_out_mprj[11] vssd vssd vccd vccd _380_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput37 la_data_out_mprj[14] vssd vssd vccd vccd _383_/C sky130_fd_sc_hd__clkbuf_4
Xinput48 la_data_out_mprj[24] vssd vssd vccd vccd _393_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_7_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput59 la_data_out_mprj[34] vssd vssd vccd vccd _403_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_45_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_177_ _177_/A _177_/B vssd vssd vccd vccd _177_/X sky130_fd_sc_hd__and2_4
XFILLER_32_1984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput408 mprj_adr_o_core[28] vssd vssd vccd vccd _333_/B sky130_fd_sc_hd__buf_8
XFILLER_44_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput419 mprj_adr_o_core[9] vssd vssd vccd vccd _314_/B sky130_fd_sc_hd__buf_8
XFILLER_2_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_100_ _100_/A vssd vssd vccd vccd _100_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_031_ _031_/A vssd vssd vccd vccd _031_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2306 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2317 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2328 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2339 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1605 _608_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1616 _620_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1627 _543_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1638 _570_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1649 _587_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_430 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_229_ _229_/A _229_/B vssd vssd vccd vccd _229_/X sky130_fd_sc_hd__and2_2
XFILLER_7_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[82\] la_data_out_core[82] _245_/X vssd vssd vccd vccd _065_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_44_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_739 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2803 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1832 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput205 la_iena_mprj[50] vssd vssd vccd vccd _213_/B sky130_fd_sc_hd__buf_4
XFILLER_22_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput216 la_iena_mprj[60] vssd vssd vccd vccd _223_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_41_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput227 la_iena_mprj[70] vssd vssd vccd vccd _233_/B sky130_fd_sc_hd__buf_4
XTAP_4704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput238 la_iena_mprj[80] vssd vssd vccd vccd _243_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput249 la_iena_mprj[90] vssd vssd vccd vccd _253_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_580_ _580_/A _580_/B vssd vssd vccd vccd _580_/X sky130_fd_sc_hd__and2_4
XFILLER_44_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_97 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_014_ _014_/A vssd vssd vccd vccd _014_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_46_4565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2103 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2114 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2125 _171_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2136 _260_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2147 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1402 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2158 _278_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1413 _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1424 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2169 _280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1435 _369_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1446 _372_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1457 _374_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1468 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1479 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1242 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_gates\[10\] mprj_dat_i_user[10] _294_/X vssd vssd vccd vccd _124_/A sky130_fd_sc_hd__nand2_1
XFILLER_45_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_4351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_1980 _362_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1991 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4024 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2779 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1830 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_800 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_811 _609_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_822 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_563_ _563_/A _563_/B vssd vssd vccd vccd _563_/X sky130_fd_sc_hd__and2_4
XTAP_3888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_833 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_844 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_855 _614_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_866 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_877 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_494_ _622_/A _494_/B _494_/C vssd vssd vccd vccd _494_/X sky130_fd_sc_hd__and3b_4
XANTENNA_888 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_899 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput509 _395_/X vssd vssd vccd vccd la_data_in_core[26] sky130_fd_sc_hd__buf_8
XFILLER_46_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1210 _246_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1221 _259_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1232 _262_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1243 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1254 _272_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1265 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1276 _275_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1287 _276_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1298 _279_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[45\] la_data_out_core[45] _208_/X vssd vssd vccd vccd _028_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_4355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[7\] la_data_out_core[7] _170_/X vssd vssd vccd vccd _154_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_5_3817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_118 mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 mprj_dat_i_user[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2819 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_615_ _615_/A _615_/B vssd vssd vccd vccd _615_/X sky130_fd_sc_hd__and2_4
XTAP_3663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_630 _549_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_641 _566_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_546_ _546_/A _546_/B vssd vssd vccd vccd _546_/X sky130_fd_sc_hd__and2_4
XANTENNA_652 _568_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_663 _570_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_674 _574_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_685 _578_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_696 _582_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_477_ _605_/A _477_/B _477_/C vssd vssd vccd vccd _477_/X sky130_fd_sc_hd__and3b_4
XFILLER_38_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1040 _165_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1051 _168_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1062 _176_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1073 _182_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1084 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1095 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3468 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput840 _591_/X vssd vssd vccd vccd la_oenb_core[94] sky130_fd_sc_hd__buf_8
XFILLER_5_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput851 _317_/X vssd vssd vccd vccd mprj_adr_o_user[12] sky130_fd_sc_hd__buf_8
XFILLER_43_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput862 _327_/X vssd vssd vccd vccd mprj_adr_o_user[22] sky130_fd_sc_hd__buf_8
XFILLER_25_4287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput873 _308_/X vssd vssd vccd vccd mprj_adr_o_user[3] sky130_fd_sc_hd__buf_8
Xoutput884 _126_/Y vssd vssd vccd vccd mprj_dat_i_core[12] sky130_fd_sc_hd__buf_8
Xoutput895 _136_/Y vssd vssd vccd vccd mprj_dat_i_core[22] sky130_fd_sc_hd__buf_8
XFILLER_43_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2863 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_400_ _528_/A _400_/B _400_/C vssd vssd vccd vccd _400_/X sky130_fd_sc_hd__and3b_4
XTAP_2247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_331_ _331_/A _331_/B vssd vssd vccd vccd _331_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_262_ _262_/A _262_/B vssd vssd vccd vccd _262_/X sky130_fd_sc_hd__and2_4
XFILLER_52_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_4545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_193_ _193_/A _193_/B vssd vssd vccd vccd _193_/X sky130_fd_sc_hd__and2_2
XFILLER_52_1570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_460 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_471 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_529_ _529_/A _529_/B vssd vssd vccd vccd _529_/X sky130_fd_sc_hd__and2_4
XFILLER_15_3733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_482 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_493 _488_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3788 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_18 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_29 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_4162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1699 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[119\] la_data_out_core[119] _282_/X vssd vssd vccd vccd _102_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_20_3494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_910 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4270 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4538 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1809 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput670 _039_/Y vssd vssd vccd vccd la_data_in_mprj[56] sky130_fd_sc_hd__buf_8
XFILLER_25_4095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput681 _049_/Y vssd vssd vccd vccd la_data_in_mprj[66] sky130_fd_sc_hd__buf_8
XFILLER_47_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput692 _059_/Y vssd vssd vccd vccd la_data_in_mprj[76] sky130_fd_sc_hd__buf_8
XFILLER_40_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_314_ _314_/A _314_/B vssd vssd vccd vccd _314_/X sky130_fd_sc_hd__and2_4
XTAP_1387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_245_ _245_/A _245_/B vssd vssd vccd vccd _245_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput16 la_data_out_mprj[110] vssd vssd vccd vccd _479_/C sky130_fd_sc_hd__clkbuf_4
Xinput27 la_data_out_mprj[120] vssd vssd vccd vccd _489_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_45_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput38 la_data_out_mprj[15] vssd vssd vccd vccd _384_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_6_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput49 la_data_out_mprj[25] vssd vssd vccd vccd _394_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3674 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_176_ _176_/A _176_/B vssd vssd vccd vccd _176_/X sky130_fd_sc_hd__and2_4
XFILLER_13_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_290 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput409 mprj_adr_o_core[29] vssd vssd vccd vccd _334_/B sky130_fd_sc_hd__buf_8
XFILLER_5_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4075 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_910 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_030_ _030_/A vssd vssd vccd vccd _030_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_3972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2307 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2318 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2329 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1606 _612_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1617 _621_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1628 _543_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1639 _570_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_228_ _228_/A _228_/B vssd vssd vccd vccd _228_/X sky130_fd_sc_hd__and2_2
XFILLER_7_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3482 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_159_ _159_/A vssd vssd vccd vccd _159_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[75\] la_data_out_core[75] _238_/X vssd vssd vccd vccd _058_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3683 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3382 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput206 la_iena_mprj[51] vssd vssd vccd vccd _214_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput217 la_iena_mprj[61] vssd vssd vccd vccd _224_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_48_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput228 la_iena_mprj[71] vssd vssd vccd vccd _234_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput239 la_iena_mprj[81] vssd vssd vccd vccd _244_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_013_ _013_/A vssd vssd vccd vccd _013_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2104 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2115 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2126 _187_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2137 _260_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2148 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1403 _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2159 _278_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1414 _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1425 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1436 _369_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1447 _372_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1458 _375_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1469 _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1254 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1970 _350_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1981 _363_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1992 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[101\] la_data_out_core[101] _264_/X vssd vssd vccd vccd _084_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_52_4036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_801 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_562_ _562_/A _562_/B vssd vssd vccd vccd _562_/X sky130_fd_sc_hd__and2_2
XTAP_3878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_812 _609_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_823 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_834 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_845 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_856 _326_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_493_ _621_/A _493_/B _493_/C vssd vssd vccd vccd _493_/X sky130_fd_sc_hd__and3b_4
XFILLER_44_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_867 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_878 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_889 _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1200 _233_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1211 _247_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1222 _260_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1233 _337_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1244 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1255 _272_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1266 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1277 _275_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1288 _278_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1299 _279_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[38\] la_data_out_core[38] _201_/X vssd vssd vccd vccd _021_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_18_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1516 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2490 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_846 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_108 mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_119 mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_614_ _614_/A _614_/B vssd vssd vccd vccd _614_/X sky130_fd_sc_hd__and2_4
XTAP_4398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_620 _517_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_631 _552_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_545_ _545_/A _545_/B vssd vssd vccd vccd _545_/X sky130_fd_sc_hd__and2_4
XANTENNA_642 _566_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_653 _568_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_664 _571_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_675 _576_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_686 _579_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_476_ _604_/A _476_/B _476_/C vssd vssd vccd vccd _476_/X sky130_fd_sc_hd__and3b_4
XANTENNA_697 _582_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1030 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1041 _165_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1052 _169_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1063 _177_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1074 _182_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1085 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1096 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput830 _582_/X vssd vssd vccd vccd la_oenb_core[85] sky130_fd_sc_hd__buf_8
XFILLER_25_4255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput841 _592_/X vssd vssd vccd vccd la_oenb_core[95] sky130_fd_sc_hd__buf_8
Xoutput852 _318_/X vssd vssd vccd vccd mprj_adr_o_user[13] sky130_fd_sc_hd__buf_8
XFILLER_47_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput863 _328_/X vssd vssd vccd vccd mprj_adr_o_user[23] sky130_fd_sc_hd__buf_8
Xoutput874 _309_/X vssd vssd vccd vccd mprj_adr_o_user[4] sky130_fd_sc_hd__buf_8
XFILLER_8_2037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput885 _127_/Y vssd vssd vccd vccd mprj_dat_i_core[13] sky130_fd_sc_hd__buf_8
XFILLER_8_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput896 _137_/Y vssd vssd vccd vccd mprj_dat_i_core[23] sky130_fd_sc_hd__buf_8
XFILLER_25_2831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2875 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_698 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_43 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_330_ _330_/A _330_/B vssd vssd vccd vccd _330_/X sky130_fd_sc_hd__and2_4
XFILLER_42_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_261_ _261_/A _261_/B vssd vssd vccd vccd _261_/X sky130_fd_sc_hd__and2_4
XFILLER_39_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_192_ _192_/A _192_/B vssd vssd vccd vccd _192_/X sky130_fd_sc_hd__and2_2
XFILLER_48_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_731 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_450 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_461 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_472 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_528_ _528_/A _528_/B vssd vssd vccd vccd _528_/X sky130_fd_sc_hd__and2_4
XFILLER_50_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_483 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_494 _488_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_459_ _587_/A _459_/B _459_/C vssd vssd vccd vccd _459_/X sky130_fd_sc_hd__and3b_4
XANTENNA_19 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_3200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2576 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4282 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4063 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput660 _030_/Y vssd vssd vccd vccd la_data_in_mprj[47] sky130_fd_sc_hd__buf_8
XFILLER_25_3340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput671 _040_/Y vssd vssd vccd vccd la_data_in_mprj[57] sky130_fd_sc_hd__buf_8
Xoutput682 _050_/Y vssd vssd vccd vccd la_data_in_mprj[67] sky130_fd_sc_hd__buf_8
XFILLER_21_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput693 _060_/Y vssd vssd vccd vccd la_data_in_mprj[77] sky130_fd_sc_hd__buf_8
XFILLER_8_1111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_313_ _313_/A _313_/B vssd vssd vccd vccd _313_/X sky130_fd_sc_hd__and2_4
XFILLER_30_616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2080 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_244_ _244_/A _244_/B vssd vssd vccd vccd _244_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput17 la_data_out_mprj[111] vssd vssd vccd vccd _480_/C sky130_fd_sc_hd__buf_4
XFILLER_32_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput28 la_data_out_mprj[121] vssd vssd vccd vccd _490_/C sky130_fd_sc_hd__clkbuf_4
Xinput39 la_data_out_mprj[16] vssd vssd vccd vccd _385_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_45_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_175_ _175_/A _175_/B vssd vssd vccd vccd _175_/X sky130_fd_sc_hd__and2_4
XFILLER_6_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[3\] mprj_dat_i_user[3] _294_/X vssd vssd vccd vccd _117_/A sky130_fd_sc_hd__nand2_1
XFILLER_10_3686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_280 _449_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_291 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[20\] la_data_out_core[20] _183_/X vssd vssd vccd vccd _003_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_15_3564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4018 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_410 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2308 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2319 mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1607 _612_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1618 _623_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1629 _551_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput490 _493_/X vssd vssd vccd vccd la_data_in_core[124] sky130_fd_sc_hd__buf_8
XFILLER_43_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_227_ _227_/A _227_/B vssd vssd vccd vccd _227_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_158_ _158_/A vssd vssd vccd vccd _158_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_089_ _089_/A vssd vssd vccd vccd _089_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4280 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[68\] la_data_out_core[68] _231_/X vssd vssd vccd vccd _051_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_22_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_516 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3394 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_4191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4066 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput207 la_iena_mprj[52] vssd vssd vccd vccd _215_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput218 la_iena_mprj[62] vssd vssd vccd vccd _225_/B sky130_fd_sc_hd__buf_4
XFILLER_41_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput229 la_iena_mprj[72] vssd vssd vccd vccd _235_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2012 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_012_ _012_/A vssd vssd vccd vccd _012_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2105 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2116 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2127 _193_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2138 _260_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2149 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1404 _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1415 _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1426 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1437 _369_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1448 _372_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1459 _375_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1266 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_490 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1960 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1971 _351_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1982 _366_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1993 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_4168 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_802 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_561_ _561_/A _561_/B vssd vssd vccd vccd _561_/X sky130_fd_sc_hd__and2_4
XTAP_3868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_813 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_824 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_835 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_846 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_492_ _620_/A _492_/B _492_/C vssd vssd vccd vccd _492_/X sky130_fd_sc_hd__and3b_4
XANTENNA_857 _615_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_868 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_879 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3040 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1936 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1201 _233_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1212 _248_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1223 _261_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1234 _266_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1245 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1256 _272_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1267 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1278 _275_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1289 _278_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_4466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1052 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2480 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2491 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1790 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_858 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_613_ _613_/A _613_/B vssd vssd vccd vccd _613_/X sky130_fd_sc_hd__and2_4
XTAP_4388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_610 _511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_621 _518_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_632 _552_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_544_ _544_/A _544_/B vssd vssd vccd vccd _544_/X sky130_fd_sc_hd__and2_4
XTAP_2942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_643 _567_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_654 _568_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_665 _574_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_676 _576_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_687 _579_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_475_ _603_/A _475_/B _475_/C vssd vssd vccd vccd _475_/X sky130_fd_sc_hd__and3b_4
XFILLER_15_3949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_698 _583_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3830 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1020 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1031 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1042 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1053 _170_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1064 _178_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1075 _182_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1086 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1097 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3738 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput390 mprj_adr_o_core[11] vssd vssd vccd vccd _316_/B sky130_fd_sc_hd__buf_8
XFILLER_3_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[50\] la_data_out_core[50] _213_/X vssd vssd vccd vccd _033_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_18_4252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2026 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput820 _573_/X vssd vssd vccd vccd la_oenb_core[76] sky130_fd_sc_hd__buf_8
XFILLER_47_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput831 _583_/X vssd vssd vccd vccd la_oenb_core[86] sky130_fd_sc_hd__buf_8
XFILLER_9_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput842 _593_/X vssd vssd vccd vccd la_oenb_core[96] sky130_fd_sc_hd__buf_8
Xoutput853 _319_/X vssd vssd vccd vccd mprj_adr_o_user[14] sky130_fd_sc_hd__buf_8
XFILLER_25_3533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput864 _329_/X vssd vssd vccd vccd mprj_adr_o_user[24] sky130_fd_sc_hd__buf_8
XFILLER_43_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput875 _310_/X vssd vssd vccd vccd mprj_adr_o_user[5] sky130_fd_sc_hd__buf_8
Xoutput886 _128_/Y vssd vssd vccd vccd mprj_dat_i_core[14] sky130_fd_sc_hd__buf_8
Xoutput897 _138_/Y vssd vssd vccd vccd mprj_dat_i_core[24] sky130_fd_sc_hd__buf_8
XFILLER_5_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_260_ _260_/A _260_/B vssd vssd vccd vccd _260_/X sky130_fd_sc_hd__and2_4
XPHY_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_191_ _191_/A _191_/B vssd vssd vccd vccd _191_/X sky130_fd_sc_hd__and2_2
XFILLER_26_4009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_irq_gates\[2\] user_irq_core[2] _293_/X vssd vssd vccd vccd _113_/A sky130_fd_sc_hd__nand2_1
XFILLER_43_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_440 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_451 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_462 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_527_ _527_/A _527_/B vssd vssd vccd vccd _527_/X sky130_fd_sc_hd__and2_4
XFILLER_15_3724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_473 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_484 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_495 _488_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_458_ _586_/A _458_/B _458_/C vssd vssd vccd vccd _458_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_389_ _517_/A _389_/B _389_/C vssd vssd vccd vccd _389_/X sky130_fd_sc_hd__and3b_4
XFILLER_12_1000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[98\] la_data_out_core[98] _261_/X vssd vssd vccd vccd _081_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_29_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_831 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2588 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4294 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4075 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput650 _021_/Y vssd vssd vccd vccd la_data_in_mprj[38] sky130_fd_sc_hd__buf_8
Xoutput661 _031_/Y vssd vssd vccd vccd la_data_in_mprj[48] sky130_fd_sc_hd__buf_8
XFILLER_9_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput672 _041_/Y vssd vssd vccd vccd la_data_in_mprj[58] sky130_fd_sc_hd__buf_8
XFILLER_25_3352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput683 _051_/Y vssd vssd vccd vccd la_data_in_mprj[68] sky130_fd_sc_hd__buf_8
XFILLER_44_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput694 _061_/Y vssd vssd vccd vccd la_data_in_mprj[78] sky130_fd_sc_hd__buf_8
XFILLER_8_1123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2695 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_146 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_312_ _312_/A _312_/B vssd vssd vccd vccd _312_/X sky130_fd_sc_hd__and2_4
XFILLER_51_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_243_ _243_/A _243_/B vssd vssd vccd vccd _243_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput18 la_data_out_mprj[112] vssd vssd vccd vccd _481_/C sky130_fd_sc_hd__buf_6
XFILLER_6_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput29 la_data_out_mprj[122] vssd vssd vccd vccd _491_/C sky130_fd_sc_hd__buf_4
XFILLER_10_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_174_ _174_/A _174_/B vssd vssd vccd vccd _174_/X sky130_fd_sc_hd__and2_4
XFILLER_13_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_270 _448_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_281 _449_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_292 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[13\] la_data_out_core[13] _176_/X vssd vssd vccd vccd _160_/A
+ sky130_fd_sc_hd__nand2_4
Xuser_wb_dat_gates\[26\] mprj_dat_i_user[26] _294_/X vssd vssd vccd vccd _140_/A sky130_fd_sc_hd__nand2_2
XFILLER_31_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1202 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[124\] la_data_out_core[124] _287_/X vssd vssd vccd vccd _107_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_42_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2309 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1608 _613_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_1619 _524_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput480 _484_/X vssd vssd vccd vccd la_data_in_core[115] sky130_fd_sc_hd__buf_8
Xoutput491 _494_/X vssd vssd vccd vccd la_data_in_core[125] sky130_fd_sc_hd__buf_8
XFILLER_40_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_226_ _226_/A _226_/B vssd vssd vccd vccd _226_/X sky130_fd_sc_hd__and2_2
XFILLER_10_4196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_157_ _157_/A vssd vssd vccd vccd _157_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_6_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_088_ _088_/A vssd vssd vccd vccd _088_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_4292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1824 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_4117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_3300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2919 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput208 la_iena_mprj[53] vssd vssd vccd vccd _216_/B sky130_fd_sc_hd__clkbuf_4
Xinput219 la_iena_mprj[63] vssd vssd vccd vccd _226_/B sky130_fd_sc_hd__buf_4
XFILLER_9_1251 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1076 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_296 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_011_ _011_/A vssd vssd vccd vccd _011_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2106 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2117 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2128 _193_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2139 _260_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1405 _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1416 _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1427 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1438 _370_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1449 _372_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_209_ _209_/A _209_/B vssd vssd vccd vccd _209_/X sky130_fd_sc_hd__and2_1
XFILLER_32_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_4332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[80\] la_data_out_core[80] _243_/X vssd vssd vccd vccd _063_/A
+ sky130_fd_sc_hd__nand2_8
XTAP_734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1950 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1961 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1972 _352_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1983 _367_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1994 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3460 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_560_ _560_/A _560_/B vssd vssd vccd vccd _560_/X sky130_fd_sc_hd__and2_4
XTAP_3858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_803 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_814 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_825 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_836 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_491_ _619_/A _491_/B _491_/C vssd vssd vccd vccd _491_/X sky130_fd_sc_hd__and3b_4
XANTENNA_847 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_858 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_869 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1202 _234_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1213 _249_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1224 _261_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1235 _266_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1246 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1257 _272_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1268 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1279 _275_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4022 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2470 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2481 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2492 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1780 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1791 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_612_ _612_/A _612_/B vssd vssd vccd vccd _612_/X sky130_fd_sc_hd__and2_4
XTAP_4378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_600 _510_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_611 _511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_543_ _543_/A _543_/B vssd vssd vccd vccd _543_/X sky130_fd_sc_hd__and2_4
XTAP_2932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_622 _519_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_633 _557_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_644 _567_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_655 _568_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_666 _574_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_474_ _602_/A _474_/B _474_/C vssd vssd vccd vccd _474_/X sky130_fd_sc_hd__and3b_4
XFILLER_15_3928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_677 _576_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_688 _579_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_699 _583_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1712 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1828 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1010 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1021 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1032 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1043 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1054 _172_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1065 _179_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1076 _182_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1087 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1098 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput380 la_oenb_mprj[93] vssd vssd vccd vccd _590_/A sky130_fd_sc_hd__buf_8
XFILLER_36_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput391 mprj_adr_o_core[12] vssd vssd vccd vccd _317_/B sky130_fd_sc_hd__buf_8
XFILLER_3_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[43\] la_data_out_core[43] _206_/X vssd vssd vccd vccd _026_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_4264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput810 _564_/X vssd vssd vccd vccd la_oenb_core[67] sky130_fd_sc_hd__buf_8
Xoutput821 _574_/X vssd vssd vccd vccd la_oenb_core[77] sky130_fd_sc_hd__buf_8
Xoutput832 _584_/X vssd vssd vccd vccd la_oenb_core[87] sky130_fd_sc_hd__buf_8
XFILLER_29_3681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput843 _594_/X vssd vssd vccd vccd la_oenb_core[97] sky130_fd_sc_hd__buf_8
XFILLER_9_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput854 _320_/X vssd vssd vccd vccd mprj_adr_o_user[15] sky130_fd_sc_hd__buf_8
Xoutput865 _330_/X vssd vssd vccd vccd mprj_adr_o_user[25] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[5\] la_data_out_core[5] _168_/X vssd vssd vccd vccd _152_/A
+ sky130_fd_sc_hd__nand2_2
Xoutput876 _311_/X vssd vssd vccd vccd mprj_adr_o_user[6] sky130_fd_sc_hd__buf_8
XFILLER_8_2039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput887 _129_/Y vssd vssd vccd vccd mprj_dat_i_core[15] sky130_fd_sc_hd__buf_8
XFILLER_5_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput898 _139_/Y vssd vssd vccd vccd mprj_dat_i_core[25] sky130_fd_sc_hd__buf_8
XFILLER_25_3589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_190_ _190_/A _190_/B vssd vssd vccd vccd _190_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2194 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_430 _480_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_441 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_452 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_526_ _526_/A _526_/B vssd vssd vccd vccd _526_/X sky130_fd_sc_hd__and2_4
XFILLER_50_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_463 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_474 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_485 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_496 _488_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_457_ _585_/A _457_/B _457_/C vssd vssd vccd vccd _457_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_388_ _516_/A _388_/B _388_/C vssd vssd vccd vccd _388_/X sky130_fd_sc_hd__and3b_4
XFILLER_48_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_4526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput640 _012_/Y vssd vssd vccd vccd la_data_in_mprj[29] sky130_fd_sc_hd__buf_8
XFILLER_25_3320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput651 _022_/Y vssd vssd vccd vccd la_data_in_mprj[39] sky130_fd_sc_hd__buf_8
XFILLER_25_4087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput662 _032_/Y vssd vssd vccd vccd la_data_in_mprj[49] sky130_fd_sc_hd__buf_8
Xoutput673 _042_/Y vssd vssd vccd vccd la_data_in_mprj[59] sky130_fd_sc_hd__buf_8
Xoutput684 _052_/Y vssd vssd vccd vccd la_data_in_mprj[69] sky130_fd_sc_hd__buf_8
XFILLER_25_3364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput695 _062_/Y vssd vssd vccd vccd la_data_in_mprj[79] sky130_fd_sc_hd__buf_8
XFILLER_5_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_311_ _311_/A _311_/B vssd vssd vccd vccd _311_/X sky130_fd_sc_hd__and2_4
XFILLER_14_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_242_ _242_/A _242_/B vssd vssd vccd vccd _242_/X sky130_fd_sc_hd__and2_4
XFILLER_52_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput19 la_data_out_mprj[113] vssd vssd vccd vccd _482_/C sky130_fd_sc_hd__buf_4
XFILLER_7_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_173_ _173_/A _173_/B vssd vssd vccd vccd _173_/X sky130_fd_sc_hd__and2_4
XFILLER_32_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_260 _445_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_271 _448_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_509_ _509_/A _509_/B vssd vssd vccd vccd _509_/X sky130_fd_sc_hd__and2_4
XANTENNA_282 _449_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_293 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3290 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[19\] mprj_dat_i_user[19] _294_/X vssd vssd vccd vccd _133_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1214 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[117\] la_data_out_core[117] _280_/X vssd vssd vccd vccd _100_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_0_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput470 _475_/X vssd vssd vccd vccd la_data_in_core[106] sky130_fd_sc_hd__buf_8
XFILLER_44_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1609 _613_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput481 _485_/X vssd vssd vccd vccd la_data_in_core[116] sky130_fd_sc_hd__buf_8
Xoutput492 _495_/X vssd vssd vccd vccd la_data_in_core[126] sky130_fd_sc_hd__buf_8
XFILLER_40_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_225_ _225_/A _225_/B vssd vssd vccd vccd _225_/X sky130_fd_sc_hd__and2_4
XFILLER_11_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_156_ _156_/A vssd vssd vccd vccd _156_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_087_ _087_/A vssd vssd vccd vccd _087_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput209 la_iena_mprj[54] vssd vssd vccd vccd _217_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_010_ _010_/A vssd vssd vccd vccd _010_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2107 _538_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2118 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2129 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1406 _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1417 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1428 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1439 _370_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_208_ _208_/A _208_/B vssd vssd vccd vccd _208_/X sky130_fd_sc_hd__and2_1
XFILLER_45_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_139_ _139_/A vssd vssd vccd vccd _139_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_3_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2630 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1940 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1951 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[73\] la_data_out_core[73] _236_/X vssd vssd vccd vccd _056_/A
+ sky130_fd_sc_hd__nand2_8
XTAP_779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1962 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1973 _353_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1984 _342_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1995 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2782 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1947 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1688 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4488 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_804 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_815 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_826 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_837 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_490_ _618_/A _490_/B _490_/C vssd vssd vccd vccd _490_/X sky130_fd_sc_hd__and3b_4
XFILLER_2_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_848 _613_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_859 _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1203 _236_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1214 _250_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1225 _262_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1236 _268_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1247 _270_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1258 _272_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1269 _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4034 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3727 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4174 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2460 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3440 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2471 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2482 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2493 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1770 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1781 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1792 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2510 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1463 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_611_ _611_/A _611_/B vssd vssd vccd vccd _611_/X sky130_fd_sc_hd__and2_4
XTAP_4368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_601 _510_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_612 _511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_542_ _542_/A _542_/B vssd vssd vccd vccd _542_/X sky130_fd_sc_hd__and2_4
XTAP_3678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_623 _519_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_634 _558_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_645 _567_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_656 _568_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_473_ _601_/A _473_/B _473_/C vssd vssd vccd vccd _473_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_4321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_667 _574_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_678 _576_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_689 _580_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1702 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1000 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1011 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1022 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1033 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1044 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4358 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1055 _173_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1066 _180_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1077 _182_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1088 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_1099 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput370 la_oenb_mprj[84] vssd vssd vccd vccd _581_/A sky130_fd_sc_hd__buf_8
Xinput381 la_oenb_mprj[94] vssd vssd vccd vccd _591_/A sky130_fd_sc_hd__buf_8
XFILLER_7_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput392 mprj_adr_o_core[13] vssd vssd vccd vccd _318_/B sky130_fd_sc_hd__buf_8
XFILLER_36_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[36\] la_data_out_core[36] _199_/X vssd vssd vccd vccd _019_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput800 _555_/X vssd vssd vccd vccd la_oenb_core[58] sky130_fd_sc_hd__buf_8
XFILLER_29_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput811 _565_/X vssd vssd vccd vccd la_oenb_core[68] sky130_fd_sc_hd__buf_8
XFILLER_9_3732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput822 _575_/X vssd vssd vccd vccd la_oenb_core[78] sky130_fd_sc_hd__buf_8
Xoutput833 _585_/X vssd vssd vccd vccd la_oenb_core[88] sky130_fd_sc_hd__buf_8
Xoutput844 _595_/X vssd vssd vccd vccd la_oenb_core[98] sky130_fd_sc_hd__buf_8
XFILLER_8_2007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput855 _321_/X vssd vssd vccd vccd mprj_adr_o_user[16] sky130_fd_sc_hd__buf_8
XFILLER_42_4550 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput866 _331_/X vssd vssd vccd vccd mprj_adr_o_user[26] sky130_fd_sc_hd__buf_8
XFILLER_29_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput877 _312_/X vssd vssd vccd vccd mprj_adr_o_user[7] sky130_fd_sc_hd__buf_8
XFILLER_3_4021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput888 _130_/Y vssd vssd vccd vccd mprj_dat_i_core[16] sky130_fd_sc_hd__buf_8
XFILLER_28_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput899 _140_/Y vssd vssd vccd vccd mprj_dat_i_core[26] sky130_fd_sc_hd__buf_8
XFILLER_3_4054 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2290 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_420 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_431 _482_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_442 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_525_ _525_/A _525_/B vssd vssd vccd vccd _525_/X sky130_fd_sc_hd__and2_4
XTAP_2752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_453 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_464 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_475 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_486 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_497 _488_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_456_ _584_/A _456_/B _456_/C vssd vssd vccd vccd _456_/X sky130_fd_sc_hd__and3b_4
XFILLER_41_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_387_ _515_/A _387_/B _387_/C vssd vssd vccd vccd _387_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3811 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3708 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1576 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3432 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput630 _148_/Y vssd vssd vccd vccd la_data_in_mprj[1] sky130_fd_sc_hd__buf_8
XFILLER_27_2929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput641 _149_/Y vssd vssd vccd vccd la_data_in_mprj[2] sky130_fd_sc_hd__buf_8
Xoutput652 _150_/Y vssd vssd vccd vccd la_data_in_mprj[3] sky130_fd_sc_hd__buf_8
XFILLER_25_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput663 _151_/Y vssd vssd vccd vccd la_data_in_mprj[4] sky130_fd_sc_hd__buf_8
XFILLER_9_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput674 _152_/Y vssd vssd vccd vccd la_data_in_mprj[5] sky130_fd_sc_hd__buf_8
Xoutput685 _153_/Y vssd vssd vccd vccd la_data_in_mprj[6] sky130_fd_sc_hd__buf_8
Xoutput696 _154_/Y vssd vssd vccd vccd la_data_in_mprj[7] sky130_fd_sc_hd__buf_8
XFILLER_5_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ _310_/A _310_/B vssd vssd vccd vccd _310_/X sky130_fd_sc_hd__and2_4
XFILLER_42_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_241_ _241_/A _241_/B vssd vssd vccd vccd _241_/X sky130_fd_sc_hd__and2_4
XFILLER_51_991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3792 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_172_ _172_/A _172_/B vssd vssd vccd vccd _172_/X sky130_fd_sc_hd__and2_4
XFILLER_49_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_498 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_250 _440_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_261 _445_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_508_ _508_/A _508_/B vssd vssd vccd vccd _508_/X sky130_fd_sc_hd__and2_4
XANTENNA_272 _448_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_283 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_294 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_439_ _567_/A _439_/B _439_/C vssd vssd vccd vccd _439_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1488 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_788 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_2207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput471 _476_/X vssd vssd vccd vccd la_data_in_core[107] sky130_fd_sc_hd__buf_8
Xoutput482 _486_/X vssd vssd vccd vccd la_data_in_core[117] sky130_fd_sc_hd__buf_8
Xoutput493 _496_/X vssd vssd vccd vccd la_data_in_core[127] sky130_fd_sc_hd__buf_8
XFILLER_40_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1990 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1707 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_224_ _224_/A _224_/B vssd vssd vccd vccd _224_/X sky130_fd_sc_hd__and2_2
XFILLER_7_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_155_ _155_/A vssd vssd vccd vccd _155_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_13_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[1\] mprj_dat_i_user[1] _294_/X vssd vssd vccd vccd _115_/A sky130_fd_sc_hd__nand2_1
XFILLER_10_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_086_ _086_/A vssd vssd vccd vccd _086_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[31\] mprj_dat_i_user[31] _294_/X vssd vssd vccd vccd _145_/A sky130_fd_sc_hd__nand2_2
XFILLER_21_438 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2108 _539_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2119 _167_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1407 _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1418 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1429 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_207_ _207_/A _207_/B vssd vssd vccd vccd _207_/X sky130_fd_sc_hd__and2_1
XFILLER_50_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_138_ _138_/A vssd vssd vccd vccd _138_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_28_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_069_ _069_/A vssd vssd vccd vccd _069_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_28_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2620 _362_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2631 _362_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1930 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1941 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1952 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1963 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1974 _354_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[66\] la_data_out_core[66] _229_/X vssd vssd vccd vccd _049_/A
+ sky130_fd_sc_hd__nand2_4
XANTENNA_1985 _345_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1996 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_805 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_816 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_827 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_838 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_849 _613_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1204 _239_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1215 _251_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1226 _262_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1237 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1248 _270_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1259 _272_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4458 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4046 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1066 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3739 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2450 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2461 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4186 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2472 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2483 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2494 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1760 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1771 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1782 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1793 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1723 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3468 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_610_ _610_/A _610_/B vssd vssd vccd vccd _610_/X sky130_fd_sc_hd__and2_4
XTAP_4358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_602 _510_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_541_ _541_/A _541_/B vssd vssd vccd vccd _541_/X sky130_fd_sc_hd__and2_4
XTAP_2912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_613 _511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_624 _520_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_635 _559_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_646 _568_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_472_ _600_/A _472_/B _472_/C vssd vssd vccd vccd _472_/X sky130_fd_sc_hd__and3b_4
XANTENNA_657 _569_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_668 _574_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_679 _576_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_4393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1001 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1012 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3822 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1023 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1034 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1045 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1056 _174_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1067 _181_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1078 _182_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1089 _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput360 la_oenb_mprj[75] vssd vssd vccd vccd _572_/A sky130_fd_sc_hd__buf_8
XFILLER_42_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput371 la_oenb_mprj[85] vssd vssd vccd vccd _582_/A sky130_fd_sc_hd__buf_8
XFILLER_23_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput382 la_oenb_mprj[95] vssd vssd vccd vccd _592_/A sky130_fd_sc_hd__buf_8
Xinput393 mprj_adr_o_core[14] vssd vssd vccd vccd _319_/B sky130_fd_sc_hd__buf_8
XFILLER_36_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[29\] la_data_out_core[29] _192_/X vssd vssd vccd vccd _012_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_31_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2018 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput801 _556_/X vssd vssd vccd vccd la_oenb_core[59] sky130_fd_sc_hd__buf_8
Xoutput812 _566_/X vssd vssd vccd vccd la_oenb_core[69] sky130_fd_sc_hd__buf_8
Xoutput823 _576_/X vssd vssd vccd vccd la_oenb_core[79] sky130_fd_sc_hd__buf_8
XFILLER_9_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput834 _586_/X vssd vssd vccd vccd la_oenb_core[89] sky130_fd_sc_hd__buf_8
Xoutput845 _596_/X vssd vssd vccd vccd la_oenb_core[99] sky130_fd_sc_hd__buf_8
Xoutput856 _322_/X vssd vssd vccd vccd mprj_adr_o_user[17] sky130_fd_sc_hd__buf_8
XFILLER_8_2019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput867 _332_/X vssd vssd vccd vccd mprj_adr_o_user[27] sky130_fd_sc_hd__buf_8
XFILLER_42_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput878 _313_/X vssd vssd vccd vccd mprj_adr_o_user[8] sky130_fd_sc_hd__buf_8
XFILLER_47_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput889 _131_/Y vssd vssd vccd vccd mprj_dat_i_core[17] sky130_fd_sc_hd__buf_8
XTAP_330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4066 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_2280 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2291 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1590 _439_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_102 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_410 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_421 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_524_ _524_/A _524_/B vssd vssd vccd vccd _524_/X sky130_fd_sc_hd__and2_4
XTAP_2742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_432 _482_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_443 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_454 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_465 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_476 _486_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_455_ _583_/A _455_/B _455_/C vssd vssd vccd vccd _455_/X sky130_fd_sc_hd__and3b_4
XTAP_2797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_487 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_498 _488_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3440 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_386_ _514_/A _386_/B _386_/C vssd vssd vccd vccd _386_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1150 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3823 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1588 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput190 la_iena_mprj[37] vssd vssd vccd vccd _200_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput620 _109_/Y vssd vssd vccd vccd la_data_in_mprj[126] sky130_fd_sc_hd__buf_8
XFILLER_47_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_4128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput631 _003_/Y vssd vssd vccd vccd la_data_in_mprj[20] sky130_fd_sc_hd__buf_8
XFILLER_9_3552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput642 _013_/Y vssd vssd vccd vccd la_data_in_mprj[30] sky130_fd_sc_hd__buf_8
XFILLER_43_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput653 _023_/Y vssd vssd vccd vccd la_data_in_mprj[40] sky130_fd_sc_hd__buf_8
XFILLER_47_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput664 _033_/Y vssd vssd vccd vccd la_data_in_mprj[50] sky130_fd_sc_hd__buf_8
XFILLER_28_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput675 _043_/Y vssd vssd vccd vccd la_data_in_mprj[60] sky130_fd_sc_hd__buf_8
XFILLER_9_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput686 _053_/Y vssd vssd vccd vccd la_data_in_mprj[70] sky130_fd_sc_hd__buf_8
Xoutput697 _063_/Y vssd vssd vccd vccd la_data_in_mprj[80] sky130_fd_sc_hd__buf_8
XFILLER_28_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_240_ _240_/A _240_/B vssd vssd vccd vccd _240_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_171_ _171_/A _171_/B vssd vssd vccd vccd _171_/X sky130_fd_sc_hd__and2_4
XFILLER_32_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1080 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_irq_gates\[0\] user_irq_core[0] _291_/X vssd vssd vccd vccd _111_/A sky130_fd_sc_hd__nand2_1
XFILLER_43_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1671 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_240 _435_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 _440_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_507_ _507_/A _507_/B vssd vssd vccd vccd _507_/X sky130_fd_sc_hd__and2_4
XANTENNA_262 _445_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_273 _448_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4550 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_284 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_295 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_438_ _566_/A _438_/B _438_/C vssd vssd vccd vccd _438_/X sky130_fd_sc_hd__and3b_4
XFILLER_18_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_369_ _497_/A _369_/B _369_/C vssd vssd vccd vccd _369_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[96\] la_data_out_core[96] _259_/X vssd vssd vccd vccd _079_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_6_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2147 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_2219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput472 _477_/X vssd vssd vccd vccd la_data_in_core[108] sky130_fd_sc_hd__buf_8
XFILLER_47_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput483 _487_/X vssd vssd vccd vccd la_data_in_core[118] sky130_fd_sc_hd__buf_8
Xoutput494 _381_/X vssd vssd vccd vccd la_data_in_core[12] sky130_fd_sc_hd__buf_8
XFILLER_5_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_296 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_223_ _223_/A _223_/B vssd vssd vccd vccd _223_/X sky130_fd_sc_hd__and2_2
XFILLER_50_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_154_ _154_/A vssd vssd vccd vccd _154_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_085_ _085_/A vssd vssd vccd vccd _085_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_49_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[11\] la_data_out_core[11] _174_/X vssd vssd vccd vccd _158_/A
+ sky130_fd_sc_hd__nand2_4
Xuser_wb_dat_gates\[24\] mprj_dat_i_user[24] _294_/X vssd vssd vccd vccd _138_/A sky130_fd_sc_hd__nand2_2
XFILLER_50_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[122\] la_data_out_core[122] _285_/X vssd vssd vccd vccd _105_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_29_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2109 _546_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1408 _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1419 _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_206_ _206_/A _206_/B vssd vssd vccd vccd _206_/X sky130_fd_sc_hd__and2_1
X_137_ _137_/A vssd vssd vccd vccd _137_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_068_ _068_/A vssd vssd vccd vccd _068_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2610 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2621 la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1920 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1931 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1942 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1953 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1964 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1975 _355_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1986 _346_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1997 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[59\] la_data_out_core[59] _222_/X vssd vssd vccd vccd _042_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2708 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_806 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1858 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_817 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_828 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_839 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1205 _240_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1216 _252_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1227 _262_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1238 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1249 _271_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3736 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3460 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1056 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2440 _454_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2451 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2462 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2473 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2484 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1750 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2495 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1761 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1772 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1783 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1794 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2458 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_906 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_540_ _540_/A _540_/B vssd vssd vccd vccd _540_/X sky130_fd_sc_hd__and2_4
XTAP_2913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_603 _511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_614 _511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_625 _521_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_840 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_636 _321_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_471_ _599_/A _471_/B _471_/C vssd vssd vccd vccd _471_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_647 _568_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_658 _569_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_669 _574_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1002 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1013 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1024 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1035 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1046 _167_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1057 _175_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1068 _182_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1079 _329_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput350 la_oenb_mprj[66] vssd vssd vccd vccd _563_/A sky130_fd_sc_hd__buf_6
Xinput361 la_oenb_mprj[76] vssd vssd vccd vccd _573_/A sky130_fd_sc_hd__buf_8
Xinput372 la_oenb_mprj[86] vssd vssd vccd vccd _583_/A sky130_fd_sc_hd__buf_8
XFILLER_40_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput383 la_oenb_mprj[96] vssd vssd vccd vccd _593_/A sky130_fd_sc_hd__buf_6
XFILLER_48_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput394 mprj_adr_o_core[15] vssd vssd vccd vccd _320_/B sky130_fd_sc_hd__buf_8
XFILLER_23_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput802 _502_/X vssd vssd vccd vccd la_oenb_core[5] sky130_fd_sc_hd__buf_8
Xoutput813 _503_/X vssd vssd vccd vccd la_oenb_core[6] sky130_fd_sc_hd__buf_8
Xoutput824 _504_/X vssd vssd vccd vccd la_oenb_core[7] sky130_fd_sc_hd__buf_8
Xoutput835 _505_/X vssd vssd vccd vccd la_oenb_core[8] sky130_fd_sc_hd__buf_8
XFILLER_6_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput846 _506_/X vssd vssd vccd vccd la_oenb_core[9] sky130_fd_sc_hd__buf_8
XFILLER_29_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput857 _323_/X vssd vssd vccd vccd mprj_adr_o_user[18] sky130_fd_sc_hd__buf_8
XFILLER_7_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput868 _333_/X vssd vssd vccd vccd mprj_adr_o_user[28] sky130_fd_sc_hd__buf_8
Xoutput879 _314_/X vssd vssd vccd vccd mprj_adr_o_user[9] sky130_fd_sc_hd__buf_8
XFILLER_25_3559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2847 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2270 _367_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2281 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2292 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1580 _296_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1591 _445_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_114 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_400 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_411 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_422 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_523_ _523_/A _523_/B vssd vssd vccd vccd _523_/X sky130_fd_sc_hd__and2_4
XTAP_3488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_433 _482_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_444 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_455 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_466 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_477 _486_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_454_ _582_/A _454_/B _454_/C vssd vssd vccd vccd _454_/X sky130_fd_sc_hd__and3b_4
XANTENNA_488 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_499 _488_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_385_ _513_/A _385_/B _385_/C vssd vssd vccd vccd _385_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_3452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1162 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput180 la_iena_mprj[28] vssd vssd vccd vccd _191_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput191 la_iena_mprj[38] vssd vssd vccd vccd _201_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[41\] la_data_out_core[41] _204_/X vssd vssd vccd vccd _024_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3352 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput610 _100_/Y vssd vssd vccd vccd la_data_in_mprj[117] sky130_fd_sc_hd__buf_8
Xoutput621 _110_/Y vssd vssd vccd vccd la_data_in_mprj[127] sky130_fd_sc_hd__buf_8
Xoutput632 _004_/Y vssd vssd vccd vccd la_data_in_mprj[21] sky130_fd_sc_hd__buf_8
XFILLER_47_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput643 _014_/Y vssd vssd vccd vccd la_data_in_mprj[31] sky130_fd_sc_hd__buf_8
XFILLER_9_3564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput654 _024_/Y vssd vssd vccd vccd la_data_in_mprj[41] sky130_fd_sc_hd__buf_8
XFILLER_5_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput665 _034_/Y vssd vssd vccd vccd la_data_in_mprj[51] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[3\] la_data_out_core[3] _166_/X vssd vssd vccd vccd _150_/A
+ sky130_fd_sc_hd__nand2_1
Xoutput676 _044_/Y vssd vssd vccd vccd la_data_in_mprj[61] sky130_fd_sc_hd__buf_8
XFILLER_28_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput687 _054_/Y vssd vssd vccd vccd la_data_in_mprj[71] sky130_fd_sc_hd__buf_8
Xoutput698 _064_/Y vssd vssd vccd vccd la_data_in_mprj[81] sky130_fd_sc_hd__buf_8
XFILLER_42_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_170_ _170_/A _170_/B vssd vssd vccd vccd _170_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4400 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1683 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_230 _434_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_241 _435_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_506_ _506_/A _506_/B vssd vssd vccd vccd _506_/X sky130_fd_sc_hd__and2_4
XANTENNA_252 _441_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_263 _445_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_274 _448_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_296 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_437_ _565_/A _437_/B _437_/C vssd vssd vccd vccd _437_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_150 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_368_ _368_/A _368_/B vssd vssd vccd vccd _368_/X sky130_fd_sc_hd__and2_4
XFILLER_31_2147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_299_ _299_/A _299_/B vssd vssd vccd vccd _299_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3643 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[89\] la_data_out_core[89] _252_/X vssd vssd vccd vccd _072_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_3687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput473 _478_/X vssd vssd vccd vccd la_data_in_core[109] sky130_fd_sc_hd__buf_8
Xoutput484 _488_/X vssd vssd vccd vccd la_data_in_core[119] sky130_fd_sc_hd__buf_8
XFILLER_43_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput495 _382_/X vssd vssd vccd vccd la_data_in_core[13] sky130_fd_sc_hd__buf_8
XFILLER_5_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_222_ _222_/A _222_/B vssd vssd vccd vccd _222_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_153_ _153_/A vssd vssd vccd vccd _153_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_084_ _084_/A vssd vssd vccd vccd _084_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[17\] mprj_dat_i_user[17] _294_/X vssd vssd vccd vccd _131_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_1806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1828 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[115\] la_data_out_core[115] _278_/X vssd vssd vccd vccd _098_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_20_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1409 _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2490 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_205_ _205_/A _205_/B vssd vssd vccd vccd _205_/X sky130_fd_sc_hd__and2_2
XFILLER_12_996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_136_ _136_/A vssd vssd vccd vccd _136_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_067_ _067_/A vssd vssd vccd vccd _067_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_1850 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2600 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_2611 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1894 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2622 _305_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1910 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1921 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1932 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1943 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1954 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1965 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1976 _357_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1987 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1998 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_807 _606_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_818 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_829 _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1206 _242_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1217 _336_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1228 _262_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1239 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_119_ _119_/A vssd vssd vccd vccd _119_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_2108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2430 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2441 _189_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2452 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2463 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2474 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1740 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2485 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[71\] la_data_out_core[71] _234_/X vssd vssd vccd vccd _054_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1751 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2496 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1762 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1773 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1784 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_1795 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1747 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1634 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_604 _511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_615 _513_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_626 _521_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_470_ _598_/A _470_/B _470_/C vssd vssd vccd vccd _470_/X sky130_fd_sc_hd__and3b_4
XFILLER_26_852 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_637 _565_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_648 _568_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_659 _569_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3960 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1003 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1014 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_1025 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1036 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1047 _167_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1058 _176_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3879 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1069 _182_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput340 la_oenb_mprj[57] vssd vssd vccd vccd _554_/A sky130_fd_sc_hd__buf_4
XFILLER_20_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput351 la_oenb_mprj[67] vssd vssd vccd vccd _564_/A sky130_fd_sc_hd__buf_6
Xinput362 la_oenb_mprj[77] vssd vssd vccd vccd _574_/A sky130_fd_sc_hd__buf_8
XFILLER_49_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput373 la_oenb_mprj[87] vssd vssd vccd vccd _584_/A sky130_fd_sc_hd__buf_8
XFILLER_2_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput384 la_oenb_mprj[97] vssd vssd vccd vccd _594_/A sky130_fd_sc_hd__buf_6
Xinput395 mprj_adr_o_core[16] vssd vssd vccd vccd _321_/B sky130_fd_sc_hd__buf_8
XFILLER_53_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_599_ _599_/A _599_/B vssd vssd vccd vccd _599_/X sky130_fd_sc_hd__and2_4
XFILLER_43_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput803 _557_/X vssd vssd vccd vccd la_oenb_core[60] sky130_fd_sc_hd__buf_8
Xoutput814 _567_/X vssd vssd vccd vccd la_oenb_core[70] sky130_fd_sc_hd__buf_8
Xoutput825 _577_/X vssd vssd vccd vccd la_oenb_core[80] sky130_fd_sc_hd__buf_8
XFILLER_47_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput836 _587_/X vssd vssd vccd vccd la_oenb_core[90] sky130_fd_sc_hd__buf_8
XFILLER_29_3685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput847 _146_/Y vssd vssd vccd vccd mprj_ack_i_core sky130_fd_sc_hd__buf_8
XFILLER_25_3527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput858 _324_/X vssd vssd vccd vccd mprj_adr_o_user[19] sky130_fd_sc_hd__buf_8
XFILLER_3_4013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput869 _334_/X vssd vssd vccd vccd mprj_adr_o_user[29] sky130_fd_sc_hd__buf_8
XFILLER_47_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2260 _302_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2271 _368_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2282 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2293 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1570 _296_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1581 _296_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_1592 _450_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_126 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_401 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_412 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_522_ _522_/A _522_/B vssd vssd vccd vccd _522_/X sky130_fd_sc_hd__and2_4
XTAP_2722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_423 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_434 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_445 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_456 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_467 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_453_ _581_/A _453_/B _453_/C vssd vssd vccd vccd _453_/X sky130_fd_sc_hd__and3b_4
XTAP_2777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_478 _486_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_489 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_384_ _512_/A _384_/B _384_/C vssd vssd vccd vccd _384_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1134 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput170 la_iena_mprj[19] vssd vssd vccd vccd _182_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_49_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput181 la_iena_mprj[29] vssd vssd vccd vccd _192_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_36_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput192 la_iena_mprj[39] vssd vssd vccd vccd _202_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_4508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[34\] la_data_out_core[34] _197_/X vssd vssd vccd vccd _017_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_990 _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput600 _091_/Y vssd vssd vccd vccd la_data_in_mprj[108] sky130_fd_sc_hd__buf_8
XFILLER_5_4108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput611 _101_/Y vssd vssd vccd vccd la_data_in_mprj[118] sky130_fd_sc_hd__buf_8
Xoutput622 _159_/Y vssd vssd vccd vccd la_data_in_mprj[12] sky130_fd_sc_hd__buf_8
XFILLER_29_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput633 _005_/Y vssd vssd vccd vccd la_data_in_mprj[22] sky130_fd_sc_hd__buf_8
XFILLER_44_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput644 _015_/Y vssd vssd vccd vccd la_data_in_mprj[32] sky130_fd_sc_hd__buf_8
Xoutput655 _025_/Y vssd vssd vccd vccd la_data_in_mprj[42] sky130_fd_sc_hd__buf_8
XFILLER_9_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput666 _035_/Y vssd vssd vccd vccd la_data_in_mprj[52] sky130_fd_sc_hd__buf_8
XFILLER_29_2770 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput677 _045_/Y vssd vssd vccd vccd la_data_in_mprj[62] sky130_fd_sc_hd__buf_8
Xoutput688 _055_/Y vssd vssd vccd vccd la_data_in_mprj[72] sky130_fd_sc_hd__buf_8
XFILLER_25_3379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput699 _065_/Y vssd vssd vccd vccd la_data_in_mprj[82] sky130_fd_sc_hd__buf_8
XFILLER_42_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2090 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3740 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_220 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 _434_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_505_ _505_/A _505_/B vssd vssd vccd vccd _505_/X sky130_fd_sc_hd__and2_4
XTAP_2552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_242 _440_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_253 _441_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_264 _447_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_275 _448_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_286 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_436_ _564_/A _436_/B _436_/C vssd vssd vccd vccd _436_/X sky130_fd_sc_hd__and3b_4
XTAP_1862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_297 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_367_ _367_/A _367_/B vssd vssd vccd vccd _367_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_298_ _298_/A _298_/B vssd vssd vccd vccd _298_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3699 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2482 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2707 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput463 _369_/X vssd vssd vccd vccd la_data_in_core[0] sky130_fd_sc_hd__buf_8
Xoutput474 _379_/X vssd vssd vccd vccd la_data_in_core[10] sky130_fd_sc_hd__buf_8
Xoutput485 _380_/X vssd vssd vccd vccd la_data_in_core[11] sky130_fd_sc_hd__buf_8
Xoutput496 _383_/X vssd vssd vccd vccd la_data_in_core[14] sky130_fd_sc_hd__buf_8
XFILLER_9_2683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_221_ _221_/A _221_/B vssd vssd vccd vccd _221_/X sky130_fd_sc_hd__and2_2
XFILLER_14_3570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_152_ _152_/A vssd vssd vccd vccd _152_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_49_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1122 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_083_ _083_/A vssd vssd vccd vccd _083_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_30_2181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_419_ _547_/A _419_/B _419_/C vssd vssd vccd vccd _419_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3463 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2795 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[108\] la_data_out_core[108] _271_/X vssd vssd vccd vccd _091_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_0_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_204_ _204_/A _204_/B vssd vssd vccd vccd _204_/X sky130_fd_sc_hd__and2_2
XFILLER_12_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_135_ _135_/A vssd vssd vccd vccd _135_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_066_ _066_/A vssd vssd vccd vccd _066_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_1840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_4462 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2601 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2612 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2623 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3783 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1900 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1911 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1922 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1933 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1944 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1955 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1966 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1977 _358_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1988 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1999 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1918 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_808 _607_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_819 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1207 _244_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1218 _253_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1229 _262_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_82 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4502 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_118_ _118_/A vssd vssd vccd vccd _118_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_049_ _049_/A vssd vssd vccd vccd _049_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_29_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_2420 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2431 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2442 _362_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2453 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2464 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1730 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2475 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1741 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2486 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1752 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2497 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1763 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1774 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1785 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1796 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[64\] la_data_out_core[64] _227_/X vssd vssd vccd vccd _047_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_21_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_605 _511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_616 _514_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_627 _524_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_638 _565_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_649 _568_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1990 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3731 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1004 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3742 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1015 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1026 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1037 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1048 _167_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1059 _176_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput330 la_oenb_mprj[48] vssd vssd vccd vccd _545_/A sky130_fd_sc_hd__buf_6
XFILLER_0_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput341 la_oenb_mprj[58] vssd vssd vccd vccd _555_/A sky130_fd_sc_hd__buf_6
XFILLER_48_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput352 la_oenb_mprj[68] vssd vssd vccd vccd _565_/A sky130_fd_sc_hd__buf_8
Xinput363 la_oenb_mprj[78] vssd vssd vccd vccd _575_/A sky130_fd_sc_hd__buf_8
Xinput374 la_oenb_mprj[88] vssd vssd vccd vccd _585_/A sky130_fd_sc_hd__buf_8
XFILLER_29_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput385 la_oenb_mprj[98] vssd vssd vccd vccd _595_/A sky130_fd_sc_hd__buf_6
XFILLER_48_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput396 mprj_adr_o_core[17] vssd vssd vccd vccd _322_/B sky130_fd_sc_hd__buf_8
XFILLER_2_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_598_ _598_/A _598_/B vssd vssd vccd vccd _598_/X sky130_fd_sc_hd__and2_4
XFILLER_34_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1 _083_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput804 _558_/X vssd vssd vccd vccd la_oenb_core[61] sky130_fd_sc_hd__buf_8
XFILLER_29_3653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput815 _568_/X vssd vssd vccd vccd la_oenb_core[71] sky130_fd_sc_hd__buf_8
XFILLER_29_3664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput826 _578_/X vssd vssd vccd vccd la_oenb_core[81] sky130_fd_sc_hd__buf_8
Xoutput837 _588_/X vssd vssd vccd vccd la_oenb_core[91] sky130_fd_sc_hd__buf_8
XFILLER_6_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput848 _305_/X vssd vssd vccd vccd mprj_adr_o_user[0] sky130_fd_sc_hd__buf_8
XFILLER_28_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput859 _306_/X vssd vssd vccd vccd mprj_adr_o_user[1] sky130_fd_sc_hd__buf_8
XFILLER_25_2805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_4565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2250 _523_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2261 _302_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2272 _345_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2283 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2294 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1560 _391_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1571 _296_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1582 _296_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1593 _457_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_738 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1410 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_402 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_521_ _521_/A _521_/B vssd vssd vccd vccd _521_/X sky130_fd_sc_hd__and2_4
XTAP_2723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_413 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_424 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_435 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_446 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_457 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_452_ _580_/A _452_/B _452_/C vssd vssd vccd vccd _452_/X sky130_fd_sc_hd__and3b_4
XFILLER_19_3888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_468 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_479 _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_383_ _511_/A _383_/B _383_/C vssd vssd vccd vccd _383_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput160 la_iena_mprj[125] vssd vssd vccd vccd _288_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1146 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput171 la_iena_mprj[1] vssd vssd vccd vccd _164_/B sky130_fd_sc_hd__clkbuf_4
Xinput182 la_iena_mprj[2] vssd vssd vccd vccd _165_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_49_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput193 la_iena_mprj[3] vssd vssd vccd vccd _166_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_4022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_980 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[27\] la_data_out_core[27] _190_/X vssd vssd vccd vccd _010_/A
+ sky130_fd_sc_hd__nand2_2
XANTENNA_991 _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput601 _092_/Y vssd vssd vccd vccd la_data_in_mprj[109] sky130_fd_sc_hd__buf_8
XFILLER_25_4037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput612 _102_/Y vssd vssd vccd vccd la_data_in_mprj[119] sky130_fd_sc_hd__buf_8
Xoutput623 _160_/Y vssd vssd vccd vccd la_data_in_mprj[13] sky130_fd_sc_hd__buf_8
Xoutput634 _006_/Y vssd vssd vccd vccd la_data_in_mprj[23] sky130_fd_sc_hd__buf_8
Xoutput645 _016_/Y vssd vssd vccd vccd la_data_in_mprj[33] sky130_fd_sc_hd__buf_8
XFILLER_47_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput656 _026_/Y vssd vssd vccd vccd la_data_in_mprj[43] sky130_fd_sc_hd__buf_8
Xoutput667 _036_/Y vssd vssd vccd vccd la_data_in_mprj[53] sky130_fd_sc_hd__buf_8
XFILLER_29_2782 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput678 _046_/Y vssd vssd vccd vccd la_data_in_mprj[63] sky130_fd_sc_hd__buf_8
Xoutput689 _056_/Y vssd vssd vccd vccd la_data_in_mprj[73] sky130_fd_sc_hd__buf_8
XFILLER_42_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2080 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2091 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1390 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1684 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1072 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_221 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_232 _434_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_504_ _504_/A _504_/B vssd vssd vccd vccd _504_/X sky130_fd_sc_hd__and2_4
XFILLER_33_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_243 _440_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_254 _441_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 _447_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_276 _448_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_435_ _563_/A _435_/B _435_/C vssd vssd vccd vccd _435_/X sky130_fd_sc_hd__and3b_4
XANTENNA_287 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_298 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_366_ _366_/A _366_/B vssd vssd vccd vccd _366_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_297_ _297_/A _297_/B vssd vssd vccd vccd _297_/X sky130_fd_sc_hd__and2_2
XFILLER_48_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2012 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2719 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput464 _469_/X vssd vssd vccd vccd la_data_in_core[100] sky130_fd_sc_hd__buf_8
Xoutput475 _479_/X vssd vssd vccd vccd la_data_in_core[110] sky130_fd_sc_hd__buf_8
XFILLER_9_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2590 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput486 _489_/X vssd vssd vccd vccd la_data_in_core[120] sky130_fd_sc_hd__buf_8
Xoutput497 _384_/X vssd vssd vccd vccd la_data_in_core[15] sky130_fd_sc_hd__buf_8
XFILLER_5_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_406 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_220_ _220_/A _220_/B vssd vssd vccd vccd _220_/X sky130_fd_sc_hd__and2_2
XFILLER_10_4125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_151_ _151_/A vssd vssd vccd vccd _151_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_3424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_082_ _082_/A vssd vssd vccd vccd _082_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_418_ _546_/A _418_/B _418_/C vssd vssd vccd vccd _418_/X sky130_fd_sc_hd__and3b_4
XTAP_1693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_349_ _349_/A _349_/B vssd vssd vccd vccd _349_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[94\] la_data_out_core[94] _257_/X vssd vssd vccd vccd _077_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_6_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3475 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_203_ _203_/A _203_/B vssd vssd vccd vccd _203_/X sky130_fd_sc_hd__and2_4
XFILLER_49_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_134_ _134_/A vssd vssd vccd vccd _134_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_065_ _065_/A vssd vssd vccd vccd _065_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_49_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4474 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2602 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2613 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2624 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1901 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1912 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1923 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1934 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1945 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1956 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1967 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1978 _360_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1989 _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[22\] mprj_dat_i_user[22] _294_/X vssd vssd vccd vccd _136_/A sky130_fd_sc_hd__nand2_2
XFILLER_50_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[120\] la_data_out_core[120] _283_/X vssd vssd vccd vccd _103_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_6_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_809 _608_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_751 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1208 _244_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1219 _254_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_117_ _117_/A vssd vssd vccd vccd _117_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_048_ _048_/A vssd vssd vccd vccd _048_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1671 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2410 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2421 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2432 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2443 _363_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2454 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1720 _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2465 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1731 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2476 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1742 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2487 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1753 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2498 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1764 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1775 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1786 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1797 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[57\] la_data_out_core[57] _220_/X vssd vssd vccd vccd _040_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_606 _511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_617 _516_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_628 _535_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_639 _565_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2962 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1005 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1016 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1027 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1038 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1049 _167_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput320 la_oenb_mprj[39] vssd vssd vccd vccd _536_/A sky130_fd_sc_hd__clkbuf_4
Xinput331 la_oenb_mprj[49] vssd vssd vccd vccd _546_/A sky130_fd_sc_hd__buf_4
XFILLER_40_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput342 la_oenb_mprj[59] vssd vssd vccd vccd _556_/A sky130_fd_sc_hd__buf_4
XFILLER_7_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput353 la_oenb_mprj[69] vssd vssd vccd vccd _566_/A sky130_fd_sc_hd__buf_8
XFILLER_48_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput364 la_oenb_mprj[79] vssd vssd vccd vccd _576_/A sky130_fd_sc_hd__buf_8
Xinput375 la_oenb_mprj[89] vssd vssd vccd vccd _586_/A sky130_fd_sc_hd__buf_4
XFILLER_29_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput386 la_oenb_mprj[99] vssd vssd vccd vccd _596_/A sky130_fd_sc_hd__buf_6
Xinput397 mprj_adr_o_core[18] vssd vssd vccd vccd _323_/B sky130_fd_sc_hd__buf_8
XFILLER_48_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_597_ _597_/A _597_/B vssd vssd vccd vccd _597_/X sky130_fd_sc_hd__and2_4
XFILLER_43_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2 _084_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput805 _559_/X vssd vssd vccd vccd la_oenb_core[62] sky130_fd_sc_hd__buf_8
XFILLER_47_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput816 _569_/X vssd vssd vccd vccd la_oenb_core[72] sky130_fd_sc_hd__buf_8
XFILLER_42_4522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput827 _579_/X vssd vssd vccd vccd la_oenb_core[82] sky130_fd_sc_hd__buf_8
Xoutput838 _589_/X vssd vssd vccd vccd la_oenb_core[92] sky130_fd_sc_hd__buf_8
Xoutput849 _315_/X vssd vssd vccd vccd mprj_adr_o_user[10] sky130_fd_sc_hd__buf_8
XFILLER_6_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2240 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2251 _525_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2262 _358_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2273 _299_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2284 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2295 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1550 _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1561 _391_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1572 _296_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1583 _296_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1594 _213_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3923 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_520_ _520_/A _520_/B vssd vssd vccd vccd _520_/X sky130_fd_sc_hd__and2_4
XTAP_2702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_403 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_414 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1466 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_425 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_436 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_447 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_451_ _579_/A _451_/B _451_/C vssd vssd vccd vccd _451_/X sky130_fd_sc_hd__and3b_4
XTAP_2757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_458 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4270 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_469 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_382_ _510_/A _382_/B _382_/C vssd vssd vccd vccd _382_/X sky130_fd_sc_hd__and3b_4
XFILLER_15_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1018 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput150 la_iena_mprj[116] vssd vssd vccd vccd _279_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_49_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput161 la_iena_mprj[126] vssd vssd vccd vccd _289_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_48_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput172 la_iena_mprj[20] vssd vssd vccd vccd _183_/B sky130_fd_sc_hd__buf_4
XFILLER_4_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1158 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput183 la_iena_mprj[30] vssd vssd vccd vccd _193_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_37_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput194 la_iena_mprj[40] vssd vssd vccd vccd _203_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3344 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_970 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_981 _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_992 _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput602 _157_/Y vssd vssd vccd vccd la_data_in_mprj[10] sky130_fd_sc_hd__buf_8
Xoutput613 _158_/Y vssd vssd vccd vccd la_data_in_mprj[11] sky130_fd_sc_hd__buf_8
Xoutput624 _161_/Y vssd vssd vccd vccd la_data_in_mprj[14] sky130_fd_sc_hd__buf_8
XFILLER_25_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput635 _007_/Y vssd vssd vccd vccd la_data_in_mprj[24] sky130_fd_sc_hd__buf_8
Xoutput646 _017_/Y vssd vssd vccd vccd la_data_in_mprj[34] sky130_fd_sc_hd__buf_8
XFILLER_5_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput657 _027_/Y vssd vssd vccd vccd la_data_in_mprj[44] sky130_fd_sc_hd__buf_8
XFILLER_47_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput668 _037_/Y vssd vssd vccd vccd la_data_in_mprj[54] sky130_fd_sc_hd__buf_8
Xoutput679 _047_/Y vssd vssd vccd vccd la_data_in_mprj[64] sky130_fd_sc_hd__buf_8
XFILLER_29_2794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2070 la_data_out_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2081 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2092 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1380 _353_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1391 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2282 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_200 _398_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_211 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_503_ _503_/A _503_/B vssd vssd vccd vccd _503_/X sky130_fd_sc_hd__and2_4
XANTENNA_222 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_233 _434_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_244 _440_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 _441_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_266 _447_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_434_ _562_/A _434_/B _434_/C vssd vssd vccd vccd _434_/X sky130_fd_sc_hd__and3b_4
XTAP_1842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_277 _448_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_288 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_299 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_365_ _365_/A _365_/B vssd vssd vccd vccd _365_/X sky130_fd_sc_hd__and2_4
XFILLER_9_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_296_ _296_/A _296_/B vssd vssd vccd vccd _296_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2923 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_602 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[1\] la_data_out_core[1] _164_/X vssd vssd vccd vccd _148_/A
+ sky130_fd_sc_hd__nand2_1
Xoutput465 _470_/X vssd vssd vccd vccd la_data_in_core[101] sky130_fd_sc_hd__buf_8
XFILLER_5_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput476 _480_/X vssd vssd vccd vccd la_data_in_core[111] sky130_fd_sc_hd__buf_8
XFILLER_44_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput487 _490_/X vssd vssd vccd vccd la_data_in_core[121] sky130_fd_sc_hd__buf_8
XFILLER_9_2663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput498 _385_/X vssd vssd vccd vccd la_data_in_core[16] sky130_fd_sc_hd__buf_8
XFILLER_25_2444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_418 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_150_ _150_/A vssd vssd vccd vccd _150_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_14_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_081_ _081_/A vssd vssd vccd vccd _081_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_417_ _545_/A _417_/B _417_/C vssd vssd vccd vccd _417_/X sky130_fd_sc_hd__and3b_4
XTAP_1672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_348_ _348_/A _348_/B vssd vssd vccd vccd _348_/X sky130_fd_sc_hd__and2_4
XFILLER_13_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_279_ _279_/A _279_/B vssd vssd vccd vccd _279_/X sky130_fd_sc_hd__and2_4
XFILLER_48_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[87\] la_data_out_core[87] _250_/X vssd vssd vccd vccd _070_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_9_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_202_ _202_/A _202_/B vssd vssd vccd vccd _202_/X sky130_fd_sc_hd__and2_4
XFILLER_51_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_454 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_988 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_133_ _133_/A vssd vssd vccd vccd _133_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_3244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_064_ _064_/A vssd vssd vccd vccd _064_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2603 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2614 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2625 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1902 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1913 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1924 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1935 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1946 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1957 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1968 _347_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1979 _361_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[15\] mprj_dat_i_user[15] _294_/X vssd vssd vccd vccd _129_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1606 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3251 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[113\] la_data_out_core[113] _276_/X vssd vssd vccd vccd _096_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_6_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_763 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1209 _245_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4422 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3718 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_116_ _116_/A vssd vssd vccd vccd _116_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_047_ _047_/A vssd vssd vccd vccd _047_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_2400 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2411 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2422 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2433 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2444 _296_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2455 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1710 _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1721 _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2466 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1732 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2477 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1743 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2488 _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1754 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2499 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1765 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_1776 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1787 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1798 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_800 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_607 _511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_618 _516_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_629 _541_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1006 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1017 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1028 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1039 _165_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput310 la_oenb_mprj[2] vssd vssd vccd vccd _499_/A sky130_fd_sc_hd__buf_4
XFILLER_7_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput321 la_oenb_mprj[3] vssd vssd vccd vccd _500_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_3799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput332 la_oenb_mprj[4] vssd vssd vccd vccd _501_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput343 la_oenb_mprj[5] vssd vssd vccd vccd _502_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput354 la_oenb_mprj[6] vssd vssd vccd vccd _503_/A sky130_fd_sc_hd__clkbuf_4
Xinput365 la_oenb_mprj[7] vssd vssd vccd vccd _504_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput376 la_oenb_mprj[8] vssd vssd vccd vccd _505_/A sky130_fd_sc_hd__buf_4
XFILLER_40_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput387 la_oenb_mprj[9] vssd vssd vccd vccd _506_/A sky130_fd_sc_hd__clkbuf_4
Xinput398 mprj_adr_o_core[19] vssd vssd vccd vccd _324_/B sky130_fd_sc_hd__buf_8
XFILLER_21_1042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_596_ _596_/A _596_/B vssd vssd vccd vccd _596_/X sky130_fd_sc_hd__and2_4
XFILLER_16_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_3 _071_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput806 _560_/X vssd vssd vccd vccd la_oenb_core[63] sky130_fd_sc_hd__buf_8
XFILLER_42_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput817 _570_/X vssd vssd vccd vccd la_oenb_core[73] sky130_fd_sc_hd__buf_8
XFILLER_6_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput828 _580_/X vssd vssd vccd vccd la_oenb_core[83] sky130_fd_sc_hd__buf_8
Xoutput839 _590_/X vssd vssd vccd vccd la_oenb_core[93] sky130_fd_sc_hd__buf_8
XFILLER_3_4005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2807 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2230 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2241 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4038 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2252 _527_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2263 _359_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2274 la_data_out_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2285 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1540 _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2296 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1551 _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1562 _392_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_1573 _296_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1584 _477_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1595 _597_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1558 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1802 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_404 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_415 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_426 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_450_ _578_/A _450_/B _450_/C vssd vssd vccd vccd _450_/X sky130_fd_sc_hd__and3b_4
XTAP_2747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_437 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_448 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_460 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_459 _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_381_ _509_/A _381_/B _381_/C vssd vssd vccd vccd _381_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4168 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput140 la_iena_mprj[107] vssd vssd vccd vccd _270_/B sky130_fd_sc_hd__clkbuf_4
Xinput151 la_iena_mprj[117] vssd vssd vccd vccd _280_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_49_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput162 la_iena_mprj[127] vssd vssd vccd vccd _290_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput173 la_iena_mprj[21] vssd vssd vccd vccd _184_/B sky130_fd_sc_hd__buf_4
XFILLER_18_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput184 la_iena_mprj[31] vssd vssd vccd vccd _194_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput195 la_iena_mprj[41] vssd vssd vccd vccd _204_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_960 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_971 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_982 _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_579_ _579_/A _579_/B vssd vssd vccd vccd _579_/X sky130_fd_sc_hd__and2_4
XFILLER_38_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_993 _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput603 _093_/Y vssd vssd vccd vccd la_data_in_mprj[110] sky130_fd_sc_hd__buf_8
Xoutput614 _103_/Y vssd vssd vccd vccd la_data_in_mprj[120] sky130_fd_sc_hd__buf_8
XFILLER_25_4039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput625 _162_/Y vssd vssd vccd vccd la_data_in_mprj[15] sky130_fd_sc_hd__buf_8
XFILLER_47_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput636 _008_/Y vssd vssd vccd vccd la_data_in_mprj[25] sky130_fd_sc_hd__buf_8
XFILLER_29_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput647 _018_/Y vssd vssd vccd vccd la_data_in_mprj[35] sky130_fd_sc_hd__buf_8
XFILLER_42_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput658 _028_/Y vssd vssd vccd vccd la_data_in_mprj[45] sky130_fd_sc_hd__buf_8
XFILLER_25_2604 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput669 _038_/Y vssd vssd vccd vccd la_data_in_mprj[55] sky130_fd_sc_hd__buf_8
XFILLER_28_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2060 output952/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2071 la_data_out_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2082 _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2093 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1370 _342_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1381 _354_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1392 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1560 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1242 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_201 _412_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_502_ _502_/A _502_/B vssd vssd vccd vccd _502_/X sky130_fd_sc_hd__and2_4
XANTENNA_212 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_223 _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_234 _434_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_245 _440_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 _441_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_433_ _561_/A _433_/B _433_/C vssd vssd vccd vccd _433_/X sky130_fd_sc_hd__and3b_4
XTAP_1843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_267 _447_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_278 _449_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_289 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_364_ _364_/A _364_/B vssd vssd vccd vccd _364_/X sky130_fd_sc_hd__and2_4
XFILLER_35_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_295_ input3/X _295_/B vssd vssd vccd vccd _295_/X sky130_fd_sc_hd__and2b_4
XFILLER_9_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[32\] la_data_out_core[32] _195_/X vssd vssd vccd vccd _015_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_790 _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput466 _471_/X vssd vssd vccd vccd la_data_in_core[102] sky130_fd_sc_hd__buf_8
Xoutput477 _481_/X vssd vssd vccd vccd la_data_in_core[112] sky130_fd_sc_hd__buf_8
XFILLER_47_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput488 _491_/X vssd vssd vccd vccd la_data_in_core[122] sky130_fd_sc_hd__buf_8
Xoutput499 _386_/X vssd vssd vccd vccd la_data_in_core[17] sky130_fd_sc_hd__buf_8
XFILLER_9_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_080_ _080_/A vssd vssd vccd vccd _080_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_290 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_416_ _544_/A _416_/B _416_/C vssd vssd vccd vccd _416_/X sky130_fd_sc_hd__and3b_4
XTAP_1673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_347_ _347_/A _347_/B vssd vssd vccd vccd _347_/X sky130_fd_sc_hd__and2_4
XFILLER_13_3094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_278_ _278_/A _278_/B vssd vssd vccd vccd _278_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_201_ _201_/A _201_/B vssd vssd vccd vccd _201_/X sky130_fd_sc_hd__and2_2
XFILLER_11_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_132_ _132_/A vssd vssd vccd vccd _132_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_063_ _063_/A vssd vssd vccd vccd _063_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1832 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2604 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2615 _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2626 _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1903 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_1914 _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1925 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1936 _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1947 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1958 _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1969 _348_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4510 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[106\] la_data_out_core[106] _269_/X vssd vssd vccd vccd _089_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_0_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_296 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3410 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_115_ _115_/A vssd vssd vccd vccd _115_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_046_ _046_/A vssd vssd vccd vccd _046_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2401 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2412 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2423 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2434 _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_2445 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1700 _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1711 _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2456 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1722 _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2467 _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1733 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2478 _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1744 _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2489 _592_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1755 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1766 _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1777 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1788 _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1799 _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2306 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_608 _511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_619 _517_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3730 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2683 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3964 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1007 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_1018 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_1029 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput300 la_oenb_mprj[20] vssd vssd vccd vccd _517_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput311 la_oenb_mprj[30] vssd vssd vccd vccd _527_/A sky130_fd_sc_hd__buf_6
Xinput322 la_oenb_mprj[40] vssd vssd vccd vccd _537_/A sky130_fd_sc_hd__buf_8
XFILLER_40_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput333 la_oenb_mprj[50] vssd vssd vccd vccd _547_/A sky130_fd_sc_hd__clkbuf_8
Xinput344 la_oenb_mprj[60] vssd vssd vccd vccd _557_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput355 la_oenb_mprj[70] vssd vssd vccd vccd _567_/A sky130_fd_sc_hd__buf_8
Xinput366 la_oenb_mprj[80] vssd vssd vccd vccd _577_/A sky130_fd_sc_hd__buf_8
Xinput377 la_oenb_mprj[90] vssd vssd vccd vccd _587_/A sky130_fd_sc_hd__buf_4
XFILLER_48_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput388 mprj_adr_o_core[0] vssd vssd vccd vccd _305_/B sky130_fd_sc_hd__buf_8
XFILLER_40_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput399 mprj_adr_o_core[1] vssd vssd vccd vccd _306_/B sky130_fd_sc_hd__buf_8
XFILLER_29_650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1190 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3516 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_595_ _595_/A _595_/B vssd vssd vccd vccd _595_/X sky130_fd_sc_hd__and2_2
XFILLER_31_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_4 _072_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput807 _561_/X vssd vssd vccd vccd la_oenb_core[64] sky130_fd_sc_hd__buf_8
Xoutput818 _571_/X vssd vssd vccd vccd la_oenb_core[74] sky130_fd_sc_hd__buf_8
XFILLER_49_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput829 _581_/X vssd vssd vccd vccd la_oenb_core[84] sky130_fd_sc_hd__buf_8
XFILLER_6_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_029_ _029_/A vssd vssd vccd vccd _029_/Y sky130_fd_sc_hd__inv_2
XANTENNA_2220 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_2231 _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2819 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2242 _382_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2253 _547_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2264 _361_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1530 _384_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2275 la_data_out_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2286 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1541 _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2297 mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1552 _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1563 _392_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1574 _296_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_1585 _491_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[62\] la_data_out_core[62] _225_/X vssd vssd vccd vccd _045_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_39_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1596 _598_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_405 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_416 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_427 _479_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_438 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_449 _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_380_ _508_/A _380_/B _380_/C vssd vssd vccd vccd _380_/X sky130_fd_sc_hd__and3b_4
XFILLER_25_185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput130 la_data_out_mprj[99] vssd vssd vccd vccd _468_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput141 la_iena_mprj[108] vssd vssd vccd vccd _271_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput152 la_iena_mprj[118] vssd vssd vccd vccd _281_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput163 la_iena_mprj[12] vssd vssd vccd vccd _175_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput174 la_iena_mprj[22] vssd vssd vccd vccd _185_/B sky130_fd_sc_hd__buf_4
Xinput185 la_iena_mprj[32] vssd vssd vccd vccd _195_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput196 la_iena_mprj[42] vssd vssd vccd vccd _205_/B sky130_fd_sc_hd__buf_4
XTAP_4673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_4036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_950 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_961 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_578_ _578_/A _578_/B vssd vssd vccd vccd _578_/X sky130_fd_sc_hd__and2_4
XANTENNA_972 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_983 _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_994 _327_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput604 _094_/Y vssd vssd vccd vccd la_data_in_mprj[111] sky130_fd_sc_hd__buf_8
XFILLER_29_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput615 _104_/Y vssd vssd vccd vccd la_data_in_mprj[121] sky130_fd_sc_hd__buf_8
XFILLER_44_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput626 _163_/Y vssd vssd vccd vccd la_data_in_mprj[16] sky130_fd_sc_hd__buf_8
XFILLER_47_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput637 _009_/Y vssd vssd vccd vccd la_data_in_mprj[26] sky130_fd_sc_hd__buf_8
Xoutput648 _019_/Y vssd vssd vccd vccd la_data_in_mprj[36] sky130_fd_sc_hd__buf_8
XFILLER_25_3328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput659 _029_/Y vssd vssd vccd vccd la_data_in_mprj[46] sky130_fd_sc_hd__buf_8
XFILLER_42_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2616 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2050 _351_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2061 output953/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2072 mprj_dat_i_user[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_2083 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_2094 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
.ends

