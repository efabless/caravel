* NGSPICE file created from mgmt_protect.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufbuf_8 abstract view
.subckt sky130_fd_sc_hd__bufbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for mprj2_logic_high abstract view
.subckt mprj2_logic_high HI vccd2 vssd2
.ends

* Black-box entry subcircuit for mprj_logic_high abstract view
.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[287] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295]
+ HI[296] HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304]
+ HI[305] HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314]
+ HI[315] HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334]
+ HI[335] HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344]
+ HI[345] HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354]
+ HI[355] HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374]
+ HI[375] HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384]
+ HI[385] HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394]
+ HI[395] HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403]
+ HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413]
+ HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423]
+ HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[42] HI[430] HI[431] HI[432] HI[433]
+ HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443]
+ HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453]
+ HI[454] HI[455] HI[456] HI[457] HI[458] HI[459] HI[45] HI[460] HI[461] HI[462] HI[46]
+ HI[47] HI[48] HI[49] HI[4] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57]
+ HI[58] HI[59] HI[5] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68]
+ HI[69] HI[6] HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79]
+ HI[7] HI[80] HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8]
+ HI[90] HI[91] HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1
+ vssd1
.ends

* Black-box entry subcircuit for mgmt_protect_hv abstract view
.subckt mgmt_protect_hv vccd vssd vdda1 vssa1 vdda2 vssa2 mprj2_vdd_logic1 mprj_vdd_logic1
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102]
+ la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107]
+ la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[10] la_iena_mprj[110] la_iena_mprj[111]
+ la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116]
+ la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[11] la_iena_mprj[120]
+ la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125]
+ la_iena_mprj[126] la_iena_mprj[127] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14]
+ la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19]
+ la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23]
+ la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28]
+ la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32]
+ la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37]
+ la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3] la_iena_mprj[40] la_iena_mprj[41]
+ la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46]
+ la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[4] la_iena_mprj[50]
+ la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55]
+ la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[5]
+ la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64]
+ la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69]
+ la_iena_mprj[6] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73]
+ la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78]
+ la_iena_mprj[79] la_iena_mprj[7] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82]
+ la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87]
+ la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[8] la_iena_mprj[90] la_iena_mprj[91]
+ la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96]
+ la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[9] la_oenb_core[0]
+ la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104]
+ la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109]
+ la_oenb_core[10] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113]
+ la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118]
+ la_oenb_core[119] la_oenb_core[11] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122]
+ la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127]
+ la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16]
+ la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[1] la_oenb_core[20]
+ la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25]
+ la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[2]
+ la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34]
+ la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39]
+ la_oenb_core[3] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43]
+ la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48]
+ la_oenb_core[49] la_oenb_core[4] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52]
+ la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57]
+ la_oenb_core[58] la_oenb_core[59] la_oenb_core[5] la_oenb_core[60] la_oenb_core[61]
+ la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66]
+ la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[6] la_oenb_core[70]
+ la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75]
+ la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[7]
+ la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84]
+ la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89]
+ la_oenb_core[8] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93]
+ la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98]
+ la_oenb_core[99] la_oenb_core[9] la_oenb_mprj[0] la_oenb_mprj[100] la_oenb_mprj[101]
+ la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106]
+ la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[10] la_oenb_mprj[110]
+ la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115]
+ la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[11]
+ la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124]
+ la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] la_oenb_mprj[12] la_oenb_mprj[13]
+ la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18]
+ la_oenb_mprj[19] la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22]
+ la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27]
+ la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31]
+ la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36]
+ la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40]
+ la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45]
+ la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4]
+ la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54]
+ la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59]
+ la_oenb_mprj[5] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63]
+ la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68]
+ la_oenb_mprj[69] la_oenb_mprj[6] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72]
+ la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77]
+ la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[7] la_oenb_mprj[80] la_oenb_mprj[81]
+ la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86]
+ la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[8] la_oenb_mprj[90]
+ la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95]
+ la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[9]
+ mprj_ack_i_core mprj_ack_i_user mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11]
+ mprj_adr_o_core[12] mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15]
+ mprj_adr_o_core[16] mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19]
+ mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23]
+ mprj_adr_o_core[24] mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27]
+ mprj_adr_o_core[28] mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31]
+ mprj_adr_o_core[3] mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7]
+ mprj_adr_o_core[8] mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11]
+ mprj_adr_o_user[12] mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15]
+ mprj_adr_o_user[16] mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19]
+ mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23]
+ mprj_adr_o_user[24] mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27]
+ mprj_adr_o_user[28] mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31]
+ mprj_adr_o_user[3] mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7]
+ mprj_adr_o_user[8] mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0]
+ mprj_dat_i_core[10] mprj_dat_i_core[11] mprj_dat_i_core[12] mprj_dat_i_core[13]
+ mprj_dat_i_core[14] mprj_dat_i_core[15] mprj_dat_i_core[16] mprj_dat_i_core[17]
+ mprj_dat_i_core[18] mprj_dat_i_core[19] mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21]
+ mprj_dat_i_core[22] mprj_dat_i_core[23] mprj_dat_i_core[24] mprj_dat_i_core[25]
+ mprj_dat_i_core[26] mprj_dat_i_core[27] mprj_dat_i_core[28] mprj_dat_i_core[29]
+ mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31] mprj_dat_i_core[3] mprj_dat_i_core[4]
+ mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7] mprj_dat_i_core[8] mprj_dat_i_core[9]
+ mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11] mprj_dat_i_user[12] mprj_dat_i_user[13]
+ mprj_dat_i_user[14] mprj_dat_i_user[15] mprj_dat_i_user[16] mprj_dat_i_user[17]
+ mprj_dat_i_user[18] mprj_dat_i_user[19] mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21]
+ mprj_dat_i_user[22] mprj_dat_i_user[23] mprj_dat_i_user[24] mprj_dat_i_user[25]
+ mprj_dat_i_user[26] mprj_dat_i_user[27] mprj_dat_i_user[28] mprj_dat_i_user[29]
+ mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31] mprj_dat_i_user[3] mprj_dat_i_user[4]
+ mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7] mprj_dat_i_user[8] mprj_dat_i_user[9]
+ mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13]
+ mprj_dat_o_core[14] mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17]
+ mprj_dat_o_core[18] mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21]
+ mprj_dat_o_core[22] mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25]
+ mprj_dat_o_core[26] mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29]
+ mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4]
+ mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9]
+ mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13]
+ mprj_dat_o_user[14] mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17]
+ mprj_dat_o_user[18] mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21]
+ mprj_dat_o_user[22] mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25]
+ mprj_dat_o_user[26] mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29]
+ mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4]
+ mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9]
+ mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2] mprj_sel_o_core[3]
+ mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3] mprj_stb_o_core
+ mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood user1_vdd_powergood
+ user2_vcc_powergood user2_vdd_powergood user_clock user_clock2 user_irq[0] user_irq[1]
+ user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2] user_irq_ena[0] user_irq_ena[1]
+ user_irq_ena[2] user_reset vccd vccd1_uq1 vccd2_uq0 vdda1_uq0 vdda2_uq0 vssd vssd1_uq1
+ vssa1_uq0 vssa2_uq0 vssd2_uq0
XTAP_188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[34\]_A la_data_out_core[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__203__B _203_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_406 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input127_A la_data_out_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_501_ _501_/A _501_/B vssd vssd vccd vccd _501_/X sky130_fd_sc_hd__and2_4
XTAP_2512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_432_ _560_/A _432_/B _432_/C vssd vssd vccd vccd _432_/X sky130_fd_sc_hd__and3b_4
XTAP_2567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_363_ _363_/A _363_/B vssd vssd vccd vccd _363_/X sky130_fd_sc_hd__and2_4
XTAP_1888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input92_A la_data_out_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_294_ _294_/A _294_/B vssd vssd vccd vccd _294_/X sky130_fd_sc_hd__and2_4
XFILLER_13_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xrebuffer7 wire1248/X vssd vssd vccd vccd rebuffer7/X sky130_fd_sc_hd__bufbuf_8
Xuser_wb_dat_gates\[8\] mprj_dat_i_user[8] wire1245/X vssd vssd vccd vccd wire993/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_6_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[25\]_A la_data_out_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output513_A _371_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1144_A wire1145/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output882_A wire976/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[25\] la_data_out_core[25] _188_/X vssd vssd vccd vccd _008_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_36_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1680_A wire1681/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[16\]_A la_data_out_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[100\]_A la_data_out_core[100] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__304__A _304_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput467 wire1057/X vssd vssd vccd vccd la_data_in_core[103] sky130_fd_sc_hd__buf_8
Xoutput478 _482_/X vssd vssd vccd vccd la_data_in_core[113] sky130_fd_sc_hd__buf_8
Xoutput489 _492_/X vssd vssd vccd vccd la_data_in_core[123] sky130_fd_sc_hd__buf_8
XFILLER_5_2507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1209 _317_/X vssd vssd vccd vccd wire1209/X sky130_fd_sc_hd__buf_6
XFILLER_25_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__490__A_N _618_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__214__A _214_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input244_A la_iena_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1710 wire1710/A vssd vssd vccd vccd _459_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1721 wire1721/A vssd vssd vccd vccd _448_/B sky130_fd_sc_hd__buf_6
Xwire1732 wire1732/A vssd vssd vccd vccd wire1732/X sky130_fd_sc_hd__buf_6
XFILLER_1_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input411_A mprj_adr_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_415_ _543_/A _415_/B _415_/C vssd vssd vccd vccd _415_/X sky130_fd_sc_hd__and3b_4
XTAP_1652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_346_ _346_/A _346_/B vssd vssd vccd vccd _346_/X sky130_fd_sc_hd__and2_4
XFILLER_35_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_277_ _277_/A _277_/B vssd vssd vccd vccd _277_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output463_A _369_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__124__A _124_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output728_A wire1043/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1359_A wire1359/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1526_A wire1526/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire979_A _121_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__034__A _034_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2390 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_max_cap1246_A split13/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1006 wire1006/A vssd vssd vccd vccd wire1006/X sky130_fd_sc_hd__buf_6
Xwire1017 wire1018/X vssd vssd vccd vccd _134_/A sky130_fd_sc_hd__buf_6
XFILLER_5_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1028 wire1028/A vssd vssd vccd vccd _125_/A sky130_fd_sc_hd__buf_8
XFILLER_38_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1039 _615_/X vssd vssd vccd vccd wire1039/X sky130_fd_sc_hd__buf_6
XFILLER_0_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__209__A _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_762 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_200_ _200_/A _200_/B vssd vssd vccd vccd _200_/X sky130_fd_sc_hd__and2_2
XFILLER_23_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_131_ _131_/A vssd vssd vccd vccd _131_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_32_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input194_A la_iena_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_062_ _062_/A vssd vssd vccd vccd _062_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_3_600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__386__A_N _514_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input361_A la_oenb_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input459_A mprj_we_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input55_A la_data_out_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__598__B _598_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1540 wire1540/A vssd vssd vccd vccd _174_/A sky130_fd_sc_hd__buf_6
Xwire1551 wire1551/A vssd vssd vccd vccd _625_/A sky130_fd_sc_hd__buf_6
XFILLER_1_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1562 wire1563/X vssd vssd vccd vccd _619_/B sky130_fd_sc_hd__buf_6
Xwire1573 wire1573/A vssd vssd vccd vccd wire1573/X sky130_fd_sc_hd__buf_6
XFILLER_19_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1584 wire1585/X vssd vssd vccd vccd _607_/B sky130_fd_sc_hd__buf_6
Xwire1595 wire1595/A vssd vssd vccd vccd _598_/B sky130_fd_sc_hd__buf_6
XFILLER_0_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__119__A _119_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output580_A wire1066/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output678_A _046_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_329_ _329_/A _329_/B vssd vssd vccd vccd _329_/X sky130_fd_sc_hd__and2_1
XFILLER_32_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output845_A _596_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1476_A wire1476/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2839 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[92\] la_data_out_core[92] _255_/X vssd vssd vccd vccd _075_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_45_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3314 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3358 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__301__B _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__029__A _029_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3695 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input207_A la_iena_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_114_ _114_/A vssd vssd vccd vccd _114_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_32_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_045_ _045_/A vssd vssd vccd vccd _045_/Y sky130_fd_sc_hd__inv_2
XTAP_507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1057_A _472_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__401__A_N _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1370 wire1371/X vssd vssd vccd vccd _334_/B sky130_fd_sc_hd__buf_6
Xwire1381 wire1381/A vssd vssd vccd vccd wire1381/X sky130_fd_sc_hd__buf_6
XFILLER_39_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1392 wire1393/X vssd vssd vccd vccd wire1392/X sky130_fd_sc_hd__buf_6
XFILLER_21_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1224_A _307_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output795_A _550_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[20\] mprj_dat_i_user[20] split13/A vssd vssd vccd vccd wire1018/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA_wire1593_A wire1593/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__312__A _312_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2684 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__222__A _222_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input157_A la_iena_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput301 la_oenb_mprj[21] vssd vssd vccd vccd _518_/A sky130_fd_sc_hd__buf_4
XANTENNA__424__A_N _552_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput312 la_oenb_mprj[31] vssd vssd vccd vccd _528_/A sky130_fd_sc_hd__buf_4
XFILLER_0_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput323 la_oenb_mprj[41] vssd vssd vccd vccd _538_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput334 la_oenb_mprj[51] vssd vssd vccd vccd _548_/A sky130_fd_sc_hd__buf_6
Xinput345 la_oenb_mprj[61] vssd vssd vccd vccd _558_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput356 la_oenb_mprj[71] vssd vssd vccd vccd _568_/A sky130_fd_sc_hd__buf_4
Xinput367 la_oenb_mprj[81] vssd vssd vccd vccd _578_/A sky130_fd_sc_hd__buf_4
XFILLER_22_3492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input324_A la_oenb_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput378 la_oenb_mprj[91] vssd vssd vccd vccd _588_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput389 mprj_adr_o_core[10] vssd vssd vccd vccd wire1417/A sky130_fd_sc_hd__buf_6
XFILLER_40_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input18_A la_data_out_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_594_ _594_/A _594_/B vssd vssd vccd vccd _594_/X sky130_fd_sc_hd__and2_4
XFILLER_16_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_2404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_5 _439_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput808 _562_/X vssd vssd vccd vccd la_oenb_core[65] sky130_fd_sc_hd__buf_8
Xoutput819 _572_/X vssd vssd vccd vccd la_oenb_core[75] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[70\]_B _233_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_028_ _028_/A vssd vssd vccd vccd _028_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_3971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output543_A wire1078/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__132__A _132_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1174_A wire1175/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output710_A _075_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output808_A _562_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1341_A wire1341/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1439_A wire1439/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[55\] la_data_out_core[55] _218_/X vssd vssd vccd vccd _038_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_26_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1606_A wire1606/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__307__A _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire961_A _146_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[61\]_B _224_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__447__A_N _575_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__042__A _042_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__217__A _217_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input274_A la_oenb_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[52\]_B _215_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_rebuffer10_A wire1245/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input441_A mprj_dat_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput120 la_data_out_mprj[8] vssd vssd vccd vccd _377_/C sky130_fd_sc_hd__clkbuf_4
Xinput131 la_data_out_mprj[9] vssd vssd vccd vccd _378_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput142 la_iena_mprj[109] vssd vssd vccd vccd _272_/B sky130_fd_sc_hd__clkbuf_4
Xinput153 la_iena_mprj[119] vssd vssd vccd vccd _282_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput164 la_iena_mprj[13] vssd vssd vccd vccd _176_/B sky130_fd_sc_hd__clkbuf_4
Xinput175 la_iena_mprj[23] vssd vssd vccd vccd _186_/B sky130_fd_sc_hd__clkbuf_4
Xinput186 la_iena_mprj[33] vssd vssd vccd vccd _196_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput197 la_iena_mprj[43] vssd vssd vccd vccd _206_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_577_ _577_/A _577_/B vssd vssd vccd vccd _577_/X sky130_fd_sc_hd__and2_4
XFILLER_18_2635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output493_A wire1054/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__127__A _127_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output660_A _030_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output758_A _498_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1291_A wire1291/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1389_A wire1390/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput605 _095_/Y vssd vssd vccd vccd la_data_in_mprj[112] sky130_fd_sc_hd__buf_8
XFILLER_9_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput616 _105_/Y vssd vssd vccd vccd la_data_in_mprj[122] sky130_fd_sc_hd__buf_8
XFILLER_9_3537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput627 _000_/Y vssd vssd vccd vccd la_data_in_mprj[17] sky130_fd_sc_hd__buf_8
Xoutput638 _010_/Y vssd vssd vccd vccd la_data_in_mprj[27] sky130_fd_sc_hd__buf_8
XFILLER_29_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output925_A wire1134/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput649 _020_/Y vssd vssd vccd vccd la_data_in_mprj[37] sky130_fd_sc_hd__buf_8
XFILLER_28_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1556_A wire1557/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3086 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1723_A wire1723/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__037__A _037_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__500__A _500_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_500_ _500_/A _500_/B vssd vssd vccd vccd _500_/X sky130_fd_sc_hd__and2_4
XFILLER_19_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_431_ _559_/A _431_/B _431_/C vssd vssd vccd vccd _431_/X sky130_fd_sc_hd__and3b_2
XFILLER_26_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_362_ _362_/A _362_/B vssd vssd vccd vccd _362_/X sky130_fd_sc_hd__and2_4
XTAP_1867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_293_ _293_/A _293_/B vssd vssd vccd vccd _293_/X sky130_fd_sc_hd__and2_4
XFILLER_35_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input391_A mprj_adr_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input85_A la_data_out_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xrebuffer8 wire1248/X vssd vssd vccd vccd rebuffer8/X sky130_fd_sc_hd__bufbuf_8
XFILLER_13_2598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[25\]_B _188_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2672 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output506_A _392_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1137_A _356_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1304_A wire1305/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output875_A wire1221/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[18\] la_data_out_core[18] _181_/X vssd vssd vccd vccd _001_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_31_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[100\]_B wire1257/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__304__B _304_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput468 _473_/X vssd vssd vccd vccd la_data_in_core[104] sky130_fd_sc_hd__buf_8
Xoutput479 _483_/X vssd vssd vccd vccd la_data_in_core[114] sky130_fd_sc_hd__buf_8
XFILLER_5_2519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__320__A _320_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_rebuffer8_A wire1248/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__214__B _214_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__230__A _230_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1700 wire1700/A vssd vssd vccd vccd _469_/B sky130_fd_sc_hd__buf_6
XFILLER_1_3618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1711 wire1711/A vssd vssd vccd vccd _458_/B sky130_fd_sc_hd__buf_6
XFILLER_28_1392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1722 wire1722/A vssd vssd vccd vccd _447_/B sky130_fd_sc_hd__buf_6
XANTENNA_input237_A la_iena_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input404_A mprj_adr_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_414_ _542_/A _414_/B _414_/C vssd vssd vccd vccd _414_/X sky130_fd_sc_hd__and3b_4
XTAP_1642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_345_ _345_/A _345_/B vssd vssd vccd vccd _345_/X sky130_fd_sc_hd__and2_4
XFILLER_41_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_276_ _276_/A _276_/B vssd vssd vccd vccd _276_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1087_A _417_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__140__A _140_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_402 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__315__A _315_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__050__A _050_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1007 wire1008/X vssd vssd vccd vccd _140_/A sky130_fd_sc_hd__buf_6
XFILLER_2_3938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1018 wire1018/A vssd vssd vccd vccd wire1018/X sky130_fd_sc_hd__buf_6
XFILLER_2_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1029 wire1029/A vssd vssd vccd vccd _124_/A sky130_fd_sc_hd__buf_8
XFILLER_38_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__209__B _209_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_130_ _130_/A vssd vssd vccd vccd _130_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_7_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_061_ _061_/A vssd vssd vccd vccd _061_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_input187_A la_iena_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input354_A la_oenb_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input48_A la_data_out_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1530 wire1530/A vssd vssd vccd vccd _184_/A sky130_fd_sc_hd__buf_6
Xwire1541 wire1541/A vssd vssd vccd vccd _173_/A sky130_fd_sc_hd__buf_6
Xwire1552 wire1553/X vssd vssd vccd vccd _624_/B sky130_fd_sc_hd__buf_6
XFILLER_46_321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1563 wire1563/A vssd vssd vccd vccd wire1563/X sky130_fd_sc_hd__buf_6
XFILLER_4_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1574 wire1575/X vssd vssd vccd vccd _613_/B sky130_fd_sc_hd__buf_6
Xwire1585 wire1585/A vssd vssd vccd vccd wire1585/X sky130_fd_sc_hd__buf_6
XFILLER_19_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1596 wire1596/A vssd vssd vccd vccd _597_/B sky130_fd_sc_hd__buf_6
XFILLER_46_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_328_ _328_/A _328_/B vssd vssd vccd vccd _328_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1002_A wire1002/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output573_A _453_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__135__A _135_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_259_ _259_/A _259_/B vssd vssd vccd vccd _259_/X sky130_fd_sc_hd__and2_1
XFILLER_31_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output740_A wire1038/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output838_A _589_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1371_A wire1371/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3326 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__480__A_N _608_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2542 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[85\] la_data_out_core[85] _248_/X vssd vssd vccd vccd _068_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_44_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1636_A wire1636/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__045__A _045_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input102_A la_data_out_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_113_ _113_/A vssd vssd vccd vccd _113_/Y sky130_fd_sc_hd__clkinv_2
X_044_ _044_/A vssd vssd vccd vccd _044_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__402__B _402_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1126 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1360 wire1361/X vssd vssd vccd vccd _308_/B sky130_fd_sc_hd__buf_6
Xwire1371 wire1371/A vssd vssd vccd vccd wire1371/X sky130_fd_sc_hd__buf_6
XFILLER_21_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_3289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1382 wire1383/X vssd vssd vccd vccd _328_/B sky130_fd_sc_hd__buf_6
Xwire1393 wire1393/A vssd vssd vccd vccd wire1393/X sky130_fd_sc_hd__buf_6
XFILLER_19_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output690_A _057_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1217_A _313_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output788_A _544_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output955_A wire1242/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[13\] mprj_dat_i_user[13] rebuffer11/X vssd vssd vccd vccd wire1026/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA_wire1586_A wire1586/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__312__B _312_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[1\]_A mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[111\] la_data_out_core[111] _274_/X vssd vssd vccd vccd _094_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_2909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__376__A_N _504_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[1\]_A la_data_out_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__503__A _503_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput302 la_oenb_mprj[22] vssd vssd vccd vccd _519_/A sky130_fd_sc_hd__buf_4
Xinput313 la_oenb_mprj[32] vssd vssd vccd vccd _529_/A sky130_fd_sc_hd__buf_4
XFILLER_27_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput324 la_oenb_mprj[42] vssd vssd vccd vccd _539_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput335 la_oenb_mprj[52] vssd vssd vccd vccd _549_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput346 la_oenb_mprj[62] vssd vssd vccd vccd _559_/A sky130_fd_sc_hd__clkbuf_4
Xinput357 la_oenb_mprj[72] vssd vssd vccd vccd _569_/A sky130_fd_sc_hd__buf_4
Xinput368 la_oenb_mprj[82] vssd vssd vccd vccd _579_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput379 la_oenb_mprj[92] vssd vssd vccd vccd _589_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input317_A la_oenb_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_593_ _593_/A _593_/B vssd vssd vccd vccd _593_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_6 wire1706/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput809 _563_/X vssd vssd vccd vccd la_oenb_core[66] sky130_fd_sc_hd__buf_8
X_027_ _027_/A vssd vssd vccd vccd _027_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output536_A wire1085/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1167_A _341_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output703_A _069_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__399__A_N _527_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1334_A wire1335/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1190 wire1191/X vssd vssd vccd vccd wire1190/X sky130_fd_sc_hd__buf_6
XFILLER_39_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[48\] la_data_out_core[48] _211_/X vssd vssd vccd vccd _031_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_34_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1501_A wire1501/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__307__B _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__323__A _323_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3852 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__217__B _217_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__233__A _233_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input267_A la_oenb_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input434_A mprj_dat_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput110 la_data_out_mprj[80] vssd vssd vccd vccd _449_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput121 la_data_out_mprj[90] vssd vssd vccd vccd _459_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_input30_A la_data_out_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput132 la_iena_mprj[0] vssd vssd vccd vccd _625_/B sky130_fd_sc_hd__clkbuf_4
Xinput143 la_iena_mprj[10] vssd vssd vccd vccd _173_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput154 la_iena_mprj[11] vssd vssd vccd vccd _174_/B sky130_fd_sc_hd__buf_4
XFILLER_2_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput165 la_iena_mprj[14] vssd vssd vccd vccd _177_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput176 la_iena_mprj[24] vssd vssd vccd vccd _187_/B sky130_fd_sc_hd__clkbuf_4
Xinput187 la_iena_mprj[34] vssd vssd vccd vccd _197_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput198 la_iena_mprj[44] vssd vssd vccd vccd _207_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_36_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_576_ _576_/A _576_/B vssd vssd vccd vccd _576_/X sky130_fd_sc_hd__and2_4
XFILLER_16_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output486_A _489_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput606 _096_/Y vssd vssd vccd vccd la_data_in_mprj[113] sky130_fd_sc_hd__buf_8
XANTENNA__143__A _143_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput617 _106_/Y vssd vssd vccd vccd la_data_in_mprj[123] sky130_fd_sc_hd__buf_8
Xoutput628 _001_/Y vssd vssd vccd vccd la_data_in_mprj[18] sky130_fd_sc_hd__buf_8
XANTENNA_wire1284_A wire1285/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput639 _011_/Y vssd vssd vccd vccd la_data_in_mprj[28] sky130_fd_sc_hd__buf_8
XFILLER_45_2011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output820_A _573_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output918_A wire1146/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1451_A wire1451/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1549_A wire1549/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1716_A wire1716/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__318__A _318_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__414__A_N _542_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__053__A _053_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__500__B _500_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_430_ _558_/A _430_/B _430_/C vssd vssd vccd vccd _430_/X sky130_fd_sc_hd__and3b_2
XFILLER_19_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__228__A _228_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_361_ _361_/A _361_/B vssd vssd vccd vccd _361_/X sky130_fd_sc_hd__and2_4
XTAP_1868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_292_ _292_/A _292_/B vssd vssd vccd vccd _292_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input384_A la_oenb_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xrebuffer9 wire1245/A vssd vssd vccd vccd rebuffer9/X sky130_fd_sc_hd__bufbuf_8
XANTENNA_input78_A la_data_out_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__410__B _410_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__437__A_N _565_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__138__A _138_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_559_ _559_/A _559_/B vssd vssd vccd vccd _559_/X sky130_fd_sc_hd__and2_4
XFILLER_31_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output770_A _527_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output868_A wire1182/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1499_A wire1499/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1666_A wire1667/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput469 wire1056/X vssd vssd vccd vccd la_data_in_core[105] sky130_fd_sc_hd__buf_8
XANTENNA__601__A _601_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__320__B _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__048__A _048_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_628 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__511__A _511_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__230__B _230_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1701 wire1701/A vssd vssd vccd vccd _468_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1712 wire1712/A vssd vssd vccd vccd _457_/B sky130_fd_sc_hd__buf_6
Xwire1723 wire1723/A vssd vssd vccd vccd _446_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input132_A la_iena_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_413_ _541_/A _413_/B _413_/C vssd vssd vccd vccd _413_/X sky130_fd_sc_hd__and3b_4
XTAP_2377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_344_ _344_/A _344_/B vssd vssd vccd vccd _344_/X sky130_fd_sc_hd__and2_4
XTAP_1698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_275_ _275_/A _275_/B vssd vssd vccd vccd _275_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__405__B _405_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output616_A _105_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1414_A wire1414/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[30\] la_data_out_core[30] _193_/X vssd vssd vccd vccd _013_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_17_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__315__B _315_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1150 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__331__A _331_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2835 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1008 wire1008/A vssd vssd vccd vccd wire1008/X sky130_fd_sc_hd__buf_6
Xwire1019 wire1019/A vssd vssd vccd vccd _115_/A sky130_fd_sc_hd__buf_8
XFILLER_25_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_ack_gate_A mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__506__A _506_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_060_ _060_/A vssd vssd vccd vccd _060_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_20_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__241__A _241_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input347_A la_oenb_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1520 wire1520/A vssd vssd vccd vccd _234_/A sky130_fd_sc_hd__buf_6
Xwire1531 wire1531/A vssd vssd vccd vccd _183_/A sky130_fd_sc_hd__buf_6
XFILLER_21_3377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1542 wire1542/A vssd vssd vccd vccd _172_/A sky130_fd_sc_hd__buf_6
XFILLER_21_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1553 wire1553/A vssd vssd vccd vccd wire1553/X sky130_fd_sc_hd__buf_6
Xwire1564 wire1565/X vssd vssd vccd vccd _618_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1076 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1575 wire1575/A vssd vssd vccd vccd wire1575/X sky130_fd_sc_hd__buf_6
Xwire1586 wire1586/A vssd vssd vccd vccd _606_/B sky130_fd_sc_hd__buf_6
Xwire1597 wire1597/A vssd vssd vccd vccd _596_/B sky130_fd_sc_hd__buf_6
XFILLER_46_377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_327_ _327_/A _327_/B vssd vssd vccd vccd _327_/X sky130_fd_sc_hd__and2_4
X_258_ _258_/A _258_/B vssd vssd vccd vccd _258_/X sky130_fd_sc_hd__and2_1
XFILLER_10_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output566_A _447_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_189_ _189_/A _189_/B vssd vssd vccd vccd _189_/X sky130_fd_sc_hd__and2_2
XFILLER_45_3823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1197_A wire1198/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output733_A _609_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1364_A wire1364/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output900_A _141_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[78\] la_data_out_core[78] _241_/X vssd vssd vccd vccd _061_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_6_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_3972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire984_A _116_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__326__A _326_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1879 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[91\]_A la_data_out_core[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__061__A _061_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__236__A _236_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input297_A la_oenb_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_112_ _112_/A vssd vssd vccd vccd _112_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[82\]_A la_data_out_core[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_043_ _043_/A vssd vssd vccd vccd _043_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input60_A la_data_out_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1350 wire1351/X vssd vssd vccd vccd wire1350/X sky130_fd_sc_hd__buf_6
XFILLER_5_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1361 wire1362/X vssd vssd vccd vccd wire1361/X sky130_fd_sc_hd__buf_6
XFILLER_19_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_3279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1372 wire1373/X vssd vssd vccd vccd _333_/B sky130_fd_sc_hd__buf_6
Xwire1383 wire1383/A vssd vssd vccd vccd wire1383/X sky130_fd_sc_hd__buf_6
XFILLER_46_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1394 wire1395/X vssd vssd vccd vccd _324_/B sky130_fd_sc_hd__buf_6
XFILLER_1_1866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1112_A wire1113/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output683_A _051_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__146__A _146_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output850_A wire1210/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[73\]_A la_data_out_core[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output948_A wire1227/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1481_A wire1481/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1579_A wire1579/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[104\] la_data_out_core[104] wire1253/X vssd vssd vccd vccd
+ _087_/A sky130_fd_sc_hd__nand2_4
XFILLER_26_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[1\]_B _164_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__056__A _056_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[64\]_A la_data_out_core[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__503__B _503_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput303 la_oenb_mprj[23] vssd vssd vccd vccd _520_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_1_969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput314 la_oenb_mprj[33] vssd vssd vccd vccd _530_/A sky130_fd_sc_hd__clkbuf_4
Xinput325 la_oenb_mprj[43] vssd vssd vccd vccd _540_/A sky130_fd_sc_hd__buf_4
Xinput336 la_oenb_mprj[53] vssd vssd vccd vccd _550_/A sky130_fd_sc_hd__clkbuf_4
Xinput347 la_oenb_mprj[63] vssd vssd vccd vccd _560_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_40_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput358 la_oenb_mprj[73] vssd vssd vccd vccd _570_/A sky130_fd_sc_hd__buf_4
XFILLER_2_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput369 la_oenb_mprj[83] vssd vssd vccd vccd _580_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input212_A la_iena_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_592_ _592_/A _592_/B vssd vssd vccd vccd _592_/X sky130_fd_sc_hd__and2_2
XFILLER_38_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3254 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__470__A_N _598_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[55\]_A la_data_out_core[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_7 wire1706/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_026_ _026_/A vssd vssd vccd vccd _026_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_4123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__413__B _413_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output529_A wire1091/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1180 wire1181/X vssd vssd vccd vccd wire1180/X sky130_fd_sc_hd__buf_6
XFILLER_1_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1191 _329_/X vssd vssd vccd vccd wire1191/X sky130_fd_sc_hd__buf_6
XANTENNA_wire1327_A wire1327/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output898_A _139_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1696_A wire1696/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[46\]_A la_data_out_core[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__604__A _604_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__323__B _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__493__A_N _621_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[37\]_A la_data_out_core[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[121\]_A la_data_out_core[121] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__514__A _514_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__233__B _233_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input162_A la_iena_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput100 la_data_out_mprj[71] vssd vssd vccd vccd _440_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput111 la_data_out_mprj[81] vssd vssd vccd vccd _450_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput122 la_data_out_mprj[91] vssd vssd vccd vccd _460_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput133 la_iena_mprj[100] vssd vssd vccd vccd _263_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input427_A mprj_dat_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput144 la_iena_mprj[110] vssd vssd vccd vccd _273_/B sky130_fd_sc_hd__clkbuf_4
Xinput155 la_iena_mprj[120] vssd vssd vccd vccd _283_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput166 la_iena_mprj[15] vssd vssd vccd vccd _178_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_input23_A la_data_out_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput177 la_iena_mprj[25] vssd vssd vccd vccd _188_/B sky130_fd_sc_hd__clkbuf_4
Xinput188 la_iena_mprj[35] vssd vssd vccd vccd _198_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput199 la_iena_mprj[45] vssd vssd vccd vccd _208_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_575_ _575_/A _575_/B vssd vssd vccd vccd _575_/X sky130_fd_sc_hd__and2_4
XFILLER_44_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__408__B _408_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[28\]_A la_data_out_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output479_A _483_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[112\]_A la_data_out_core[112] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_8_376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput607 _097_/Y vssd vssd vccd vccd la_data_in_mprj[114] sky130_fd_sc_hd__buf_8
XFILLER_9_3528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput618 _107_/Y vssd vssd vccd vccd la_data_in_mprj[124] sky130_fd_sc_hd__buf_8
XFILLER_29_3467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput629 _002_/Y vssd vssd vccd vccd la_data_in_mprj[19] sky130_fd_sc_hd__buf_8
XANTENNA_output646_A _017_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_009_ _009_/A vssd vssd vccd vccd _009_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1277_A wire1277/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output813_A _503_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1444_A wire1445/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[60\] la_data_out_core[60] _223_/X vssd vssd vccd vccd _043_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_3_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1758 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1611_A wire1611/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1709_A wire1709/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__318__B _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[19\]_A la_data_out_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__334__A _334_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_A la_data_out_core[103] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_30_2358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__509__A _509_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__228__B _228_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_360_ _360_/A _360_/B vssd vssd vccd vccd _360_/X sky130_fd_sc_hd__and2_4
XFILLER_17_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_291_ _291_/A _291_/B vssd vssd vccd vccd _291_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__244__A _244_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__389__A_N _517_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input377_A la_oenb_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_558_ _558_/A _558_/B vssd vssd vccd vccd _558_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1025_A wire1025/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output596_A _087_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_489_ _617_/A _489_/B _489_/C vssd vssd vccd vccd _489_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output763_A _521_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__154__A _154_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1394_A wire1395/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output930_A wire1124/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1561_A wire1561/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1659_A wire1659/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__601__B _601_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__329__A _329_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__064__A _064_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput960 wire1243/X vssd vssd vccd vccd user_reset sky130_fd_sc_hd__buf_8
XANTENNA__511__B _511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1702 wire1702/A vssd vssd vccd vccd _467_/B sky130_fd_sc_hd__buf_6
Xwire1713 wire1713/A vssd vssd vccd vccd _456_/B sky130_fd_sc_hd__buf_6
Xwire1724 wire1724/A vssd vssd vccd vccd _445_/B sky130_fd_sc_hd__buf_6
XFILLER_19_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input125_A la_data_out_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__239__A _239_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_412_ _540_/A _412_/B _412_/C vssd vssd vccd vccd _412_/X sky130_fd_sc_hd__and3b_4
XTAP_2367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_968 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_343_ _343_/A _343_/B vssd vssd vccd vccd _343_/X sky130_fd_sc_hd__and2_4
XTAP_1688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input90_A la_data_out_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_274_ _274_/A _274_/B vssd vssd vccd vccd _274_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__405__C _405_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[6\] mprj_dat_i_user[6] rebuffer2/X vssd vssd vccd vccd wire995/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_6_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__404__A_N _532_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output511_A wire1107/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output609_A _099_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1142_A wire1143/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1407_A wire1408/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output880_A wire1239/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[23\] la_data_out_core[23] _186_/X vssd vssd vccd vccd _006_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_36_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3122 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__612__A _612_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2803 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__331__B _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2847 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1009 wire1009/A vssd vssd vccd vccd _139_/A sky130_fd_sc_hd__buf_6
XFILLER_3_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__059__A _059_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__506__B _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3238 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__522__A _522_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__241__B _241_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__427__A_N _555_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput790 _546_/X vssd vssd vccd vccd la_oenb_core[49] sky130_fd_sc_hd__buf_8
XANTENNA_input242_A la_iena_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1510 wire1510/A vssd vssd vccd vccd _260_/A sky130_fd_sc_hd__buf_6
Xwire1521 wire1521/A vssd vssd vccd vccd _193_/A sky130_fd_sc_hd__buf_4
XFILLER_5_2863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1532 wire1532/A vssd vssd vccd vccd _182_/A sky130_fd_sc_hd__buf_6
XFILLER_5_2874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1543 wire1543/A vssd vssd vccd vccd _171_/A sky130_fd_sc_hd__buf_6
XFILLER_1_2727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1554 wire1555/X vssd vssd vccd vccd _623_/B sky130_fd_sc_hd__buf_6
Xwire1565 wire1565/A vssd vssd vccd vccd wire1565/X sky130_fd_sc_hd__buf_6
XFILLER_4_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1576 wire1577/X vssd vssd vccd vccd _612_/B sky130_fd_sc_hd__buf_6
XFILLER_0_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1587 wire1588/X vssd vssd vccd vccd _605_/B sky130_fd_sc_hd__buf_6
Xwire1598 wire1598/A vssd vssd vccd vccd _595_/B sky130_fd_sc_hd__buf_6
XTAP_2120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1438 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_326_ _326_/A _326_/B vssd vssd vccd vccd _326_/X sky130_fd_sc_hd__and2_4
XFILLER_9_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__416__B _416_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_257_ _257_/A _257_/B vssd vssd vccd vccd _257_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_188_ _188_/A _188_/B vssd vssd vccd vccd _188_/X sky130_fd_sc_hd__and2_2
XANTENNA_output559_A wire1068/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1092_A _412_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2522 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output726_A _603_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1357_A wire1358/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1524_A wire1524/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__607__A _607_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__326__B _326_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire977_A _123_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[91\]_B _254_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__517__A _517_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__236__B _236_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_111_ _111_/A vssd vssd vccd vccd _111_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input192_A la_iena_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[82\]_B _245_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_042_ _042_/A vssd vssd vccd vccd _042_/Y sky130_fd_sc_hd__inv_2
XANTENNA__252__A _252_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input457_A mprj_sel_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input53_A la_data_out_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1340 wire1341/X vssd vssd vccd vccd _337_/B sky130_fd_sc_hd__buf_6
Xwire1351 wire1351/A vssd vssd vccd vccd wire1351/X sky130_fd_sc_hd__buf_6
XFILLER_1_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1362 wire1362/A vssd vssd vccd vccd wire1362/X sky130_fd_sc_hd__buf_6
XFILLER_1_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1373 wire1373/A vssd vssd vccd vccd wire1373/X sky130_fd_sc_hd__buf_6
Xwire1384 wire1385/X vssd vssd vccd vccd _327_/B sky130_fd_sc_hd__buf_6
Xwire1395 wire1395/A vssd vssd vccd vccd wire1395/X sky130_fd_sc_hd__buf_6
XFILLER_21_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1878 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_309_ _309_/A _309_/B vssd vssd vccd vccd _309_/X sky130_fd_sc_hd__and2_4
XFILLER_30_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[73\]_B _236_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output843_A _594_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1474_A wire1475/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[90\] la_data_out_core[90] _253_/X vssd vssd vccd vccd _073_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_6_3125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3158 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1641_A wire1641/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__337__A _337_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[64\]_B _227_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__072__A _072_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput304 la_oenb_mprj[24] vssd vssd vccd vccd _521_/A sky130_fd_sc_hd__buf_4
XFILLER_2_3512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput315 la_oenb_mprj[34] vssd vssd vccd vccd _531_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput326 la_oenb_mprj[44] vssd vssd vccd vccd _541_/A sky130_fd_sc_hd__clkbuf_4
Xinput337 la_oenb_mprj[54] vssd vssd vccd vccd _551_/A sky130_fd_sc_hd__buf_4
XFILLER_29_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput348 la_oenb_mprj[64] vssd vssd vccd vccd _561_/A sky130_fd_sc_hd__buf_4
Xinput359 la_oenb_mprj[74] vssd vssd vccd vccd _571_/A sky130_fd_sc_hd__buf_4
XFILLER_40_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_591_ _591_/A _591_/B vssd vssd vccd vccd _591_/X sky130_fd_sc_hd__and2_4
XFILLER_29_687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input205_A la_iena_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__247__A _247_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[55\]_B _218_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_025_ _025_/A vssd vssd vccd vccd _025_/Y sky130_fd_sc_hd__inv_2
XANTENNA_8 _314_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2650 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1170 wire1171/X vssd vssd vccd vccd wire1170/X sky130_fd_sc_hd__buf_6
XFILLER_19_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1181 _334_/X vssd vssd vccd vccd wire1181/X sky130_fd_sc_hd__buf_6
XFILLER_39_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1192 wire1193/X vssd vssd vccd vccd wire1192/X sky130_fd_sc_hd__buf_6
XFILLER_1_1631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__295__A_N _295_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1222_A _309_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output793_A _548_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output960_A wire1243/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1591_A wire1591/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1689_A wire1690/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__604__B _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__620__A _620_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1946 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__067__A _067_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[121\]_B _284_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__514__B _514_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__530__A _530_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input155_A la_iena_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput101 la_data_out_mprj[72] vssd vssd vccd vccd _441_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput112 la_data_out_mprj[82] vssd vssd vccd vccd _451_/C sky130_fd_sc_hd__clkbuf_4
Xinput123 la_data_out_mprj[92] vssd vssd vccd vccd _461_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput134 la_iena_mprj[101] vssd vssd vccd vccd _264_/B sky130_fd_sc_hd__clkbuf_4
Xinput145 la_iena_mprj[111] vssd vssd vccd vccd _274_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput156 la_iena_mprj[121] vssd vssd vccd vccd _284_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input322_A la_oenb_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput167 la_iena_mprj[16] vssd vssd vccd vccd _179_/B sky130_fd_sc_hd__clkbuf_4
Xinput178 la_iena_mprj[26] vssd vssd vccd vccd _189_/B sky130_fd_sc_hd__clkbuf_4
Xinput189 la_iena_mprj[36] vssd vssd vccd vccd _199_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input16_A la_data_out_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_574_ _574_/A _574_/B vssd vssd vccd vccd _574_/X sky130_fd_sc_hd__and2_4
XANTENNA_user_wb_dat_gates\[30\]_A mprj_dat_i_user[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[112\]_B _275_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput608 _098_/Y vssd vssd vccd vccd la_data_in_mprj[115] sky130_fd_sc_hd__buf_8
Xoutput619 _108_/Y vssd vssd vccd vccd la_data_in_mprj[125] sky130_fd_sc_hd__buf_8
X_008_ _008_/A vssd vssd vccd vccd _008_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output541_A wire1080/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output639_A _011_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1172_A wire1173/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output806_A _560_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1437_A wire1437/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_4129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[53\] la_data_out_core[53] _216_/X vssd vssd vccd vccd _036_/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA_wire1604_A wire1604/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[21\]_A mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__615__A _615_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[19\]_B _182_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__334__B _334_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_B wire1254/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__460__A_N _588_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input8_A la_data_out_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3684 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__509__B _509_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[12\]_A mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_290_ _290_/A _290_/B vssd vssd vccd vccd _290_/X sky130_fd_sc_hd__and2_4
XFILLER_13_3225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__525__A _525_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__244__B _244_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input272_A la_oenb_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__260__A _260_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__419__B _419_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_557_ _557_/A _557_/B vssd vssd vccd vccd _557_/X sky130_fd_sc_hd__and2_2
XFILLER_44_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_488_ _616_/A _488_/B _488_/C vssd vssd vccd vccd _488_/X sky130_fd_sc_hd__and3b_4
XANTENNA_output491_A _494_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output589_A _468_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output756_A _515_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1387_A wire1388/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__483__A_N _611_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output923_A wire1136/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__170__A _170_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1554_A wire1555/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1721_A wire1721/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__329__B _329_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__080__A _080_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput950 wire1235/X vssd vssd vccd vccd mprj_we_o_user sky130_fd_sc_hd__buf_8
XFILLER_25_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1703 wire1703/A vssd vssd vccd vccd _466_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1714 wire1714/A vssd vssd vccd vccd _455_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1725 wire1725/A vssd vssd vccd vccd _444_/B sky130_fd_sc_hd__buf_6
XFILLER_4_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__239__B _239_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input118_A la_data_out_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_411_ _539_/A _411_/B _411_/C vssd vssd vccd vccd _411_/X sky130_fd_sc_hd__and3b_4
XFILLER_14_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_342_ _342_/A _342_/B vssd vssd vccd vccd _342_/X sky130_fd_sc_hd__and2_4
XTAP_1678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__255__A _255_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_273_ _273_/A _273_/B vssd vssd vccd vccd _273_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input83_A la_data_out_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output504_A _390_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1135_A _357_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_609_ _609_/A _609_/B vssd vssd vccd vccd _609_/X sky130_fd_sc_hd__and2_4
XFILLER_33_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1302_A wire1303/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output873_A wire1223/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__165__A _165_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[16\] la_data_out_core[16] _179_/X vssd vssd vccd vccd _163_/A
+ sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_gates\[29\] mprj_dat_i_user[29] wire1248/X vssd vssd vccd vccd wire1002/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_31_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1671_A wire1671/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__612__B _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2859 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[127\] la_data_out_core[127] _290_/X vssd vssd vccd vccd _110_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_3_1331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__379__A_N _507_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__075__A _075_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_rebuffer6_A wire1248/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__522__B _522_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput780 _500_/X vssd vssd vccd vccd la_oenb_core[3] sky130_fd_sc_hd__buf_8
XFILLER_21_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput791 _501_/X vssd vssd vccd vccd la_oenb_core[4] sky130_fd_sc_hd__buf_8
XFILLER_40_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1500 wire1500/A vssd vssd vccd vccd _270_/A sky130_fd_sc_hd__buf_6
XFILLER_21_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1511 wire1511/A vssd vssd vccd vccd _259_/A sky130_fd_sc_hd__buf_6
XFILLER_21_3357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input235_A la_iena_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1522 wire1522/A vssd vssd vccd vccd _192_/A sky130_fd_sc_hd__buf_6
XFILLER_4_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1533 wire1533/A vssd vssd vccd vccd _181_/A sky130_fd_sc_hd__buf_6
XFILLER_19_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1544 wire1544/A vssd vssd vccd vccd _170_/A sky130_fd_sc_hd__buf_6
XFILLER_8_1286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1555 wire1555/A vssd vssd vccd vccd wire1555/X sky130_fd_sc_hd__buf_6
XFILLER_46_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1566 wire1567/X vssd vssd vccd vccd _617_/B sky130_fd_sc_hd__buf_6
Xwire1577 wire1577/A vssd vssd vccd vccd wire1577/X sky130_fd_sc_hd__buf_6
XFILLER_21_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1588 wire1588/A vssd vssd vccd vccd wire1588/X sky130_fd_sc_hd__buf_6
XFILLER_21_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1599 wire1600/X vssd vssd vccd vccd _297_/A sky130_fd_sc_hd__buf_6
XFILLER_19_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input402_A mprj_adr_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_325_ _325_/A _325_/B vssd vssd vccd vccd _325_/X sky130_fd_sc_hd__and2_4
XFILLER_30_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_256_ _256_/A _256_/B vssd vssd vccd vccd _256_/X sky130_fd_sc_hd__and2_1
XFILLER_7_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_187_ _187_/A _187_/B vssd vssd vccd vccd _187_/X sky130_fd_sc_hd__and2_1
XFILLER_45_3803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__432__B _432_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1085_A _419_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output621_A _110_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output719_A _497_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__607__B _607_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__623__A _623_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__342__B _342_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[4\]_A mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[4\]_A la_data_out_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__517__B _517_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_574 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_110_ _110_/A vssd vssd vccd vccd _110_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__533__A _533_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_041_ _041_/A vssd vssd vccd vccd _041_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input185_A la_iena_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__252__B _252_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input352_A la_oenb_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_4063 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input46_A la_data_out_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1330 wire1331/X vssd vssd vccd vccd _351_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1341 wire1341/A vssd vssd vccd vccd wire1341/X sky130_fd_sc_hd__buf_6
Xwire1352 wire1353/X vssd vssd vccd vccd _311_/B sky130_fd_sc_hd__buf_6
XFILLER_46_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1363 wire1364/X vssd vssd vccd vccd _336_/B sky130_fd_sc_hd__buf_6
Xwire1374 wire1375/X vssd vssd vccd vccd _332_/B sky130_fd_sc_hd__buf_6
Xwire1385 wire1385/A vssd vssd vccd vccd wire1385/X sky130_fd_sc_hd__buf_6
XFILLER_1_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1396 wire1397/X vssd vssd vccd vccd _323_/B sky130_fd_sc_hd__buf_6
XFILLER_21_1752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_308_ _308_/A _308_/B vssd vssd vccd vccd _308_/X sky130_fd_sc_hd__and2_4
XFILLER_15_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1000_A wire1000/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output571_A _451_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output669_A _038_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_239_ _239_/A _239_/B vssd vssd vccd vccd _239_/X sky130_fd_sc_hd__and2_4
XFILLER_13_1291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output836_A _587_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1467_A wire1468/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[83\] la_data_out_core[83] _246_/X vssd vssd vccd vccd _066_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_44_1218 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1634_A wire1634/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__618__A _618_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__337__B _337_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__417__A_N _545_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_894 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput305 la_oenb_mprj[25] vssd vssd vccd vccd _522_/A sky130_fd_sc_hd__buf_4
Xinput316 la_oenb_mprj[35] vssd vssd vccd vccd _532_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput327 la_oenb_mprj[45] vssd vssd vccd vccd _542_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput338 la_oenb_mprj[55] vssd vssd vccd vccd _552_/A sky130_fd_sc_hd__buf_4
XFILLER_5_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput349 la_oenb_mprj[65] vssd vssd vccd vccd _562_/A sky130_fd_sc_hd__buf_4
XFILLER_6_2970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_590_ _590_/A _590_/B vssd vssd vccd vccd _590_/X sky130_fd_sc_hd__and2_4
XFILLER_2_2889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_699 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__528__A _528_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__247__B _247_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input100_A la_data_out_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__263__A _263_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_9 _314_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_024_ _024_/A vssd vssd vccd vccd _024_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_2504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1160 wire1161/X vssd vssd vccd vccd wire1160/X sky130_fd_sc_hd__buf_6
Xwire1171 _339_/X vssd vssd vccd vccd wire1171/X sky130_fd_sc_hd__buf_6
XFILLER_1_3089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1182 wire1183/X vssd vssd vccd vccd wire1182/X sky130_fd_sc_hd__buf_6
XFILLER_19_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1193 _328_/X vssd vssd vccd vccd wire1193/X sky130_fd_sc_hd__buf_6
XFILLER_36_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1215_A wire1216/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output786_A wire1052/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output953_A wire1729/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__173__A _173_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[11\] mprj_dat_i_user[11] wire1245/X vssd vssd vccd vccd wire1028/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_30_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1584_A wire1585/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__620__B _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2110 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_374 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__083__A _083_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__530__B _530_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput102 la_data_out_mprj[73] vssd vssd vccd vccd _442_/C sky130_fd_sc_hd__clkbuf_4
Xinput113 la_data_out_mprj[83] vssd vssd vccd vccd _452_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput124 la_data_out_mprj[93] vssd vssd vccd vccd _462_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input148_A la_iena_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput135 la_iena_mprj[102] vssd vssd vccd vccd _265_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput146 la_iena_mprj[112] vssd vssd vccd vccd _275_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput157 la_iena_mprj[122] vssd vssd vccd vccd _285_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput168 la_iena_mprj[17] vssd vssd vccd vccd _180_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput179 la_iena_mprj[27] vssd vssd vccd vccd _190_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_29_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input315_A la_oenb_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__258__A _258_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_573_ _573_/A _573_/B vssd vssd vccd vccd _573_/X sky130_fd_sc_hd__and2_4
XFILLER_18_2606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[30\]_B wire1248/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3086 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput609 _099_/Y vssd vssd vccd vccd la_data_in_mprj[116] sky130_fd_sc_hd__buf_8
XFILLER_29_2724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_007_ _007_/A vssd vssd vccd vccd _007_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__440__B _440_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output534_A wire1086/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1165_A _342_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output701_A _067_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1332_A wire1333/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__168__A _168_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[46\] la_data_out_core[46] _209_/X vssd vssd vccd vccd _029_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[21\]_B split13/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__615__B _615_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[8\] la_data_out_core[8] _171_/X vssd vssd vccd vccd _155_/A
+ sky130_fd_sc_hd__nand2_2
XANTENNA__350__B _350_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__078__A _078_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[12\]_B wire1245/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__525__B _525_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1250 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__541__A _541_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input265_A la_oenb_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input432_A mprj_dat_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_625_ _625_/A _625_/B vssd vssd vccd vccd _625_/X sky130_fd_sc_hd__and2_2
XFILLER_29_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__419__C _419_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_556_ _556_/A _556_/B vssd vssd vccd vccd _556_/X sky130_fd_sc_hd__and2_4
XFILLER_17_488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_487_ _615_/A _487_/B _487_/C vssd vssd vccd vccd _487_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__435__B _435_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output484_A _488_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output749_A wire1032/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1282_A wire1283/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__170__B _170_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output916_A wire1150/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1547_A wire1547/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1430 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1714_A wire1714/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__345__B _345_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__361__A _361_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput940 wire1164/X vssd vssd vccd vccd mprj_dat_o_user[5] sky130_fd_sc_hd__buf_8
XFILLER_28_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput951 wire1467/X vssd vssd vccd vccd user1_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_5_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1330 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1704 wire1704/A vssd vssd vccd vccd _465_/B sky130_fd_sc_hd__buf_6
XFILLER_25_2963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1715 wire1715/A vssd vssd vccd vccd _454_/B sky130_fd_sc_hd__buf_6
XFILLER_41_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1726 wire1726/A vssd vssd vccd vccd _443_/B sky130_fd_sc_hd__buf_6
XTAP_491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_410_ _538_/A _410_/B _410_/C vssd vssd vccd vccd _410_/X sky130_fd_sc_hd__and3b_2
XTAP_1602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__536__A _536_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_341_ _341_/A _341_/B vssd vssd vccd vccd _341_/X sky130_fd_sc_hd__and2_4
XFILLER_36_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_272_ _272_/A _272_/B vssd vssd vccd vccd _272_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input382_A la_oenb_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input76_A la_data_out_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__271__A _271_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_608_ _608_/A _608_/B vssd vssd vccd vccd _608_/X sky130_fd_sc_hd__and2_4
XTAP_3593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1030_A wire1030/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1128_A wire1129/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output699_A _065_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_539_ _539_/A _539_/B vssd vssd vccd vccd _539_/X sky130_fd_sc_hd__and2_4
XFILLER_15_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__165__B _165_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__450__A_N _578_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output866_A wire1186/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1497_A wire1497/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__181__A _181_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1664_A wire1665/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3572 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__356__A _356_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[94\]_A la_data_out_core[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput770 _527_/X vssd vssd vccd vccd la_oenb_core[30] sky130_fd_sc_hd__buf_8
XFILLER_5_3522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput781 _537_/X vssd vssd vccd vccd la_oenb_core[40] sky130_fd_sc_hd__buf_8
XFILLER_25_3461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput792 wire1051/X vssd vssd vccd vccd la_oenb_core[50] sky130_fd_sc_hd__buf_8
XFILLER_8_1221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1501 wire1501/A vssd vssd vccd vccd _269_/A sky130_fd_sc_hd__buf_6
XFILLER_5_3588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1512 wire1512/A vssd vssd vccd vccd _258_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1523 wire1523/A vssd vssd vccd vccd _191_/A sky130_fd_sc_hd__buf_6
XFILLER_21_3369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1534 wire1534/A vssd vssd vccd vccd _180_/A sky130_fd_sc_hd__buf_6
XFILLER_4_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1545 wire1545/A vssd vssd vccd vccd _169_/A sky130_fd_sc_hd__buf_6
XFILLER_19_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input130_A la_data_out_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1556 wire1557/X vssd vssd vccd vccd _622_/B sky130_fd_sc_hd__buf_6
Xwire1567 wire1567/A vssd vssd vccd vccd wire1567/X sky130_fd_sc_hd__buf_6
Xwire1578 wire1579/X vssd vssd vccd vccd _611_/B sky130_fd_sc_hd__buf_6
XANTENNA_input228_A la_iena_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1589 wire1589/A vssd vssd vccd vccd _604_/B sky130_fd_sc_hd__buf_6
XFILLER_21_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_2531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__473__A_N _601_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__266__A _266_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_324_ _324_/A _324_/B vssd vssd vccd vccd _324_/X sky130_fd_sc_hd__and2_2
XFILLER_32_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[85\]_A la_data_out_core[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1142 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_255_ _255_/A _255_/B vssd vssd vccd vccd _255_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_186_ _186_/A _186_/B vssd vssd vccd vccd _186_/X sky130_fd_sc_hd__and2_2
XFILLER_6_4009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__432__C _432_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1078_A _426_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output614_A _103_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1245_A wire1245/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_594 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__176__A _176_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_A la_data_out_core[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__623__B _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__496__A_N _624_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[4\]_B _167_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__086__A _086_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[67\]_A la_data_out_core[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_040_ _040_/A vssd vssd vccd vccd _040_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__533__B _533_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input178_A la_iena_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input345_A la_oenb_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4075 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input39_A la_data_out_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1320 wire1321/X vssd vssd vccd vccd _356_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1331 wire1331/A vssd vssd vccd vccd wire1331/X sky130_fd_sc_hd__buf_6
XFILLER_1_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1342 wire1343/X vssd vssd vccd vccd _298_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1353 wire1353/A vssd vssd vccd vccd wire1353/X sky130_fd_sc_hd__buf_6
Xwire1364 wire1364/A vssd vssd vccd vccd wire1364/X sky130_fd_sc_hd__buf_6
XFILLER_21_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1375 wire1375/A vssd vssd vccd vccd wire1375/X sky130_fd_sc_hd__buf_6
Xwire1386 wire1387/X vssd vssd vccd vccd _326_/B sky130_fd_sc_hd__buf_6
Xwire1397 wire1398/X vssd vssd vccd vccd wire1397/X sky130_fd_sc_hd__buf_6
XFILLER_1_2559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[58\]_A la_data_out_core[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_307_ _307_/A _307_/B vssd vssd vccd vccd _307_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_238_ _238_/A _238_/B vssd vssd vccd vccd _238_/X sky130_fd_sc_hd__and2_4
XANTENNA__443__B _443_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output564_A _445_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__369__A_N _497_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_169_ _169_/A _169_/B vssd vssd vccd vccd _169_/X sky130_fd_sc_hd__and2_2
XANTENNA_wire1195_A _327_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output731_A wire1042/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output829_A _581_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[76\] la_data_out_core[76] _239_/X vssd vssd vccd vccd _059_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_23_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__618__B _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire982_A _118_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[49\]_A la_data_out_core[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__353__B _353_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput306 la_oenb_mprj[26] vssd vssd vccd vccd _523_/A sky130_fd_sc_hd__clkbuf_4
Xinput317 la_oenb_mprj[36] vssd vssd vccd vccd _533_/A sky130_fd_sc_hd__buf_4
XFILLER_2_3525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput328 la_oenb_mprj[46] vssd vssd vccd vccd _543_/A sky130_fd_sc_hd__clkbuf_4
Xinput339 la_oenb_mprj[56] vssd vssd vccd vccd _553_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__528__B _528_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[124\]_A la_data_out_core[124] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__544__A _544_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input295_A la_oenb_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_023_ _023_/A vssd vssd vccd vccd _023_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_46_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input462_A user_irq_ena[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1150 wire1151/X vssd vssd vccd vccd wire1150/X sky130_fd_sc_hd__buf_6
Xwire1161 _344_/X vssd vssd vccd vccd wire1161/X sky130_fd_sc_hd__buf_6
XFILLER_1_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1172 wire1173/X vssd vssd vccd vccd wire1172/X sky130_fd_sc_hd__buf_6
XFILLER_40_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1183 _333_/X vssd vssd vccd vccd wire1183/X sky130_fd_sc_hd__buf_6
XFILLER_34_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1194 wire1195/X vssd vssd vccd vccd wire1194/X sky130_fd_sc_hd__buf_6
XANTENNA__438__B _438_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1208_A wire1209/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output681_A _049_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output779_A _536_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[115\]_A la_data_out_core[115] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__173__B _173_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1354 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output946_A wire1231/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1577_A wire1577/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[102\] la_data_out_core[102] wire1255/X vssd vssd vccd vccd
+ _085_/A sky130_fd_sc_hd__nand2_4
XFILLER_26_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__348__B _348_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__364__A _364_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_A la_data_out_core[106] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_11_3121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput103 la_data_out_mprj[74] vssd vssd vccd vccd _443_/C sky130_fd_sc_hd__clkbuf_4
Xinput114 la_data_out_mprj[84] vssd vssd vccd vccd _453_/C sky130_fd_sc_hd__clkbuf_4
Xinput125 la_data_out_mprj[94] vssd vssd vccd vccd _463_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput136 la_iena_mprj[103] vssd vssd vccd vccd _266_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput147 la_iena_mprj[113] vssd vssd vccd vccd _276_/B sky130_fd_sc_hd__clkbuf_4
Xinput158 la_iena_mprj[123] vssd vssd vccd vccd _286_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput169 la_iena_mprj[18] vssd vssd vccd vccd _181_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__539__A _539_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input210_A la_iena_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_572_ _572_/A _572_/B vssd vssd vccd vccd _572_/X sky130_fd_sc_hd__and2_4
XFILLER_44_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input308_A la_oenb_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__274__A _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_006_ _006_/A vssd vssd vccd vccd _006_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__440__C _440_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__407__A_N _535_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output527_A wire1093/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1158_A wire1159/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__168__B _168_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1325_A wire1325/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output896_A wire963/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[39\] la_data_out_core[39] _202_/X vssd vssd vccd vccd _022_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_36_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__184__A _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1694_A wire1695/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__359__A _359_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__541__B _541_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input160_A la_iena_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input258_A la_iena_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2070 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input425_A mprj_dat_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input21_A la_data_out_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__269__A _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_624_ _624_/A _624_/B vssd vssd vccd vccd _624_/X sky130_fd_sc_hd__and2_2
XFILLER_44_220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_555_ _555_/A _555_/B vssd vssd vccd vccd _555_/X sky130_fd_sc_hd__and2_2
XFILLER_18_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_486_ _614_/A _486_/B _486_/C vssd vssd vccd vccd _486_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__435__C _435_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output477_A _481_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_4102 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__451__B _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output644_A _015_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1275_A wire1276/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3074 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output811_A _565_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output909_A wire980/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1442_A wire1443/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__179__A _179_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1442 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1707_A wire1707/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__361__B _361_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput930 wire1124/X vssd vssd vccd vccd mprj_dat_o_user[25] sky130_fd_sc_hd__buf_8
Xoutput941 wire1162/X vssd vssd vccd vccd mprj_dat_o_user[6] sky130_fd_sc_hd__buf_8
XFILLER_9_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput952 output952/A vssd vssd vccd vccd user1_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_43_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1342 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1705 wire1705/A vssd vssd vccd vccd _464_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1716 wire1716/A vssd vssd vccd vccd _453_/B sky130_fd_sc_hd__buf_6
XTAP_470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1727 wire1727/A vssd vssd vccd vccd _442_/B sky130_fd_sc_hd__buf_6
XFILLER_3_3461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__089__A _089_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_340_ _340_/A _340_/B vssd vssd vccd vccd _340_/X sky130_fd_sc_hd__and2_4
XFILLER_39_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__536__B _536_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_271_ _271_/A _271_/B vssd vssd vccd vccd _271_/X sky130_fd_sc_hd__and2_4
XFILLER_39_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__552__A _552_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input375_A la_oenb_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input69_A la_data_out_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_607_ _607_/A _607_/B vssd vssd vccd vccd _607_/X sky130_fd_sc_hd__and2_1
XFILLER_37_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__446__B _446_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_538_ _538_/A _538_/B vssd vssd vccd vccd _538_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1023_A wire1023/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output594_A wire987/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_469_ _597_/A _469_/B _469_/C vssd vssd vccd vccd _469_/X sky130_fd_sc_hd__and3b_2
XFILLER_32_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1700 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output761_A _519_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output859_A wire1225/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1110 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1392_A wire1393/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1657_A wire1657/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__356__B _356_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[94\]_B _257_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput760 _518_/X vssd vssd vccd vccd la_oenb_core[21] sky130_fd_sc_hd__buf_8
XFILLER_21_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput771 _528_/X vssd vssd vccd vccd la_oenb_core[31] sky130_fd_sc_hd__buf_8
XFILLER_40_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput782 _538_/X vssd vssd vccd vccd la_oenb_core[41] sky130_fd_sc_hd__buf_8
XFILLER_8_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput793 _548_/X vssd vssd vccd vccd la_oenb_core[51] sky130_fd_sc_hd__buf_8
XFILLER_28_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2822 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1502 wire1502/A vssd vssd vccd vccd _268_/A sky130_fd_sc_hd__buf_6
Xwire1513 wire1513/A vssd vssd vccd vccd _257_/A sky130_fd_sc_hd__buf_4
Xwire1524 wire1524/A vssd vssd vccd vccd _190_/A sky130_fd_sc_hd__buf_6
Xwire1535 wire1535/A vssd vssd vccd vccd _179_/A sky130_fd_sc_hd__buf_6
Xwire1546 wire1546/A vssd vssd vccd vccd _168_/A sky130_fd_sc_hd__buf_6
XFILLER_21_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1557 wire1557/A vssd vssd vccd vccd wire1557/X sky130_fd_sc_hd__buf_6
Xwire1568 wire1569/X vssd vssd vccd vccd _616_/B sky130_fd_sc_hd__buf_6
XFILLER_46_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1579 wire1579/A vssd vssd vccd vccd wire1579/X sky130_fd_sc_hd__buf_6
XANTENNA_input123_A la_data_out_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__547__A _547_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_323_ _323_/A _323_/B vssd vssd vccd vccd _323_/X sky130_fd_sc_hd__and2_4
XFILLER_42_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[85\]_B _248_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_254_ _254_/A _254_/B vssd vssd vccd vccd _254_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1154 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__282__A _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_185_ _185_/A _185_/B vssd vssd vccd vccd _185_/X sky130_fd_sc_hd__and2_1
XFILLER_13_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[4\] mprj_dat_i_user[4] max_cap1244/X vssd vssd vccd vccd wire997/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_6_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output607_A _097_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1140_A wire1141/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_540 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1238_A _299_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_562 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__176__B _176_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1405_A wire1406/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[21\] la_data_out_core[21] _184_/X vssd vssd vccd vccd _004_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_37_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3664 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[76\]_B _239_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__192__A _192_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1902 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__367__A _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3406 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[67\]_B _230_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput590 _378_/X vssd vssd vccd vccd la_data_in_core[9] sky130_fd_sc_hd__buf_8
XFILLER_5_4087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input240_A la_iena_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input338_A la_oenb_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1310 wire1311/X vssd vssd vccd vccd _360_/B sky130_fd_sc_hd__buf_6
XFILLER_40_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1321 wire1321/A vssd vssd vccd vccd wire1321/X sky130_fd_sc_hd__buf_6
XANTENNA__440__A_N _568_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1332 wire1333/X vssd vssd vccd vccd _350_/B sky130_fd_sc_hd__buf_6
Xwire1343 wire1343/A vssd vssd vccd vccd wire1343/X sky130_fd_sc_hd__buf_6
Xwire1354 wire1355/X vssd vssd vccd vccd _310_/B sky130_fd_sc_hd__buf_6
Xwire1365 wire1366/X vssd vssd vccd vccd _335_/B sky130_fd_sc_hd__buf_6
XFILLER_19_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1376 wire1377/X vssd vssd vccd vccd _331_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1387 wire1388/X vssd vssd vccd vccd wire1387/X sky130_fd_sc_hd__buf_6
Xwire1398 wire1398/A vssd vssd vccd vccd wire1398/X sky130_fd_sc_hd__buf_6
XANTENNA__277__A _277_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[58\]_B _221_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_306_ _306_/A _306_/B vssd vssd vccd vccd _306_/X sky130_fd_sc_hd__and2_4
XFILLER_12_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_237_ _237_/A _237_/B vssd vssd vccd vccd _237_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__443__C _443_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_168_ _168_/A _168_/B vssd vssd vccd vccd _168_/X sky130_fd_sc_hd__and2_2
XFILLER_13_1271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output557_A wire1111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_099_ _099_/A vssd vssd vccd vccd _099_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_wire1090_A _414_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1188_A wire1189/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output724_A _601_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1355_A wire1356/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_4107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[69\] la_data_out_core[69] _232_/X vssd vssd vccd vccd _052_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_39_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__187__A _187_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire975_A _125_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__463__A_N _591_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput307 la_oenb_mprj[27] vssd vssd vccd vccd _524_/A sky130_fd_sc_hd__clkbuf_4
Xinput318 la_oenb_mprj[37] vssd vssd vccd vccd _534_/A sky130_fd_sc_hd__buf_4
Xinput329 la_oenb_mprj[47] vssd vssd vccd vccd _544_/A sky130_fd_sc_hd__buf_4
XFILLER_44_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__097__A _097_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[124\]_B _287_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__544__B _544_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_506 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input190_A la_iena_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input288_A la_oenb_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_022_ _022_/A vssd vssd vccd vccd _022_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_6_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__560__A _560_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input455_A mprj_sel_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input51_A la_data_out_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1140 wire1141/X vssd vssd vccd vccd wire1140/X sky130_fd_sc_hd__buf_6
XFILLER_40_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1151 _349_/X vssd vssd vccd vccd wire1151/X sky130_fd_sc_hd__buf_6
Xwire1162 wire1163/X vssd vssd vccd vccd wire1162/X sky130_fd_sc_hd__buf_6
XFILLER_1_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1173 _338_/X vssd vssd vccd vccd wire1173/X sky130_fd_sc_hd__buf_6
XFILLER_40_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1184 wire1185/X vssd vssd vccd vccd wire1184/X sky130_fd_sc_hd__buf_6
XFILLER_1_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1195 _327_/X vssd vssd vccd vccd wire1195/X sky130_fd_sc_hd__buf_6
XANTENNA__438__C _438_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__454__B _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[115\]_B _278_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__486__A_N _614_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output841_A wire1047/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output939_A wire1166/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1472_A wire1473/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1716 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[24\]_A mprj_dat_i_user[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__364__B _364_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_B wire1251/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput104 la_data_out_mprj[75] vssd vssd vccd vccd _444_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput115 la_data_out_mprj[85] vssd vssd vccd vccd _454_/C sky130_fd_sc_hd__clkbuf_4
Xinput126 la_data_out_mprj[95] vssd vssd vccd vccd _464_/C sky130_fd_sc_hd__clkbuf_4
Xinput137 la_iena_mprj[104] vssd vssd vccd vccd _267_/B sky130_fd_sc_hd__clkbuf_4
Xinput148 la_iena_mprj[114] vssd vssd vccd vccd _277_/B sky130_fd_sc_hd__clkbuf_4
Xinput159 la_iena_mprj[124] vssd vssd vccd vccd _287_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__539__B _539_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[15\]_A mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_571_ _571_/A _571_/B vssd vssd vccd vccd _571_/X sky130_fd_sc_hd__and2_4
XFILLER_38_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input203_A la_iena_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__555__A _555_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__274__B _274_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input99_A la_data_out_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__290__A _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_005_ _005_/A vssd vssd vccd vccd _005_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__449__B _449_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output791_A _501_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1318_A wire1319/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output889_A wire969/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__184__B _184_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1687_A wire1688/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__359__B _359_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input153_A la_iena_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input320_A la_oenb_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input418_A mprj_adr_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_623_ _623_/A _623_/B vssd vssd vccd vccd _623_/X sky130_fd_sc_hd__and2_2
XFILLER_29_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input14_A la_data_out_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_554_ _554_/A _554_/B vssd vssd vccd vccd _554_/X sky130_fd_sc_hd__and2_4
XANTENNA__285__A _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_485_ _613_/A _485_/B _485_/C vssd vssd vccd vccd _485_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__451__C _451_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output637_A _009_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1170_A wire1171/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1268_A wire1268/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output804_A _558_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__179__B _179_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1435_A wire1435/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[51\] la_data_out_core[51] _214_/X vssd vssd vccd vccd _034_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_40_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1602_A wire1602/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__195__A _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput920 wire1142/X vssd vssd vccd vccd mprj_dat_o_user[16] sky130_fd_sc_hd__buf_8
XFILLER_2_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput931 wire1122/X vssd vssd vccd vccd mprj_dat_o_user[26] sky130_fd_sc_hd__buf_8
Xoutput942 wire1160/X vssd vssd vccd vccd mprj_dat_o_user[7] sky130_fd_sc_hd__buf_8
Xoutput953 wire1729/X vssd vssd vccd vccd user2_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_25_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A la_data_out_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1706 wire1706/A vssd vssd vccd vccd _463_/B sky130_fd_sc_hd__buf_6
XTAP_471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1717 wire1717/A vssd vssd vccd vccd _452_/B sky130_fd_sc_hd__buf_6
XFILLER_25_2987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1728 wire1728/A vssd vssd vccd vccd _441_/B sky130_fd_sc_hd__buf_6
XFILLER_3_3473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_270_ _270_/A _270_/B vssd vssd vccd vccd _270_/X sky130_fd_sc_hd__and2_1
XFILLER_41_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input270_A la_oenb_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input368_A la_oenb_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_606_ _606_/A _606_/B vssd vssd vccd vccd _606_/X sky130_fd_sc_hd__and2_4
XTAP_3573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_537_ _537_/A _537_/B vssd vssd vccd vccd _537_/X sky130_fd_sc_hd__and2_4
XTAP_2872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__446__C _446_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_468_ _596_/A _468_/B _468_/C vssd vssd vccd vccd _468_/X sky130_fd_sc_hd__and3b_4
XFILLER_14_983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output587_A wire1061/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_399_ _527_/A _399_/B _399_/C vssd vssd vccd vccd _399_/X sky130_fd_sc_hd__and3b_2
XFILLER_31_1712 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__462__B _462_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output754_A _513_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1385_A wire1385/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output921_A wire1140/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[99\] la_data_out_core[99] wire1258/X vssd vssd vccd vccd _082_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_29_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2206 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1552_A wire1553/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__372__B _372_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[7\]_A mprj_dat_i_user[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput750 _509_/X vssd vssd vccd vccd la_oenb_core[12] sky130_fd_sc_hd__buf_8
XFILLER_25_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput761 _519_/X vssd vssd vccd vccd la_oenb_core[22] sky130_fd_sc_hd__buf_8
XFILLER_21_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput772 _529_/X vssd vssd vccd vccd la_oenb_core[32] sky130_fd_sc_hd__buf_8
Xoutput783 _539_/X vssd vssd vccd vccd la_oenb_core[42] sky130_fd_sc_hd__buf_8
XFILLER_40_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput794 _549_/X vssd vssd vccd vccd la_oenb_core[52] sky130_fd_sc_hd__buf_8
XFILLER_43_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1503 wire1503/A vssd vssd vccd vccd _267_/A sky130_fd_sc_hd__buf_6
XFILLER_5_2845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1026 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1514 wire1514/A vssd vssd vccd vccd _256_/A sky130_fd_sc_hd__buf_4
XFILLER_21_3349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1525 wire1525/A vssd vssd vccd vccd _189_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1536 wire1536/A vssd vssd vccd vccd _178_/A sky130_fd_sc_hd__buf_6
XANTENNA_user_to_mprj_in_gates\[7\]_A la_data_out_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1547 wire1547/A vssd vssd vccd vccd _167_/A sky130_fd_sc_hd__buf_6
XFILLER_21_2648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1558 wire1559/X vssd vssd vccd vccd _621_/B sky130_fd_sc_hd__buf_6
Xwire1569 wire1569/A vssd vssd vccd vccd wire1569/X sky130_fd_sc_hd__buf_6
XFILLER_46_349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__547__B _547_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input116_A la_data_out_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_322_ _322_/A _322_/B vssd vssd vccd vccd _322_/X sky130_fd_sc_hd__and2_4
XTAP_1467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__563__A _563_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_253_ _253_/A _253_/B vssd vssd vccd vccd _253_/X sky130_fd_sc_hd__and2_4
XFILLER_14_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__282__B _282_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input81_A la_data_out_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_184_ _184_/A _184_/B vssd vssd vccd vccd _184_/X sky130_fd_sc_hd__and2_1
XFILLER_11_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output502_A _370_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__457__B _457_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1133_A _358_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1300_A wire1301/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output871_A wire1178/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3676 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[14\] la_data_out_core[14] _177_/X vssd vssd vccd vccd _161_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_31_2210 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[27\] mprj_dat_i_user[27] rebuffer6/X vssd vssd vccd vccd wire1006/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_33_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3811 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1914 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[125\] la_data_out_core[125] _288_/X vssd vssd vccd vccd _108_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_5_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__367__B _367_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3418 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__392__A_N _520_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_rebuffer4_A split13/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput580 wire1066/X vssd vssd vccd vccd la_data_in_core[90] sky130_fd_sc_hd__buf_8
XFILLER_40_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput591 _147_/Y vssd vssd vccd vccd la_data_in_mprj[0] sky130_fd_sc_hd__buf_8
XFILLER_43_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1300 wire1301/X vssd vssd vccd vccd _365_/B sky130_fd_sc_hd__buf_6
XFILLER_5_3387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1311 wire1311/A vssd vssd vccd vccd wire1311/X sky130_fd_sc_hd__buf_6
XFILLER_25_2581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1322 wire1323/X vssd vssd vccd vccd _355_/B sky130_fd_sc_hd__buf_6
Xwire1333 wire1333/A vssd vssd vccd vccd wire1333/X sky130_fd_sc_hd__buf_6
XANTENNA_input233_A la_iena_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1344 wire1345/X vssd vssd vccd vccd _314_/B sky130_fd_sc_hd__buf_6
XFILLER_46_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1355 wire1356/X vssd vssd vccd vccd wire1355/X sky130_fd_sc_hd__buf_6
XANTENNA__558__A _558_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1366 wire1366/A vssd vssd vccd vccd wire1366/X sky130_fd_sc_hd__buf_6
XFILLER_46_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1377 wire1377/A vssd vssd vccd vccd wire1377/X sky130_fd_sc_hd__buf_6
XFILLER_19_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1388 wire1388/A vssd vssd vccd vccd wire1388/X sky130_fd_sc_hd__buf_6
XFILLER_35_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1399 wire1400/X vssd vssd vccd vccd _322_/B sky130_fd_sc_hd__buf_6
XFILLER_28_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input400_A mprj_adr_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__277__B _277_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__293__A _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_305_ _305_/A _305_/B vssd vssd vccd vccd _305_/X sky130_fd_sc_hd__and2_4
XFILLER_15_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_236_ _236_/A _236_/B vssd vssd vccd vccd _236_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_167_ _167_/A _167_/B vssd vssd vccd vccd _167_/X sky130_fd_sc_hd__and2_4
XFILLER_6_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_098_ _098_/A vssd vssd vccd vccd _098_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output717_A wire990/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1348_A wire1348/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__187__B _187_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_382 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire968_A _132_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1722 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput308 la_oenb_mprj[28] vssd vssd vccd vccd _525_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput319 la_oenb_mprj[38] vssd vssd vccd vccd _535_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_518 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_021_ _021_/A vssd vssd vccd vccd _021_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input183_A la_iena_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__560__B _560_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input350_A la_oenb_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input448_A mprj_dat_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input44_A la_data_out_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1130 wire1131/X vssd vssd vccd vccd wire1130/X sky130_fd_sc_hd__buf_6
XANTENNA__288__A _288_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1141 _354_/X vssd vssd vccd vccd wire1141/X sky130_fd_sc_hd__buf_6
XFILLER_40_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1152 wire1153/X vssd vssd vccd vccd wire1152/X sky130_fd_sc_hd__buf_6
XFILLER_38_4141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1163 _343_/X vssd vssd vccd vccd wire1163/X sky130_fd_sc_hd__buf_6
XFILLER_19_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1174 wire1175/X vssd vssd vccd vccd wire1174/X sky130_fd_sc_hd__buf_6
XFILLER_21_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1185 _332_/X vssd vssd vccd vccd wire1185/X sky130_fd_sc_hd__buf_6
XFILLER_34_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1196 _326_/X vssd vssd vccd vccd wire1196/X sky130_fd_sc_hd__buf_6
XFILLER_35_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__454__C _454_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output667_A _036_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_219_ _219_/A _219_/B vssd vssd vccd vccd _219_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1298_A wire1299/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__470__B _470_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output834_A _586_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1465_A wire1465/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[81\] la_data_out_core[81] _244_/X vssd vssd vccd vccd _064_/A
+ sky130_fd_sc_hd__nand2_8
XTAP_823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__198__A _198_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[24\]_B split13/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3502 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__430__A_N _558_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__380__B _380_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput105 la_data_out_mprj[76] vssd vssd vccd vccd _445_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput116 la_data_out_mprj[86] vssd vssd vccd vccd _455_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_44_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput127 la_data_out_mprj[96] vssd vssd vccd vccd _465_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput138 la_iena_mprj[105] vssd vssd vccd vccd _268_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput149 la_iena_mprj[115] vssd vssd vccd vccd _278_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_570_ _570_/A _570_/B vssd vssd vccd vccd _570_/X sky130_fd_sc_hd__and2_4
XFILLER_0_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__555__B _555_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input398_A mprj_adr_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__571__A _571_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_004_ _004_/A vssd vssd vccd vccd _004_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2738 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__449__C _449_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_gates\[0\]_A user_irq_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__465__B _465_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1213_A wire1214/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__453__A_N _581_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output784_A _540_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output951_A wire1467/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1582_A wire1582/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__375__B _375_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input146_A la_iena_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_622_ _622_/A _622_/B vssd vssd vccd vccd _622_/X sky130_fd_sc_hd__and2_2
XANTENNA_input313_A la_oenb_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__476__A_N _604_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__566__A _566_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_553_ _553_/A _553_/B vssd vssd vccd vccd _553_/X sky130_fd_sc_hd__and2_1
XFILLER_26_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_484_ _612_/A _484_/B _484_/C vssd vssd vccd vccd _484_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output532_A wire1088/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1163_A _343_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1330_A wire1331/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1428_A wire1428/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[44\] la_data_out_core[44] _207_/X vssd vssd vccd vccd _027_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_24_918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput910 wire979/X vssd vssd vccd vccd mprj_dat_i_core[7] sky130_fd_sc_hd__buf_8
Xoutput921 wire1140/X vssd vssd vccd vccd mprj_dat_o_user[17] sky130_fd_sc_hd__buf_8
Xoutput932 wire1120/X vssd vssd vccd vccd mprj_dat_o_user[27] sky130_fd_sc_hd__buf_8
Xoutput943 wire1158/X vssd vssd vccd vccd mprj_dat_o_user[8] sky130_fd_sc_hd__buf_8
XFILLER_9_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[6\] la_data_out_core[6] _169_/X vssd vssd vccd vccd _153_/A
+ sky130_fd_sc_hd__nand2_1
Xoutput954 output954/A vssd vssd vccd vccd user2_vdd_powergood sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[30\]_A la_data_out_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1707 wire1707/A vssd vssd vccd vccd _462_/B sky130_fd_sc_hd__buf_6
XFILLER_28_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1718 wire1718/A vssd vssd vccd vccd _451_/B sky130_fd_sc_hd__buf_6
XTAP_472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1729 wire1730/X vssd vssd vccd vccd wire1729/X sky130_fd_sc_hd__buf_6
XTAP_494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_A la_data_out_core[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input263_A la_oenb_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[21\]_A la_data_out_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input430_A mprj_dat_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__296__A _296_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_605_ _605_/A _605_/B vssd vssd vccd vccd _605_/X sky130_fd_sc_hd__and2_2
XTAP_3574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_536_ _536_/A _536_/B vssd vssd vccd vccd _536_/X sky130_fd_sc_hd__and2_4
XTAP_2862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[88\]_A la_data_out_core[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_467_ _595_/A _467_/B _467_/C vssd vssd vccd vccd _467_/X sky130_fd_sc_hd__and3b_2
XFILLER_31_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_398_ _526_/A _398_/B _398_/C vssd vssd vccd vccd _398_/X sky130_fd_sc_hd__and3b_2
XANTENNA_output482_A _486_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1009_A wire1009/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__462__C _462_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1768 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output747_A wire1034/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1280_A wire1281/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1378_A wire1379/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2218 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output914_A wire1154/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[12\]_A la_data_out_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1545_A wire1545/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1712_A wire1712/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire998_A wire998/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[79\]_A la_data_out_core[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1056 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_2509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__372__C _372_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput740 wire1038/X vssd vssd vccd vccd la_oenb_core[119] sky130_fd_sc_hd__buf_8
Xoutput751 _510_/X vssd vssd vccd vccd la_oenb_core[13] sky130_fd_sc_hd__buf_8
Xoutput762 _520_/X vssd vssd vccd vccd la_oenb_core[23] sky130_fd_sc_hd__buf_8
XFILLER_5_3514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput773 _530_/X vssd vssd vccd vccd la_oenb_core[33] sky130_fd_sc_hd__buf_8
XFILLER_9_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput784 _540_/X vssd vssd vccd vccd la_oenb_core[43] sky130_fd_sc_hd__buf_8
XFILLER_40_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput795 _550_/X vssd vssd vccd vccd la_oenb_core[53] sky130_fd_sc_hd__buf_8
XFILLER_5_2802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1504 wire1504/A vssd vssd vccd vccd _266_/A sky130_fd_sc_hd__buf_6
XFILLER_21_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1515 wire1515/A vssd vssd vccd vccd _253_/A sky130_fd_sc_hd__buf_6
XFILLER_41_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1526 wire1526/A vssd vssd vccd vccd _188_/A sky130_fd_sc_hd__buf_6
XTAP_280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1537 wire1537/A vssd vssd vccd vccd _177_/A sky130_fd_sc_hd__buf_6
XANTENNA_user_to_mprj_in_gates\[7\]_B _170_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1548 wire1548/A vssd vssd vccd vccd _166_/A sky130_fd_sc_hd__buf_6
Xwire1559 wire1559/A vssd vssd vccd vccd wire1559/X sky130_fd_sc_hd__buf_6
XFILLER_41_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input109_A la_data_out_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_321_ _321_/A _321_/B vssd vssd vccd vccd _321_/X sky130_fd_sc_hd__and2_4
XFILLER_19_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_252_ _252_/A _252_/B vssd vssd vccd vccd _252_/X sky130_fd_sc_hd__and2_4
XANTENNA__563__B _563_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_183_ _183_/A _183_/B vssd vssd vccd vccd _183_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input380_A la_oenb_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input74_A la_data_out_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__457__C _457_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1126_A wire1127/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output697_A _063_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_519_ _519_/A _519_/B vssd vssd vccd vccd _519_/X sky130_fd_sc_hd__and2_4
XFILLER_37_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__473__B _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2222 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output864_A wire1190/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1495_A wire1495/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1662_A wire1663/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3823 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1494 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[118\] la_data_out_core[118] _281_/X vssd vssd vccd vccd _101_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_3_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__383__B _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput570 _450_/X vssd vssd vccd vccd la_data_in_core[81] sky130_fd_sc_hd__buf_8
Xoutput581 wire1065/X vssd vssd vccd vccd la_data_in_core[91] sky130_fd_sc_hd__buf_8
XFILLER_25_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput592 wire989/X vssd vssd vccd vccd la_data_in_mprj[100] sky130_fd_sc_hd__buf_8
XFILLER_43_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1301 wire1301/A vssd vssd vccd vccd wire1301/X sky130_fd_sc_hd__buf_6
XFILLER_8_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1312 wire1313/X vssd vssd vccd vccd _359_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2643 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1323 wire1323/A vssd vssd vccd vccd wire1323/X sky130_fd_sc_hd__buf_6
XFILLER_5_3399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1334 wire1335/X vssd vssd vccd vccd _349_/B sky130_fd_sc_hd__buf_6
Xwire1345 wire1345/A vssd vssd vccd vccd wire1345/X sky130_fd_sc_hd__buf_6
XFILLER_8_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1356 wire1356/A vssd vssd vccd vccd wire1356/X sky130_fd_sc_hd__buf_6
XFILLER_5_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__558__B _558_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input226_A la_iena_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1367 wire1368/X vssd vssd vccd vccd _307_/B sky130_fd_sc_hd__buf_6
XFILLER_21_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1378 wire1379/X vssd vssd vccd vccd _330_/B sky130_fd_sc_hd__buf_6
XFILLER_46_147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1389 wire1390/X vssd vssd vccd vccd _325_/B sky130_fd_sc_hd__buf_6
XFILLER_34_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[127\]_A la_data_out_core[127] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__574__A _574_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_304_ _304_/A _304_/B vssd vssd vccd vccd _304_/X sky130_fd_sc_hd__and2_4
XANTENNA__293__B _293_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_235_ _235_/A _235_/B vssd vssd vccd vccd _235_/X sky130_fd_sc_hd__and2_4
XFILLER_6_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_166_ _166_/A _166_/B vssd vssd vccd vccd _166_/X sky130_fd_sc_hd__and2_4
XFILLER_32_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_097_ _097_/A vssd vssd vccd vccd _097_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_6_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output612_A _102_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__468__B _468_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1410_A wire1411/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_394 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1508_A wire1508/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_A la_data_out_core[118] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_15_3452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1162 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput309 la_oenb_mprj[29] vssd vssd vccd vccd _526_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1734 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__378__B _378_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[109\]_A la_data_out_core[109] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_25_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_020_ _020_/A vssd vssd vccd vccd _020_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input176_A la_iena_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input343_A la_oenb_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__569__A _569_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input37_A la_data_out_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1120 wire1121/X vssd vssd vccd vccd wire1120/X sky130_fd_sc_hd__buf_6
Xwire1131 _359_/X vssd vssd vccd vccd wire1131/X sky130_fd_sc_hd__buf_6
XFILLER_1_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1142 wire1143/X vssd vssd vccd vccd wire1142/X sky130_fd_sc_hd__buf_6
XFILLER_19_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1153 _348_/X vssd vssd vccd vccd wire1153/X sky130_fd_sc_hd__buf_6
XFILLER_40_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1164 wire1165/X vssd vssd vccd vccd wire1164/X sky130_fd_sc_hd__buf_6
Xwire1175 _337_/X vssd vssd vccd vccd wire1175/X sky130_fd_sc_hd__buf_6
Xwire1186 wire1187/X vssd vssd vccd vccd wire1186/X sky130_fd_sc_hd__buf_6
XFILLER_1_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1197 wire1198/X vssd vssd vccd vccd wire1197/X sky130_fd_sc_hd__buf_6
XFILLER_34_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_218_ _218_/A _218_/B vssd vssd vccd vccd _218_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output562_A _443_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_149_ _149_/A vssd vssd vccd vccd _149_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_13_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__470__C _470_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1193_A _328_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3467 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output827_A _579_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__382__A_N _510_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1360_A wire1361/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1458_A wire1459/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[74\] la_data_out_core[74] _237_/X vssd vssd vccd vccd _057_/A
+ sky130_fd_sc_hd__nand2_8
XTAP_879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1625_A wire1625/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_824 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire980_A _120_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__380__C _380_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput106 la_data_out_mprj[77] vssd vssd vccd vccd _446_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_41_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput117 la_data_out_mprj[87] vssd vssd vccd vccd _456_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput128 la_data_out_mprj[97] vssd vssd vccd vccd _466_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput139 la_iena_mprj[106] vssd vssd vccd vccd _269_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input293_A la_oenb_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__571__B _571_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_90 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_003_ _003_/A vssd vssd vccd vccd _003_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input460_A user_irq_ena[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__299__A _299_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_irq_gates\[0\]_B _291_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__465__C _465_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1206_A _319_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output777_A _534_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_698 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__481__B _481_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output944_A wire1156/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1575_A wire1575/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[100\] la_data_out_core[100] wire1257/X vssd vssd vccd vccd
+ _083_/A sky130_fd_sc_hd__nand2_4
XFILLER_27_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__375__C _375_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__391__B _391_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_4005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2614 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input139_A la_iena_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_621_ _621_/A _621_/B vssd vssd vccd vccd _621_/X sky130_fd_sc_hd__and2_1
XFILLER_35_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_552_ _552_/A _552_/B vssd vssd vccd vccd _552_/X sky130_fd_sc_hd__and2_4
XANTENNA__566__B _566_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input306_A la_oenb_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1110 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_483_ _611_/A _483_/B _483_/C vssd vssd vccd vccd _483_/X sky130_fd_sc_hd__and3b_4
XFILLER_26_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__582__A _582_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output525_A wire1095/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1156_A wire1157/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__420__A_N _548_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__476__B _476_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1323_A wire1323/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output894_A wire965/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[37\] la_data_out_core[37] _200_/X vssd vssd vccd vccd _020_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_36_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput900 _141_/Y vssd vssd vccd vccd mprj_dat_i_core[27] sky130_fd_sc_hd__buf_8
Xoutput911 wire978/X vssd vssd vccd vccd mprj_dat_i_core[8] sky130_fd_sc_hd__buf_8
XFILLER_9_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput922 wire1138/X vssd vssd vccd vccd mprj_dat_o_user[18] sky130_fd_sc_hd__buf_8
Xoutput933 wire1118/X vssd vssd vccd vccd mprj_dat_o_user[28] sky130_fd_sc_hd__buf_8
Xoutput944 wire1156/X vssd vssd vccd vccd mprj_dat_o_user[9] sky130_fd_sc_hd__buf_8
Xoutput955 wire1242/X vssd vssd vccd vccd user_clock sky130_fd_sc_hd__buf_8
XFILLER_9_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1708 wire1708/A vssd vssd vccd vccd _461_/B sky130_fd_sc_hd__buf_6
XTAP_473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1719 wire1719/A vssd vssd vccd vccd _450_/B sky130_fd_sc_hd__buf_6
XFILLER_45_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__386__B _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_930 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_B _260_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3174 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input256_A la_iena_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__443__A_N _571_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input423_A mprj_dat_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__577__A _577_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__296__B _296_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_604_ _604_/A _604_/B vssd vssd vccd vccd _604_/X sky130_fd_sc_hd__and2_4
XTAP_3553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_535_ _535_/A _535_/B vssd vssd vccd vccd _535_/X sky130_fd_sc_hd__and2_4
XFILLER_33_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[88\]_B _251_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_466_ _594_/A _466_/B _466_/C vssd vssd vccd vccd _466_/X sky130_fd_sc_hd__and3b_2
XFILLER_35_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_397_ _525_/A _397_/B _397_/C vssd vssd vccd vccd _397_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output475_A _479_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1168 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output642_A _013_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1273_A wire1274/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[12\]_B _175_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1518 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output907_A wire982/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1440_A wire1441/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1538_A wire1538/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1705_A wire1705/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[79\]_B _242_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__466__A_N _594_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput730 _507_/X vssd vssd vccd vccd la_oenb_core[10] sky130_fd_sc_hd__buf_8
Xoutput741 _508_/X vssd vssd vccd vccd la_oenb_core[11] sky130_fd_sc_hd__buf_8
Xoutput752 _511_/X vssd vssd vccd vccd la_oenb_core[14] sky130_fd_sc_hd__buf_8
Xoutput763 _521_/X vssd vssd vccd vccd la_oenb_core[24] sky130_fd_sc_hd__buf_8
Xoutput774 _531_/X vssd vssd vccd vccd la_oenb_core[34] sky130_fd_sc_hd__buf_8
Xoutput785 _541_/X vssd vssd vccd vccd la_oenb_core[44] sky130_fd_sc_hd__buf_8
Xoutput796 _551_/X vssd vssd vccd vccd la_oenb_core[54] sky130_fd_sc_hd__buf_8
XFILLER_5_3559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1505 wire1505/A vssd vssd vccd vccd _265_/A sky130_fd_sc_hd__buf_6
XFILLER_5_2858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1516 wire1516/A vssd vssd vccd vccd _252_/A sky130_fd_sc_hd__buf_6
XFILLER_21_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1527 wire1527/A vssd vssd vccd vccd _187_/A sky130_fd_sc_hd__buf_6
XFILLER_41_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1538 wire1538/A vssd vssd vccd vccd _176_/A sky130_fd_sc_hd__buf_6
Xwire1549 wire1549/A vssd vssd vccd vccd _165_/A sky130_fd_sc_hd__buf_6
XFILLER_21_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_320_ _320_/A _320_/B vssd vssd vccd vccd _320_/X sky130_fd_sc_hd__and2_4
XFILLER_42_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_251_ _251_/A _251_/B vssd vssd vccd vccd _251_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_182_ _182_/A _182_/B vssd vssd vccd vccd _182_/X sky130_fd_sc_hd__and2_4
XFILLER_13_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input373_A la_oenb_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input67_A la_data_out_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__100__A _100_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_518_ _518_/A _518_/B vssd vssd vccd vccd _518_/X sky130_fd_sc_hd__and2_4
XFILLER_18_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1021_A wire1021/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output592_A wire989/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1119_A _365_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__473__C _473_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_449_ _577_/A _449_/B _449_/C vssd vssd vccd vccd _449_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__489__A_N _617_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output857_A wire1201/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1390_A wire1390/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3307 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1655_A wire1655/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3879 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__010__A _010_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__383__C _383_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput560 _441_/X vssd vssd vccd vccd la_data_in_core[72] sky130_fd_sc_hd__buf_8
XFILLER_40_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput571 _451_/X vssd vssd vccd vccd la_data_in_core[82] sky130_fd_sc_hd__buf_8
XFILLER_43_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput582 wire1064/X vssd vssd vccd vccd la_data_in_core[92] sky130_fd_sc_hd__buf_8
Xoutput593 wire988/X vssd vssd vccd vccd la_data_in_mprj[101] sky130_fd_sc_hd__buf_8
XFILLER_5_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1302 wire1303/X vssd vssd vccd vccd _364_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1313 wire1313/A vssd vssd vccd vccd wire1313/X sky130_fd_sc_hd__buf_6
XFILLER_8_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1324 wire1325/X vssd vssd vccd vccd _354_/B sky130_fd_sc_hd__buf_6
Xwire1335 wire1335/A vssd vssd vccd vccd wire1335/X sky130_fd_sc_hd__buf_6
XFILLER_1_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1702 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1346 wire1347/X vssd vssd vccd vccd _313_/B sky130_fd_sc_hd__buf_6
Xwire1357 wire1358/X vssd vssd vccd vccd _309_/B sky130_fd_sc_hd__buf_6
XFILLER_3_3091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1368 wire1369/X vssd vssd vccd vccd wire1368/X sky130_fd_sc_hd__buf_6
Xwire1379 wire1379/A vssd vssd vccd vccd wire1379/X sky130_fd_sc_hd__buf_6
XANTENNA_input121_A la_data_out_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input219_A la_iena_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[127\]_B _290_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__574__B _574_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_303_ _303_/A _303_/B vssd vssd vccd vccd _303_/X sky130_fd_sc_hd__and2_4
XTAP_1288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_234_ _234_/A _234_/B vssd vssd vccd vccd _234_/X sky130_fd_sc_hd__and2_4
XFILLER_7_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__590__A _590_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_165_ _165_/A _165_/B vssd vssd vccd vccd _165_/X sky130_fd_sc_hd__and2_2
XFILLER_6_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[2\] mprj_dat_i_user[2] max_cap1244/X vssd vssd vccd vccd wire1001/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_13_1263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_096_ _096_/A vssd vssd vccd vccd _096_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_6_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_powergood_check_mprj_vdd_logic1 output952/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__468__C _468_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output605_A _095_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1236_A _300_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_800 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__484__B _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_B _281_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2307 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1174 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__005__A _005_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3643 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1746 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[27\]_A mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__378__C _378_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__394__B _394_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[109\]_B _272_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input169_A la_iena_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__569__B _569_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input336_A la_oenb_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[18\]_A mprj_dat_i_user[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1110 _377_/X vssd vssd vccd vccd wire1110/X sky130_fd_sc_hd__buf_6
XFILLER_5_3197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1121 _364_/X vssd vssd vccd vccd wire1121/X sky130_fd_sc_hd__buf_6
XFILLER_25_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1132 wire1133/X vssd vssd vccd vccd wire1132/X sky130_fd_sc_hd__buf_6
XFILLER_1_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1143 _353_/X vssd vssd vccd vccd wire1143/X sky130_fd_sc_hd__buf_6
Xwire1154 wire1155/X vssd vssd vccd vccd wire1154/X sky130_fd_sc_hd__buf_6
XFILLER_43_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1165 _342_/X vssd vssd vccd vccd wire1165/X sky130_fd_sc_hd__buf_6
Xwire1176 wire1177/X vssd vssd vccd vccd wire1176/X sky130_fd_sc_hd__buf_6
Xwire1187 _331_/X vssd vssd vccd vccd wire1187/X sky130_fd_sc_hd__buf_6
Xwire1198 _325_/X vssd vssd vccd vccd wire1198/X sky130_fd_sc_hd__buf_6
XFILLER_34_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__585__A _585_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1358 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_217_ _217_/A _217_/B vssd vssd vccd vccd _217_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_148_ _148_/A vssd vssd vccd vccd _148_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output555_A wire1070/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2682 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_079_ _079_/A vssd vssd vccd vccd _079_/Y sky130_fd_sc_hd__inv_4
XANTENNA_wire1186_A wire1187/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3700 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output722_A _599_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__479__B _479_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1353_A wire1353/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[67\] la_data_out_core[67] _230_/X vssd vssd vccd vccd _050_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_22_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire973_A _127_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput107 la_data_out_mprj[78] vssd vssd vccd vccd _447_/C sky130_fd_sc_hd__clkbuf_4
Xinput118 la_data_out_mprj[88] vssd vssd vccd vccd _457_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__389__B _389_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1554 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput129 la_data_out_mprj[98] vssd vssd vccd vccd _467_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input286_A la_oenb_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_80 _169_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_390 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_002_ _002_/A vssd vssd vccd vccd _002_/Y sky130_fd_sc_hd__inv_2
XANTENNA_91 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input453_A mprj_iena_wb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__299__B _299_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__481__C _481_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output937_A wire1112/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1470_A wire1471/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1568_A wire1569/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__391__C _391_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_620_ _620_/A _620_/B vssd vssd vccd vccd _620_/X sky130_fd_sc_hd__and2_2
XTAP_3713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_551_ _551_/A _551_/B vssd vssd vccd vccd _551_/X sky130_fd_sc_hd__and2_4
XFILLER_44_224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input201_A la_iena_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_482_ _610_/A _482_/B _482_/C vssd vssd vccd vccd _482_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1122 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__372__A_N _500_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__582__B _582_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input97_A la_data_out_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__103__A _103_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output518_A wire1101/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput460 user_irq_ena[0] vssd vssd vccd vccd wire1264/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1149_A _350_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__476__C _476_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1316_A wire1317/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output887_A wire971/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__492__B _492_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1685_A wire1685/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput901 _142_/Y vssd vssd vccd vccd mprj_dat_i_core[28] sky130_fd_sc_hd__buf_8
Xoutput912 wire977/X vssd vssd vccd vccd mprj_dat_i_core[9] sky130_fd_sc_hd__buf_8
Xoutput923 wire1136/X vssd vssd vccd vccd mprj_dat_o_user[19] sky130_fd_sc_hd__buf_8
XFILLER_9_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput934 wire1116/X vssd vssd vccd vccd mprj_dat_o_user[29] sky130_fd_sc_hd__buf_8
XFILLER_28_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput945 wire1233/X vssd vssd vccd vccd mprj_sel_o_user[0] sky130_fd_sc_hd__buf_8
Xoutput956 wire1241/X vssd vssd vccd vccd user_clock2 sky130_fd_sc_hd__buf_8
XFILLER_9_3888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__013__A _013_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1709 wire1709/A vssd vssd vccd vccd _460_/B sky130_fd_sc_hd__buf_6
XFILLER_23_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__386__C _386_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__395__A_N _523_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3310 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input151_A la_iena_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input249_A la_iena_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__577__B _577_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input416_A mprj_adr_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_603_ _603_/A _603_/B vssd vssd vccd vccd _603_/X sky130_fd_sc_hd__and2_4
XTAP_3543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input12_A la_data_out_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_534_ _534_/A _534_/B vssd vssd vccd vccd _534_/X sky130_fd_sc_hd__and2_4
XTAP_2842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__593__A _593_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_465_ _593_/A _465_/B _465_/C vssd vssd vccd vccd _465_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_396_ _524_/A _396_/B _396_/C vssd vssd vccd vccd _396_/X sky130_fd_sc_hd__and3b_2
XFILLER_43_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output468_A _473_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output635_A _007_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1266_A wire1266/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output802_A _502_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3774 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1210 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__487__B _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1433_A wire1433/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput290 la_oenb_mprj[127] vssd vssd vccd vccd _624_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1600_A wire1601/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__008__A _008_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput720 wire1046/X vssd vssd vccd vccd la_oenb_core[100] sky130_fd_sc_hd__buf_8
Xoutput731 wire1042/X vssd vssd vccd vccd la_oenb_core[110] sky130_fd_sc_hd__buf_8
XFILLER_9_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput742 _617_/X vssd vssd vccd vccd la_oenb_core[120] sky130_fd_sc_hd__buf_8
Xoutput753 _512_/X vssd vssd vccd vccd la_oenb_core[15] sky130_fd_sc_hd__buf_8
XFILLER_43_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput764 _522_/X vssd vssd vccd vccd la_oenb_core[25] sky130_fd_sc_hd__buf_8
XFILLER_25_3455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput775 _532_/X vssd vssd vccd vccd la_oenb_core[35] sky130_fd_sc_hd__buf_8
XFILLER_9_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput786 wire1052/X vssd vssd vccd vccd la_oenb_core[45] sky130_fd_sc_hd__buf_8
Xoutput797 _552_/X vssd vssd vccd vccd la_oenb_core[55] sky130_fd_sc_hd__buf_8
XFILLER_25_2732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A la_data_out_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1506 wire1506/A vssd vssd vccd vccd _264_/A sky130_fd_sc_hd__buf_6
XFILLER_8_1259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1517 wire1517/A vssd vssd vccd vccd _250_/A sky130_fd_sc_hd__buf_6
XTAP_271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1528 wire1528/A vssd vssd vccd vccd _186_/A sky130_fd_sc_hd__buf_6
XTAP_282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1539 wire1539/A vssd vssd vccd vccd _175_/A sky130_fd_sc_hd__buf_6
XANTENNA__397__B _397_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_250_ _250_/A _250_/B vssd vssd vccd vccd _250_/X sky130_fd_sc_hd__and2_4
XFILLER_23_761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_181_ _181_/A _181_/B vssd vssd vccd vccd _181_/X sky130_fd_sc_hd__and2_2
XFILLER_10_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input199_A la_iena_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__410__A_N _538_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input366_A la_oenb_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_irq_gates\[1\] user_irq_core[1] _292_/X vssd vssd vccd vccd _112_/A sky130_fd_sc_hd__nand2_2
XFILLER_8_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__588__A _588_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_517_ _517_/A _517_/B vssd vssd vccd vccd _517_/X sky130_fd_sc_hd__and2_4
XTAP_2672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_448_ _576_/A _448_/B _448_/C vssd vssd vccd vccd _448_/X sky130_fd_sc_hd__and3b_4
XTAP_1982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1014_A wire1014/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output585_A wire1062/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_379_ _507_/A _379_/B _379_/C vssd vssd vccd vccd _379_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output752_A _511_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1383_A wire1383/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3319 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[97\] la_data_out_core[97] _260_/X vssd vssd vccd vccd _080_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_46_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1550_A wire1550/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1648_A wire1648/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__498__A _498_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__433__A_N _561_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput550 _432_/X vssd vssd vccd vccd la_data_in_core[63] sky130_fd_sc_hd__buf_8
Xoutput561 _442_/X vssd vssd vccd vccd la_data_in_core[73] sky130_fd_sc_hd__buf_8
XFILLER_25_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput572 _452_/X vssd vssd vccd vccd la_data_in_core[83] sky130_fd_sc_hd__buf_8
XFILLER_40_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput583 _462_/X vssd vssd vccd vccd la_data_in_core[93] sky130_fd_sc_hd__buf_8
XFILLER_5_3335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput594 wire987/X vssd vssd vccd vccd la_data_in_mprj[102] sky130_fd_sc_hd__buf_8
XFILLER_5_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1303 wire1303/A vssd vssd vccd vccd wire1303/X sky130_fd_sc_hd__buf_6
XFILLER_43_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1314 wire1315/X vssd vssd vccd vccd _358_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__201__A _201_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1325 wire1325/A vssd vssd vccd vccd wire1325/X sky130_fd_sc_hd__buf_6
XFILLER_5_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1336 wire1337/X vssd vssd vccd vccd _348_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1347 wire1348/X vssd vssd vccd vccd wire1347/X sky130_fd_sc_hd__buf_6
XFILLER_3_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1358 wire1359/X vssd vssd vccd vccd wire1358/X sky130_fd_sc_hd__buf_6
Xwire1369 wire1369/A vssd vssd vccd vccd wire1369/X sky130_fd_sc_hd__buf_6
XFILLER_38_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input114_A la_data_out_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_302_ _302_/A _302_/B vssd vssd vccd vccd _302_/X sky130_fd_sc_hd__and2_4
XTAP_1278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_233_ _233_/A _233_/B vssd vssd vccd vccd _233_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__590__B _590_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_164_ _164_/A _164_/B vssd vssd vccd vccd _164_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_095_ _095_/A vssd vssd vccd vccd _095_/Y sky130_fd_sc_hd__inv_4
XFILLER_40_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output500_A _387_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1131_A _359_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__456__A_N _584_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1229_A wire1230/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__484__C _484_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_170 _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[12\] la_data_out_core[12] _175_/X vssd vssd vccd vccd _159_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_33_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[25\] mprj_dat_i_user[25] rebuffer8/X vssd vssd vccd vccd wire1009/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_18_1186 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1598_A wire1598/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3699 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__021__A _021_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[123\] la_data_out_core[123] _286_/X vssd vssd vccd vccd _106_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_29_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__394__C _394_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2971 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1100 _404_/X vssd vssd vccd vccd wire1100/X sky130_fd_sc_hd__buf_6
XFILLER_40_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1111 _375_/X vssd vssd vccd vccd wire1111/X sky130_fd_sc_hd__buf_6
XFILLER_27_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1122 wire1123/X vssd vssd vccd vccd wire1122/X sky130_fd_sc_hd__buf_6
XFILLER_43_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input231_A la_iena_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1133 _358_/X vssd vssd vccd vccd wire1133/X sky130_fd_sc_hd__buf_6
XANTENNA_input329_A la_oenb_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__479__A_N _607_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1144 wire1145/X vssd vssd vccd vccd wire1144/X sky130_fd_sc_hd__buf_6
Xwire1155 _347_/X vssd vssd vccd vccd wire1155/X sky130_fd_sc_hd__buf_6
XFILLER_38_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1166 wire1167/X vssd vssd vccd vccd wire1166/X sky130_fd_sc_hd__buf_6
XFILLER_1_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1177 _336_/X vssd vssd vccd vccd wire1177/X sky130_fd_sc_hd__buf_6
XFILLER_35_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1188 wire1189/X vssd vssd vccd vccd wire1188/X sky130_fd_sc_hd__buf_6
Xwire1199 wire1200/X vssd vssd vccd vccd wire1199/X sky130_fd_sc_hd__buf_6
XFILLER_38_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__585__B _585_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_216_ _216_/A _216_/B vssd vssd vccd vccd _216_/X sky130_fd_sc_hd__and2_4
XFILLER_11_594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__106__A _106_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_147_ _147_/A vssd vssd vccd vccd _147_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_078_ _078_/A vssd vssd vccd vccd _078_/Y sky130_fd_sc_hd__inv_4
XANTENNA_output548_A wire1074/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1179_A _335_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3756 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__479__C _479_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output715_A _080_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1346_A wire1347/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__495__B _495_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1054 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__016__A _016_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[60\]_A la_data_out_core[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput108 la_data_out_mprj[79] vssd vssd vccd vccd _448_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__389__C _389_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput119 la_data_out_mprj[89] vssd vssd vccd vccd _458_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_41_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1566 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_686 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_70 _250_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_81 _169_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_001_ _001_/A vssd vssd vccd vccd _001_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_92 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input181_A la_iena_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input279_A la_oenb_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[51\]_A la_data_out_core[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input446_A mprj_dat_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input42_A la_data_out_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__596__A _596_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output498_A _385_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output665_A _034_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1470 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1296_A wire1297/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output832_A _584_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[42\]_A la_data_out_core[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1463_A wire1463/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_3299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_2380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput90 la_data_out_mprj[62] vssd vssd vccd vccd _431_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[33\]_A la_data_out_core[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_550_ _550_/A _550_/B vssd vssd vccd vccd _550_/X sky130_fd_sc_hd__and2_4
XFILLER_35_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_481_ _609_/A _481_/B _481_/C vssd vssd vccd vccd _481_/X sky130_fd_sc_hd__and3b_4
XFILLER_44_269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input396_A mprj_adr_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[24\]_A la_data_out_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3923 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput450 mprj_dat_o_core[7] vssd vssd vccd vccd wire1283/A sky130_fd_sc_hd__buf_6
XFILLER_23_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput461 user_irq_ena[1] vssd vssd vccd vccd wire1263/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1211_A _316_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output782_A _538_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1309_A wire1309/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__492__C _492_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1580_A wire1581/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1678_A wire1679/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput902 _143_/Y vssd vssd vccd vccd mprj_dat_i_core[29] sky130_fd_sc_hd__buf_8
XFILLER_29_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput913 wire1174/X vssd vssd vccd vccd mprj_dat_o_user[0] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[15\]_A la_data_out_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput924 wire1172/X vssd vssd vccd vccd mprj_dat_o_user[1] sky130_fd_sc_hd__buf_8
Xoutput935 wire1170/X vssd vssd vccd vccd mprj_dat_o_user[2] sky130_fd_sc_hd__buf_8
XFILLER_9_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput946 wire1231/X vssd vssd vccd vccd mprj_sel_o_user[1] sky130_fd_sc_hd__buf_8
XFILLER_3_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput957 _111_/Y vssd vssd vccd vccd user_irq[0] sky130_fd_sc_hd__buf_8
XFILLER_28_2059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2642 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__204__A _204_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2643 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input144_A la_iena_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_602_ _602_/A _602_/B vssd vssd vccd vccd _602_/X sky130_fd_sc_hd__and2_4
XTAP_3533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input311_A la_oenb_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input409_A mprj_adr_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_533_ _533_/A _533_/B vssd vssd vccd vccd _533_/X sky130_fd_sc_hd__and2_4
XTAP_2843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__593__B _593_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_464_ _592_/A _464_/B _464_/C vssd vssd vccd vccd _464_/X sky130_fd_sc_hd__and3b_2
XFILLER_31_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_395_ _523_/A _395_/B _395_/C vssd vssd vccd vccd _395_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_486 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__114__A _114_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output530_A wire1090/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3731 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output628_A _001_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1161_A _344_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__487__C _487_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput280 la_oenb_mprj[118] vssd vssd vccd vccd _615_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput291 la_oenb_mprj[12] vssd vssd vccd vccd _509_/A sky130_fd_sc_hd__buf_4
XFILLER_3_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1426_A input1/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[42\] la_data_out_core[42] _205_/X vssd vssd vccd vccd _025_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_3620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput710 _075_/Y vssd vssd vccd vccd la_data_in_mprj[92] sky130_fd_sc_hd__buf_8
Xoutput721 wire1045/X vssd vssd vccd vccd la_oenb_core[101] sky130_fd_sc_hd__buf_8
Xoutput732 _608_/X vssd vssd vccd vccd la_oenb_core[111] sky130_fd_sc_hd__buf_8
Xoutput743 _618_/X vssd vssd vccd vccd la_oenb_core[121] sky130_fd_sc_hd__buf_8
XFILLER_9_3664 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput754 _513_/X vssd vssd vccd vccd la_oenb_core[16] sky130_fd_sc_hd__buf_8
Xoutput765 wire1053/X vssd vssd vccd vccd la_oenb_core[26] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[4\] la_data_out_core[4] _167_/X vssd vssd vccd vccd _151_/A
+ sky130_fd_sc_hd__nand2_2
Xoutput776 _533_/X vssd vssd vccd vccd la_oenb_core[36] sky130_fd_sc_hd__buf_8
XFILLER_5_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput787 _543_/X vssd vssd vccd vccd la_oenb_core[46] sky130_fd_sc_hd__buf_8
XFILLER_5_3539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput798 wire1050/X vssd vssd vccd vccd la_oenb_core[56] sky130_fd_sc_hd__buf_8
XFILLER_5_2816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1507 wire1507/A vssd vssd vccd vccd _263_/A sky130_fd_sc_hd__buf_6
XTAP_272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1518 wire1518/A vssd vssd vccd vccd _249_/A sky130_fd_sc_hd__buf_6
XTAP_283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1529 wire1529/A vssd vssd vccd vccd _185_/A sky130_fd_sc_hd__buf_6
XFILLER_25_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_180_ _180_/A _180_/B vssd vssd vccd vccd _180_/X sky130_fd_sc_hd__and2_1
XFILLER_10_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input261_A la_oenb_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input359_A la_oenb_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__588__B _588_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_516_ _516_/A _516_/B vssd vssd vccd vccd _516_/X sky130_fd_sc_hd__and2_4
XFILLER_37_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__109__A _109_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_447_ _575_/A _447_/B _447_/C vssd vssd vccd vccd _447_/X sky130_fd_sc_hd__and3b_4
XTAP_1983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_378_ _506_/A _378_/B _378_/C vssd vssd vccd vccd _378_/X sky130_fd_sc_hd__and3b_4
XANTENNA_wire1007_A wire1008/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output480_A _484_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output578_A wire1067/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output745_A wire1036/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__385__A_N _513_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1376_A wire1377/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1442 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output912_A wire977/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__498__B _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1543_A wire1543/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire996_A wire996/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput540 wire1081/X vssd vssd vccd vccd la_data_in_core[54] sky130_fd_sc_hd__buf_8
XFILLER_5_4037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput551 wire1072/X vssd vssd vccd vccd la_data_in_core[64] sky130_fd_sc_hd__buf_8
XFILLER_9_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput562 _443_/X vssd vssd vccd vccd la_data_in_core[74] sky130_fd_sc_hd__buf_8
Xoutput573 _453_/X vssd vssd vccd vccd la_data_in_core[84] sky130_fd_sc_hd__buf_8
XFILLER_43_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput584 wire1063/X vssd vssd vccd vccd la_data_in_core[94] sky130_fd_sc_hd__buf_8
Xoutput595 _086_/Y vssd vssd vccd vccd la_data_in_mprj[103] sky130_fd_sc_hd__buf_8
XFILLER_25_3286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1304 wire1305/X vssd vssd vccd vccd _363_/B sky130_fd_sc_hd__buf_6
Xwire1315 wire1315/A vssd vssd vccd vccd wire1315/X sky130_fd_sc_hd__buf_6
XFILLER_25_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1326 wire1327/X vssd vssd vccd vccd _353_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1337 wire1337/A vssd vssd vccd vccd wire1337/X sky130_fd_sc_hd__buf_6
XFILLER_19_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1348 wire1348/A vssd vssd vccd vccd wire1348/X sky130_fd_sc_hd__buf_6
XFILLER_5_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1359 wire1359/A vssd vssd vccd vccd wire1359/X sky130_fd_sc_hd__buf_6
XFILLER_46_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input107_A la_data_out_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_301_ _301_/A _301_/B vssd vssd vccd vccd _301_/X sky130_fd_sc_hd__and2_4
XTAP_1268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_232_ _232_/A _232_/B vssd vssd vccd vccd _232_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_163_ _163_/A vssd vssd vccd vccd _163_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_3544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input72_A la_data_out_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_094_ _094_/A vssd vssd vccd vccd _094_/Y sky130_fd_sc_hd__inv_4
XFILLER_13_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__599__A _599_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1124_A wire1125/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_160 _256_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 _468_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output695_A _062_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output862_A wire1194/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[18\] mprj_dat_i_user[18] rebuffer4/X vssd vssd vccd vccd wire1021/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA_wire1493_A wire1493/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1660_A wire1661/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3139 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__302__A _302_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[116\] la_data_out_core[116] _279_/X vssd vssd vccd vccd _099_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_28_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__400__A_N _528_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2708 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__212__A _212_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1101 _403_/X vssd vssd vccd vccd wire1101/X sky130_fd_sc_hd__buf_6
XFILLER_22_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1112 wire1113/X vssd vssd vccd vccd wire1112/X sky130_fd_sc_hd__buf_6
XFILLER_5_3199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1123 _363_/X vssd vssd vccd vccd wire1123/X sky130_fd_sc_hd__buf_6
XFILLER_19_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1134 wire1135/X vssd vssd vccd vccd wire1134/X sky130_fd_sc_hd__buf_6
XFILLER_43_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1145 _352_/X vssd vssd vccd vccd wire1145/X sky130_fd_sc_hd__buf_6
XFILLER_25_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1156 wire1157/X vssd vssd vccd vccd wire1156/X sky130_fd_sc_hd__buf_6
XANTENNA_input224_A la_iena_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1167 _341_/X vssd vssd vccd vccd wire1167/X sky130_fd_sc_hd__buf_6
Xwire1178 wire1179/X vssd vssd vccd vccd wire1178/X sky130_fd_sc_hd__buf_6
Xwire1189 _330_/X vssd vssd vccd vccd wire1189/X sky130_fd_sc_hd__buf_6
XFILLER_34_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_215_ _215_/A _215_/B vssd vssd vccd vccd _215_/X sky130_fd_sc_hd__and2_2
XFILLER_11_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_146_ _146_/A vssd vssd vccd vccd _146_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_7_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_077_ _077_/A vssd vssd vccd vccd _077_/Y sky130_fd_sc_hd__inv_4
XFILLER_45_2703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__122__A _122_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__423__A_N _551_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output610_A _100_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output708_A _073_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1339_A wire1339/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1690 wire1690/A vssd vssd vccd vccd wire1690/X sky130_fd_sc_hd__buf_6
XANTENNA__495__C _495_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1066 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1506_A wire1506/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1162 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[60\]_B _223_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__032__A _032_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput109 la_data_out_mprj[7] vssd vssd vccd vccd _376_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1578 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_698 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__207__A _207_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_60 _270_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_000_ _000_/A vssd vssd vccd vccd _000_/Y sky130_fd_sc_hd__inv_2
XANTENNA_71 _187_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_82 _169_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_93 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input174_A la_iena_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__446__A_N _574_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input341_A la_oenb_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input439_A mprj_dat_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input35_A la_data_out_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__596__B _596_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__117__A _117_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output560_A _441_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output658_A _028_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_129_ _129_/A vssd vssd vccd vccd _129_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_45_3223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1289_A wire1289/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output825_A _577_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1456_A wire1457/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[72\] la_data_out_core[72] _235_/X vssd vssd vccd vccd _055_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1623_A wire1623/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__469__A_N _597_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput80 la_data_out_mprj[53] vssd vssd vccd vccd _422_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_46_2319 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput91 la_data_out_mprj[63] vssd vssd vccd vccd _432_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_43_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1386 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_480_ _608_/A _480_/B _480_/C vssd vssd vccd vccd _480_/X sky130_fd_sc_hd__and3b_4
XFILLER_0_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input291_A la_oenb_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input389_A mprj_adr_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput440 mprj_dat_o_core[27] vssd vssd vccd vccd wire1303/A sky130_fd_sc_hd__buf_6
Xinput451 mprj_dat_o_core[8] vssd vssd vccd vccd wire1281/A sky130_fd_sc_hd__buf_6
Xinput462 user_irq_ena[2] vssd vssd vccd vccd wire1262/A sky130_fd_sc_hd__buf_6
XFILLER_40_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1204_A _321_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output775_A _532_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output942_A wire1160/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2598 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput903 wire984/X vssd vssd vccd vccd mprj_dat_i_core[2] sky130_fd_sc_hd__buf_8
XFILLER_7_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput914 wire1154/X vssd vssd vccd vccd mprj_dat_o_user[10] sky130_fd_sc_hd__buf_8
Xoutput925 wire1134/X vssd vssd vccd vccd mprj_dat_o_user[20] sky130_fd_sc_hd__buf_8
Xoutput936 wire1114/X vssd vssd vccd vccd mprj_dat_o_user[30] sky130_fd_sc_hd__buf_8
Xoutput947 wire1229/X vssd vssd vccd vccd mprj_sel_o_user[2] sky130_fd_sc_hd__buf_8
XFILLER_28_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput958 _112_/Y vssd vssd vccd vccd user_irq[1] sky130_fd_sc_hd__buf_8
XFILLER_45_3075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_4052 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3467 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__204__B _204_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__220__A _220_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input137_A la_iena_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_601_ _601_/A _601_/B vssd vssd vccd vccd _601_/X sky130_fd_sc_hd__and2_4
XTAP_3523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_532_ _532_/A _532_/B vssd vssd vccd vccd _532_/X sky130_fd_sc_hd__and2_4
XTAP_2822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input304_A la_oenb_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_463_ _591_/A _463_/B _463_/C vssd vssd vccd vccd _463_/X sky130_fd_sc_hd__and3b_2
XTAP_2877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_394_ _522_/A _394_/B _394_/C vssd vssd vccd vccd _394_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output523_A wire1096/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__130__A _130_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1154_A wire1155/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput270 la_oenb_mprj[109] vssd vssd vccd vccd _606_/A sky130_fd_sc_hd__buf_4
XFILLER_3_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput281 la_oenb_mprj[119] vssd vssd vccd vccd _616_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput292 la_oenb_mprj[13] vssd vssd vccd vccd _510_/A sky130_fd_sc_hd__buf_4
XFILLER_36_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1321_A wire1321/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output892_A wire985/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1419_A wire1420/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[35\] la_data_out_core[35] _198_/X vssd vssd vccd vccd _018_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_14_3306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__305__A _305_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput700 _066_/Y vssd vssd vccd vccd la_data_in_mprj[83] sky130_fd_sc_hd__buf_8
Xoutput711 _076_/Y vssd vssd vccd vccd la_data_in_mprj[93] sky130_fd_sc_hd__buf_8
XFILLER_9_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput722 _599_/X vssd vssd vccd vccd la_oenb_core[102] sky130_fd_sc_hd__buf_8
Xoutput733 _609_/X vssd vssd vccd vccd la_oenb_core[112] sky130_fd_sc_hd__buf_8
XFILLER_25_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput744 wire1037/X vssd vssd vccd vccd la_oenb_core[122] sky130_fd_sc_hd__buf_8
Xoutput755 _514_/X vssd vssd vccd vccd la_oenb_core[17] sky130_fd_sc_hd__buf_8
XFILLER_5_3507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3676 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput766 _524_/X vssd vssd vccd vccd la_oenb_core[27] sky130_fd_sc_hd__buf_8
Xoutput777 _534_/X vssd vssd vccd vccd la_oenb_core[37] sky130_fd_sc_hd__buf_8
XFILLER_29_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput788 _544_/X vssd vssd vccd vccd la_oenb_core[47] sky130_fd_sc_hd__buf_8
Xoutput799 _554_/X vssd vssd vccd vccd la_oenb_core[57] sky130_fd_sc_hd__buf_8
XFILLER_25_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1508 wire1508/A vssd vssd vccd vccd _262_/A sky130_fd_sc_hd__buf_6
XFILLER_42_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__040__A _040_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1519 wire1519/A vssd vssd vccd vccd _244_/A sky130_fd_sc_hd__buf_4
XFILLER_3_3253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__215__A _215_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1794 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3070 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input254_A la_iena_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input421_A mprj_dat_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_515_ _515_/A _515_/B vssd vssd vccd vccd _515_/X sky130_fd_sc_hd__and2_4
XTAP_2652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_446_ _574_/A _446_/B _446_/C vssd vssd vccd vccd _446_/X sky130_fd_sc_hd__and3b_4
XTAP_1962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_377_ _505_/A _377_/B _377_/C vssd vssd vccd vccd _377_/X sky130_fd_sc_hd__and3b_2
XFILLER_35_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output473_A _478_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__125__A _125_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmax_cap1244 wire1245/X vssd vssd vccd vccd max_cap1244/X sky130_fd_sc_hd__buf_8
XFILLER_31_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output640_A _012_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output738_A _614_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1271_A wire1272/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1369_A wire1369/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output905_A _145_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1536_A wire1536/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1703_A wire1703/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__035__A _035_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3811 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput530 wire1090/X vssd vssd vccd vccd la_data_in_core[45] sky130_fd_sc_hd__buf_8
Xoutput541 wire1080/X vssd vssd vccd vccd la_data_in_core[55] sky130_fd_sc_hd__buf_8
XFILLER_44_3855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput552 wire1071/X vssd vssd vccd vccd la_data_in_core[65] sky130_fd_sc_hd__buf_8
Xoutput563 _444_/X vssd vssd vccd vccd la_data_in_core[75] sky130_fd_sc_hd__buf_8
XFILLER_9_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput574 _454_/X vssd vssd vccd vccd la_data_in_core[85] sky130_fd_sc_hd__buf_8
Xoutput585 wire1062/X vssd vssd vccd vccd la_data_in_core[95] sky130_fd_sc_hd__buf_8
Xoutput596 _087_/Y vssd vssd vccd vccd la_data_in_mprj[104] sky130_fd_sc_hd__buf_8
XFILLER_25_3276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1305 wire1305/A vssd vssd vccd vccd wire1305/X sky130_fd_sc_hd__buf_6
XFILLER_25_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1316 wire1317/X vssd vssd vccd vccd _357_/B sky130_fd_sc_hd__buf_6
Xwire1327 wire1327/A vssd vssd vccd vccd wire1327/X sky130_fd_sc_hd__buf_6
Xwire1338 wire1339/X vssd vssd vccd vccd _347_/B sky130_fd_sc_hd__buf_6
Xwire1349 wire1350/X vssd vssd vccd vccd _312_/B sky130_fd_sc_hd__buf_6
XFILLER_41_1153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_300_ _300_/A _300_/B vssd vssd vccd vccd _300_/X sky130_fd_sc_hd__and2_4
XFILLER_42_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_231_ _231_/A _231_/B vssd vssd vccd vccd _231_/X sky130_fd_sc_hd__and2_4
XFILLER_23_582 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_162_ _162_/A vssd vssd vccd vccd _162_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_093_ _093_/A vssd vssd vccd vccd _093_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input371_A la_oenb_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input65_A la_data_out_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__599__B _599_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2052 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_150 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_161 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_172 _466_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output590_A _378_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1122 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1117_A _366_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output688_A _055_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_429_ _557_/A _429_/B _429_/C vssd vssd vccd vccd _429_/X sky130_fd_sc_hd__and3b_2
XTAP_1792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output855_A wire1204/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1486_A wire1486/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1653_A wire1654/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__302__B _302_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[0\]_A mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput1 caravel_clk vssd vssd vccd vccd input1/X sky130_fd_sc_hd__buf_6
XFILLER_4_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[109\] la_data_out_core[109] _272_/X vssd vssd vccd vccd _092_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_0_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[0\]_A la_data_out_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1102 _402_/X vssd vssd vccd vccd wire1102/X sky130_fd_sc_hd__buf_6
XFILLER_44_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1113 _368_/X vssd vssd vccd vccd wire1113/X sky130_fd_sc_hd__buf_6
XFILLER_22_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1124 wire1125/X vssd vssd vccd vccd wire1124/X sky130_fd_sc_hd__buf_6
XFILLER_19_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1135 _357_/X vssd vssd vccd vccd wire1135/X sky130_fd_sc_hd__buf_6
Xwire1146 wire1147/X vssd vssd vccd vccd wire1146/X sky130_fd_sc_hd__buf_6
XFILLER_21_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1157 _346_/X vssd vssd vccd vccd wire1157/X sky130_fd_sc_hd__buf_6
XFILLER_38_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1168 wire1169/X vssd vssd vccd vccd wire1168/X sky130_fd_sc_hd__buf_6
XFILLER_19_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1179 _335_/X vssd vssd vccd vccd wire1179/X sky130_fd_sc_hd__buf_6
XFILLER_38_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input217_A la_iena_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__375__A_N _503_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_214_ _214_/A _214_/B vssd vssd vccd vccd _214_/X sky130_fd_sc_hd__and2_2
XFILLER_15_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_145_ _145_/A vssd vssd vccd vccd _145_/Y sky130_fd_sc_hd__inv_4
XFILLER_32_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[0\] mprj_dat_i_user[0] max_cap1244/X vssd vssd vccd vccd wire1030/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_7_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_076_ _076_/A vssd vssd vccd vccd _076_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_7_3911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output603_A _093_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1680 wire1681/X vssd vssd vccd vccd _482_/B sky130_fd_sc_hd__buf_6
Xwire1691 wire1692/X vssd vssd vccd vccd _476_/B sky130_fd_sc_hd__buf_6
XFILLER_20_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1234_A _301_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1401_A wire1402/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[30\] mprj_dat_i_user[30] wire1248/X vssd vssd vccd vccd wire1000/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_33_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1586 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__313__A _313_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__398__A_N _526_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_338 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__207__B _207_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_50 _375_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_61 _270_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_72 _187_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_83 _169_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_94 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input167_A la_iena_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input334_A la_oenb_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input28_A la_data_out_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_128_ _128_/A vssd vssd vccd vccd _128_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_29_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output553_A _435_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__133__A _133_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_059_ _059_/A vssd vssd vccd vccd _059_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_wire1184_A wire1185/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output720_A wire1046/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output818_A _571_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1351_A wire1351/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1449_A wire1449/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[65\] la_data_out_core[65] _228_/X vssd vssd vccd vccd _048_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_40_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1616_A wire1616/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__308__A _308_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire971_A _129_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3422 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput70 la_data_out_mprj[44] vssd vssd vccd vccd _413_/C sky130_fd_sc_hd__clkbuf_4
Xinput81 la_data_out_mprj[54] vssd vssd vccd vccd _423_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__043__A _043_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput92 la_data_out_mprj[64] vssd vssd vccd vccd _433_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1398 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__218__A _218_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__413__A_N _541_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input284_A la_oenb_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input451_A mprj_dat_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput430 mprj_dat_o_core[18] vssd vssd vccd vccd wire1323/A sky130_fd_sc_hd__buf_6
Xinput441 mprj_dat_o_core[28] vssd vssd vccd vccd wire1301/A sky130_fd_sc_hd__buf_6
XANTENNA__400__B _400_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput452 mprj_dat_o_core[9] vssd vssd vccd vccd wire1279/A sky130_fd_sc_hd__buf_6
XFILLER_2_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__128__A _128_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output670_A _039_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output768_A _526_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1399_A wire1400/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output935_A wire1170/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput904 _144_/Y vssd vssd vccd vccd mprj_dat_i_core[30] sky130_fd_sc_hd__buf_8
Xoutput915 wire1152/X vssd vssd vccd vccd mprj_dat_o_user[11] sky130_fd_sc_hd__buf_8
Xoutput926 wire1132/X vssd vssd vccd vccd mprj_dat_o_user[21] sky130_fd_sc_hd__buf_8
Xoutput937 wire1112/X vssd vssd vccd vccd mprj_dat_o_user[31] sky130_fd_sc_hd__buf_8
XANTENNA_wire1566_A wire1567/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput948 wire1227/X vssd vssd vccd vccd mprj_sel_o_user[3] sky130_fd_sc_hd__buf_8
XFILLER_25_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput959 _113_/Y vssd vssd vccd vccd user_irq[2] sky130_fd_sc_hd__buf_8
XTAP_400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__310__B _310_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__436__A_N _564_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__038__A _038_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__501__A _501_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_600_ _600_/A _600_/B vssd vssd vccd vccd _600_/X sky130_fd_sc_hd__and2_2
XFILLER_40_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_531_ _531_/A _531_/B vssd vssd vccd vccd _531_/X sky130_fd_sc_hd__and2_4
XTAP_2812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_462_ _590_/A _462_/B _462_/C vssd vssd vccd vccd _462_/X sky130_fd_sc_hd__and3b_4
XTAP_2867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_393_ _521_/A _393_/B _393_/C vssd vssd vccd vccd _393_/X sky130_fd_sc_hd__and3b_4
XFILLER_25_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input95_A la_data_out_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output516_A wire1103/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput260 la_oenb_mprj[0] vssd vssd vccd vccd _497_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_4_3799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput271 la_oenb_mprj[10] vssd vssd vccd vccd _507_/A sky130_fd_sc_hd__buf_4
Xinput282 la_oenb_mprj[11] vssd vssd vccd vccd _508_/A sky130_fd_sc_hd__buf_4
Xinput293 la_oenb_mprj[14] vssd vssd vccd vccd _511_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__459__A_N _587_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1147_A _351_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1314_A wire1315/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output885_A wire973/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[28\] la_data_out_core[28] _191_/X vssd vssd vccd vccd _011_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_20_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__305__B _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput701 _067_/Y vssd vssd vccd vccd la_data_in_mprj[84] sky130_fd_sc_hd__buf_8
XFILLER_25_4126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput712 _077_/Y vssd vssd vccd vccd la_data_in_mprj[94] sky130_fd_sc_hd__buf_8
Xoutput723 wire1044/X vssd vssd vccd vccd la_oenb_core[103] sky130_fd_sc_hd__buf_8
Xoutput734 _610_/X vssd vssd vccd vccd la_oenb_core[113] sky130_fd_sc_hd__buf_8
XFILLER_29_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput745 wire1036/X vssd vssd vccd vccd la_oenb_core[123] sky130_fd_sc_hd__buf_8
Xoutput756 _515_/X vssd vssd vccd vccd la_oenb_core[18] sky130_fd_sc_hd__buf_8
Xoutput767 _525_/X vssd vssd vccd vccd la_oenb_core[28] sky130_fd_sc_hd__buf_8
XFILLER_9_3688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput778 _535_/X vssd vssd vccd vccd la_oenb_core[38] sky130_fd_sc_hd__buf_8
XFILLER_7_4091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput789 _545_/X vssd vssd vccd vccd la_oenb_core[48] sky130_fd_sc_hd__buf_8
XANTENNA_powergood_check_mprj2_vdd_logic1 output954/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1509 wire1509/A vssd vssd vccd vccd _261_/A sky130_fd_sc_hd__buf_6
XTAP_274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__215__B _215_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__231__A _231_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input247_A la_iena_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input414_A mprj_adr_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input10_A la_data_out_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_514_ _514_/A _514_/B vssd vssd vccd vccd _514_/X sky130_fd_sc_hd__and2_4
XFILLER_33_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_445_ _573_/A _445_/B _445_/C vssd vssd vccd vccd _445_/X sky130_fd_sc_hd__and3b_4
XTAP_1963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4074 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_376_ _504_/A _376_/B _376_/C vssd vssd vccd vccd _376_/X sky130_fd_sc_hd__and3b_4
XFILLER_9_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output466_A wire1058/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output633_A _005_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__141__A _141_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output800_A wire1049/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1104 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1431_A wire1431/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1529_A wire1529/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__316__A _316_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[90\]_A la_data_out_core[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput520 wire1099/X vssd vssd vccd vccd la_data_in_core[36] sky130_fd_sc_hd__buf_8
Xoutput531 wire1089/X vssd vssd vccd vccd la_data_in_core[46] sky130_fd_sc_hd__buf_8
Xoutput542 wire1079/X vssd vssd vccd vccd la_data_in_core[56] sky130_fd_sc_hd__buf_8
XFILLER_5_4039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput553 _435_/X vssd vssd vccd vccd la_data_in_core[66] sky130_fd_sc_hd__buf_8
XFILLER_43_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput564 _445_/X vssd vssd vccd vccd la_data_in_core[76] sky130_fd_sc_hd__buf_8
Xoutput575 _455_/X vssd vssd vccd vccd la_data_in_core[86] sky130_fd_sc_hd__buf_8
XANTENNA__051__A _051_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput586 _465_/X vssd vssd vccd vccd la_data_in_core[96] sky130_fd_sc_hd__buf_8
XFILLER_8_1004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput597 _088_/Y vssd vssd vccd vccd la_data_in_mprj[105] sky130_fd_sc_hd__buf_8
Xwire1306 wire1307/X vssd vssd vccd vccd _362_/B sky130_fd_sc_hd__buf_6
XANTENNA_input2_A caravel_clk2 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1317 wire1317/A vssd vssd vccd vccd wire1317/X sky130_fd_sc_hd__buf_6
XFILLER_3_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1328 wire1329/X vssd vssd vccd vccd _352_/B sky130_fd_sc_hd__buf_6
XFILLER_25_1853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1339 wire1339/A vssd vssd vccd vccd wire1339/X sky130_fd_sc_hd__buf_6
XFILLER_21_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_230_ _230_/A _230_/B vssd vssd vccd vccd _230_/X sky130_fd_sc_hd__and2_4
XFILLER_23_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_594 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__226__A _226_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_161_ _161_/A vssd vssd vccd vccd _161_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input197_A la_iena_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_092_ _092_/A vssd vssd vccd vccd _092_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_3579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[81\]_A la_data_out_core[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input364_A la_oenb_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input58_A la_data_out_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_3736 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3560 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _213_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_173 _466_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_428_ _556_/A _428_/B _428_/C vssd vssd vccd vccd _428_/X sky130_fd_sc_hd__and3b_2
XTAP_1793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1012_A wire1013/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output583_A _462_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__136__A _136_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_359_ _359_/A _359_/B vssd vssd vccd vccd _359_/X sky130_fd_sc_hd__and2_4
XFILLER_13_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output750_A _509_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[72\]_A la_data_out_core[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output848_A wire1226/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1381_A wire1381/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_782 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1479_A wire1480/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[95\] la_data_out_core[95] wire1260/X vssd vssd vccd vccd _078_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_6_2902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput2 caravel_clk2 vssd vssd vccd vccd input2/X sky130_fd_sc_hd__buf_6
XFILLER_42_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[0\]_B _625_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__046__A _046_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[63\]_A la_data_out_core[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1103 _401_/X vssd vssd vccd vccd wire1103/X sky130_fd_sc_hd__buf_6
XFILLER_21_2204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1114 wire1115/X vssd vssd vccd vccd wire1114/X sky130_fd_sc_hd__buf_6
Xwire1125 _362_/X vssd vssd vccd vccd wire1125/X sky130_fd_sc_hd__buf_6
XFILLER_22_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1136 wire1137/X vssd vssd vccd vccd wire1136/X sky130_fd_sc_hd__buf_6
XFILLER_21_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1147 _351_/X vssd vssd vccd vccd wire1147/X sky130_fd_sc_hd__buf_6
Xwire1158 wire1159/X vssd vssd vccd vccd wire1158/X sky130_fd_sc_hd__buf_6
XFILLER_21_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1169 _340_/X vssd vssd vccd vccd wire1169/X sky130_fd_sc_hd__buf_6
XFILLER_38_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input112_A la_data_out_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_213_ _213_/A _213_/B vssd vssd vccd vccd _213_/X sky130_fd_sc_hd__and2_2
XFILLER_32_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_144_ _144_/A vssd vssd vccd vccd _144_/Y sky130_fd_sc_hd__inv_4
XFILLER_10_2620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[54\]_A la_data_out_core[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_075_ _075_/A vssd vssd vccd vccd _075_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__403__B _403_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1670 wire1671/X vssd vssd vccd vccd _487_/B sky130_fd_sc_hd__buf_6
XFILLER_20_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1681 wire1681/A vssd vssd vccd vccd wire1681/X sky130_fd_sc_hd__buf_6
XFILLER_1_2865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1692 wire1692/A vssd vssd vccd vccd wire1692/X sky130_fd_sc_hd__buf_6
XFILLER_18_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1227_A wire1228/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output798_A wire1050/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_split13_A split13/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[10\] la_data_out_core[10] _173_/X vssd vssd vccd vccd _157_/A
+ sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_gates\[23\] mprj_dat_i_user[23] split13/X vssd vssd vccd vccd wire1013/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_37_1598 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1596_A wire1596/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[45\]_A la_data_out_core[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__313__B _313_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[121\] la_data_out_core[121] _284_/X vssd vssd vccd vccd _104_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_6_2776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_40 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_51 _375_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_62 _270_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_73 _187_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_84 _169_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[36\]_A la_data_out_core[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_95 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__504__A _504_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[120\]_A la_data_out_core[120] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_14_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1912 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input327_A la_oenb_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__492__A_N _620_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[27\]_A la_data_out_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[111\]_A la_data_out_core[111] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
X_127_ _127_/A vssd vssd vccd vccd _127_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_10_3195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_058_ _058_/A vssd vssd vccd vccd _058_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_output546_A _374_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1177_A _336_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output713_A _078_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1344_A wire1345/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[58\] la_data_out_core[58] _221_/X vssd vssd vccd vccd _041_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_1_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1609_A wire1609/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3338 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__308__B _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2394 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[18\]_A la_data_out_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__324__A _324_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_A la_data_out_core[102] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xinput60 la_data_out_mprj[35] vssd vssd vccd vccd _404_/C sky130_fd_sc_hd__clkbuf_4
Xinput71 la_data_out_mprj[45] vssd vssd vccd vccd _414_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput82 la_data_out_mprj[55] vssd vssd vccd vccd _424_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput93 la_data_out_mprj[65] vssd vssd vccd vccd _434_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_2711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__234__A _234_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input277_A la_oenb_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input444_A mprj_dat_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input40_A la_data_out_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput420 mprj_cyc_o_core vssd vssd vccd vccd wire1343/A sky130_fd_sc_hd__buf_6
Xinput431 mprj_dat_o_core[19] vssd vssd vccd vccd wire1321/A sky130_fd_sc_hd__buf_6
XFILLER_40_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput442 mprj_dat_o_core[29] vssd vssd vccd vccd wire1299/A sky130_fd_sc_hd__buf_6
XANTENNA__400__C _400_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput453 mprj_iena_wb vssd vssd vccd vccd wire1277/A sky130_fd_sc_hd__buf_8
XFILLER_27_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_486 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3202 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output496_A _383_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__144__A _144_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__388__A_N _516_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1294_A wire1295/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput905 _145_/Y vssd vssd vccd vccd mprj_dat_i_core[31] sky130_fd_sc_hd__buf_8
XFILLER_45_3022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput916 wire1150/X vssd vssd vccd vccd mprj_dat_o_user[12] sky130_fd_sc_hd__buf_8
XFILLER_29_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2018 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output830_A _582_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput927 wire1130/X vssd vssd vccd vccd mprj_dat_o_user[22] sky130_fd_sc_hd__buf_8
XFILLER_10_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput938 wire1168/X vssd vssd vccd vccd mprj_dat_o_user[3] sky130_fd_sc_hd__buf_8
XFILLER_45_3055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output928_A wire1128/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput949 wire1237/X vssd vssd vccd vccd mprj_stb_o_user sky130_fd_sc_hd__buf_8
XFILLER_23_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1461_A wire1461/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1559_A wire1559/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__319__A _319_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__054__A _054_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__501__B _501_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1450 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_530_ _530_/A _530_/B vssd vssd vccd vccd _530_/X sky130_fd_sc_hd__and2_4
XTAP_3558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_461_ _589_/A _461_/B _461_/C vssd vssd vccd vccd _461_/X sky130_fd_sc_hd__and3b_2
XFILLER_32_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_392_ _520_/A _392_/B _392_/C vssd vssd vccd vccd _392_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input394_A mprj_adr_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input88_A la_data_out_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3290 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__411__B _411_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput250 la_iena_mprj[91] vssd vssd vccd vccd _254_/B sky130_fd_sc_hd__clkbuf_4
Xinput261 la_oenb_mprj[100] vssd vssd vccd vccd _597_/A sky130_fd_sc_hd__clkbuf_4
Xinput272 la_oenb_mprj[110] vssd vssd vccd vccd _607_/A sky130_fd_sc_hd__clkbuf_4
Xinput283 la_oenb_mprj[120] vssd vssd vccd vccd _617_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_output509_A wire1109/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput294 la_oenb_mprj[15] vssd vssd vccd vccd _512_/A sky130_fd_sc_hd__buf_4
XFILLER_18_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__139__A _139_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output780_A _500_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output878_A wire1217/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1676_A wire1677/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput702 _068_/Y vssd vssd vccd vccd la_data_in_mprj[85] sky130_fd_sc_hd__buf_8
Xoutput713 _078_/Y vssd vssd vccd vccd la_data_in_mprj[95] sky130_fd_sc_hd__buf_8
Xoutput724 _601_/X vssd vssd vccd vccd la_oenb_core[104] sky130_fd_sc_hd__buf_8
Xoutput735 wire1041/X vssd vssd vccd vccd la_oenb_core[114] sky130_fd_sc_hd__buf_8
XANTENNA__602__A _602_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput746 wire1035/X vssd vssd vccd vccd la_oenb_core[124] sky130_fd_sc_hd__buf_8
Xoutput757 _516_/X vssd vssd vccd vccd la_oenb_core[19] sky130_fd_sc_hd__buf_8
Xoutput768 _526_/X vssd vssd vccd vccd la_oenb_core[29] sky130_fd_sc_hd__buf_8
Xoutput779 _536_/X vssd vssd vccd vccd la_oenb_core[39] sky130_fd_sc_hd__buf_8
XANTENNA__321__B _321_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__403__A_N _531_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__049__A _049_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__512__A _512_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__231__B _231_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input142_A la_iena_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input407_A mprj_adr_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_513_ _513_/A _513_/B vssd vssd vccd vccd _513_/X sky130_fd_sc_hd__and2_4
XTAP_2632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_444_ _572_/A _444_/B _444_/C vssd vssd vccd vccd _444_/X sky130_fd_sc_hd__and3b_4
XTAP_2687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_375_ _503_/A _375_/B _375_/C vssd vssd vccd vccd _375_/X sky130_fd_sc_hd__and3b_1
XTAP_1997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__406__B _406_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmax_cap1246 split13/A vssd vssd vccd vccd wire1245/A sky130_fd_sc_hd__buf_8
XFILLER_13_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__426__A_N _554_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output626_A _163_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_802 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2070 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[40\] la_data_out_core[40] _203_/X vssd vssd vccd vccd _023_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_3230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__316__B _316_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[90\]_B _253_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput510 wire1108/X vssd vssd vccd vccd la_data_in_core[27] sky130_fd_sc_hd__buf_8
XFILLER_5_4007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__332__A _332_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput521 wire1098/X vssd vssd vccd vccd la_data_in_core[37] sky130_fd_sc_hd__buf_8
XFILLER_44_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput532 wire1088/X vssd vssd vccd vccd la_data_in_core[47] sky130_fd_sc_hd__buf_8
Xoutput543 wire1078/X vssd vssd vccd vccd la_data_in_core[57] sky130_fd_sc_hd__buf_8
Xoutput554 _436_/X vssd vssd vccd vccd la_data_in_core[67] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[2\] la_data_out_core[2] _165_/X vssd vssd vccd vccd _149_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_44_3879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput565 _446_/X vssd vssd vccd vccd la_data_in_core[77] sky130_fd_sc_hd__buf_8
Xoutput576 _456_/X vssd vssd vccd vccd la_data_in_core[87] sky130_fd_sc_hd__buf_8
Xoutput587 wire1061/X vssd vssd vccd vccd la_data_in_core[97] sky130_fd_sc_hd__buf_8
Xoutput598 _089_/Y vssd vssd vccd vccd la_data_in_mprj[106] sky130_fd_sc_hd__buf_8
XFILLER_8_1016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1307 wire1307/A vssd vssd vccd vccd wire1307/X sky130_fd_sc_hd__buf_6
XFILLER_25_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1318 wire1319/X vssd vssd vccd vccd _338_/B sky130_fd_sc_hd__buf_6
Xwire1329 wire1329/A vssd vssd vccd vccd wire1329/X sky130_fd_sc_hd__buf_6
XFILLER_3_3063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__507__A _507_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__226__B _226_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_160_ _160_/A vssd vssd vccd vccd _160_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_091_ _091_/A vssd vssd vccd vccd _091_/Y sky130_fd_sc_hd__inv_4
XFILLER_10_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[81\]_B _244_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__449__A_N _577_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__242__A _242_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input357_A la_oenb_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_130 _197_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 _213_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_152 _329_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_163 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _466_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_427_ _555_/A _427_/B _427_/C vssd vssd vccd vccd _427_/X sky130_fd_sc_hd__and3b_4
XTAP_1772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_358_ _358_/A _358_/B vssd vssd vccd vccd _358_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1005_A wire1006/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output576_A _456_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_289_ _289_/A _289_/B vssd vssd vccd vccd _289_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[72\]_B _235_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output743_A _618_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_794 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1374_A wire1375/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output910_A wire979/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[88\] la_data_out_core[88] _251_/X vssd vssd vccd vccd _071_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_9_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1541_A wire1541/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1639_A wire1639/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput3 caravel_rstn vssd vssd vccd vccd input3/X sky130_fd_sc_hd__buf_6
XFILLER_20_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire994_A wire994/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__327__A _327_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[63\]_B _226_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__062__A _062_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3643 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1104 _400_/X vssd vssd vccd vccd wire1104/X sky130_fd_sc_hd__buf_6
XFILLER_44_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1115 _367_/X vssd vssd vccd vccd wire1115/X sky130_fd_sc_hd__buf_6
XFILLER_25_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1126 wire1127/X vssd vssd vccd vccd wire1126/X sky130_fd_sc_hd__buf_6
XFILLER_38_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1137 _356_/X vssd vssd vccd vccd wire1137/X sky130_fd_sc_hd__buf_6
XFILLER_22_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1148 wire1149/X vssd vssd vccd vccd wire1148/X sky130_fd_sc_hd__buf_6
Xwire1159 _345_/X vssd vssd vccd vccd wire1159/X sky130_fd_sc_hd__buf_6
XFILLER_28_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input105_A la_data_out_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__237__A _237_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_212_ _212_/A _212_/B vssd vssd vccd vccd _212_/X sky130_fd_sc_hd__and2_2
X_143_ _143_/A vssd vssd vccd vccd _143_/Y sky130_fd_sc_hd__inv_4
XFILLER_13_1032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[54\]_B _217_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input70_A la_data_out_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_074_ _074_/A vssd vssd vccd vccd _074_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_13_1087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_3523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1660 wire1661/X vssd vssd vccd vccd _492_/B sky130_fd_sc_hd__buf_6
Xwire1671 wire1671/A vssd vssd vccd vccd wire1671/X sky130_fd_sc_hd__buf_6
XFILLER_1_3589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1682 wire1683/X vssd vssd vccd vccd _481_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1693 wire1693/A vssd vssd vccd vccd _475_/B sky130_fd_sc_hd__buf_6
XFILLER_18_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1122_A wire1123/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output693_A _060_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output860_A wire1197/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[16\] mprj_dat_i_user[16] rebuffer3/X vssd vssd vccd vccd wire1023/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_31_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1491_A wire1491/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1589_A wire1589/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire990 _082_/Y vssd vssd vccd vccd wire990/X sky130_fd_sc_hd__buf_6
XFILLER_28_2904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_3215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__610__A _610_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[114\] la_data_out_core[114] _277_/X vssd vssd vccd vccd _097_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_2_1907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__057__A _057_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_30 _202_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_41 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_52 _375_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_63 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3664 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_74 _187_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_85 _169_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[36\]_B _199_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_96 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__504__B _504_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[120\]_B _283_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3104 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__520__A _520_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input222_A la_iena_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_126_ _126_/A vssd vssd vccd vccd _126_/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__414__B _414_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[111\]_B _274_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_057_ _057_/A vssd vssd vccd vccd _057_/Y sky130_fd_sc_hd__clkinv_4
XTAP_605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3743 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output539_A wire1082/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output706_A _072_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1337_A wire1337/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1490 wire1490/A vssd vssd vccd vccd _280_/A sky130_fd_sc_hd__buf_6
XFILLER_19_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1504_A wire1504/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[20\]_A mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__605__A _605_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[18\]_B _181_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__324__B _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_B wire1255/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput50 la_data_out_mprj[26] vssd vssd vccd vccd _395_/C sky130_fd_sc_hd__clkbuf_4
Xinput61 la_data_out_mprj[36] vssd vssd vccd vccd _405_/C sky130_fd_sc_hd__clkbuf_4
Xinput72 la_data_out_mprj[46] vssd vssd vccd vccd _415_/C sky130_fd_sc_hd__clkbuf_4
Xinput83 la_data_out_mprj[56] vssd vssd vccd vccd _425_/C sky130_fd_sc_hd__clkbuf_4
Xinput94 la_data_out_mprj[66] vssd vssd vccd vccd _435_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__340__A _340_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_782 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[11\]_A mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__515__A _515_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3450 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__234__B _234_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input172_A la_iena_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__250__A _250_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input437_A mprj_dat_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput410 mprj_adr_o_core[2] vssd vssd vccd vccd wire1369/A sky130_fd_sc_hd__buf_6
Xinput421 mprj_dat_o_core[0] vssd vssd vccd vccd wire1341/A sky130_fd_sc_hd__buf_6
XANTENNA_input33_A la_data_out_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput432 mprj_dat_o_core[1] vssd vssd vccd vccd wire1319/A sky130_fd_sc_hd__buf_6
XFILLER_0_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput443 mprj_dat_o_core[2] vssd vssd vccd vccd wire1297/A sky130_fd_sc_hd__buf_6
XFILLER_40_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput454 mprj_sel_o_core[0] vssd vssd vccd vccd wire1276/A sky130_fd_sc_hd__buf_6
XFILLER_44_1890 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__409__B _409_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_498 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output489_A _492_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_109_ _109_/A vssd vssd vccd vccd _109_/Y sky130_fd_sc_hd__inv_2
Xoutput906 wire983/X vssd vssd vccd vccd mprj_dat_i_core[3] sky130_fd_sc_hd__buf_8
Xoutput917 wire1148/X vssd vssd vccd vccd mprj_dat_o_user[13] sky130_fd_sc_hd__buf_8
Xoutput928 wire1128/X vssd vssd vccd vccd mprj_dat_o_user[23] sky130_fd_sc_hd__buf_8
XFILLER_23_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1287_A wire1287/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput939 wire1166/X vssd vssd vccd vccd mprj_dat_o_user[4] sky130_fd_sc_hd__buf_8
XFILLER_45_3067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output823_A _576_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__160__A _160_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1454_A wire1455/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2850 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[70\] la_data_out_core[70] _233_/X vssd vssd vccd vccd _053_/A
+ sky130_fd_sc_hd__nand2_8
XTAP_468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1064 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1719_A wire1719/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__319__B _319_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__335__A _335_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__482__A_N _610_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__070__A _070_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1462 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_460_ _588_/A _460_/B _460_/C vssd vssd vccd vccd _460_/X sky130_fd_sc_hd__and3b_2
XTAP_2847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_391_ _519_/A _391_/B _391_/C vssd vssd vccd vccd _391_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__245__A _245_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input387_A la_oenb_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput240 la_iena_mprj[82] vssd vssd vccd vccd _245_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput251 la_iena_mprj[92] vssd vssd vccd vccd _255_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput262 la_oenb_mprj[101] vssd vssd vccd vccd _598_/A sky130_fd_sc_hd__buf_4
XFILLER_2_3470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput273 la_oenb_mprj[111] vssd vssd vccd vccd _608_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput284 la_oenb_mprj[121] vssd vssd vccd vccd _618_/A sky130_fd_sc_hd__clkbuf_4
Xinput295 la_oenb_mprj[16] vssd vssd vccd vccd _513_/A sky130_fd_sc_hd__buf_4
XFILLER_18_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_589_ _589_/A _589_/B vssd vssd vccd vccd _589_/X sky130_fd_sc_hd__and2_4
XFILLER_38_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1202_A wire1203/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output773_A _530_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output940_A wire1164/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput703 _069_/Y vssd vssd vccd vccd la_data_in_mprj[86] sky130_fd_sc_hd__buf_8
XANTENNA_wire1571_A wire1571/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput714 _079_/Y vssd vssd vccd vccd la_data_in_mprj[96] sky130_fd_sc_hd__buf_8
XANTENNA_wire1669_A wire1669/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput725 _602_/X vssd vssd vccd vccd la_oenb_core[105] sky130_fd_sc_hd__buf_8
Xoutput736 _612_/X vssd vssd vccd vccd la_oenb_core[115] sky130_fd_sc_hd__buf_8
XANTENNA__602__B _602_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput747 wire1034/X vssd vssd vccd vccd la_oenb_core[125] sky130_fd_sc_hd__buf_8
Xoutput758 _498_/X vssd vssd vccd vccd la_oenb_core[1] sky130_fd_sc_hd__buf_8
Xoutput769 _499_/X vssd vssd vccd vccd la_oenb_core[2] sky130_fd_sc_hd__buf_8
XTAP_210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__065__A _065_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__512__B _512_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input135_A la_iena_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__378__A_N _506_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_512_ _512_/A _512_/B vssd vssd vccd vccd _512_/X sky130_fd_sc_hd__and2_4
XTAP_2622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input302_A la_oenb_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_443_ _571_/A _443_/B _443_/C vssd vssd vccd vccd _443_/X sky130_fd_sc_hd__and3b_4
XTAP_1943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_374_ _502_/A _374_/B _374_/C vssd vssd vccd vccd _374_/X sky130_fd_sc_hd__and3b_4
XTAP_1987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmax_cap1247 wire1248/X vssd vssd vccd vccd split13/A sky130_fd_sc_hd__buf_8
XFILLER_29_2114 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output521_A wire1098/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output619_A _108_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1152_A wire1153/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1417_A wire1417/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output890_A wire968/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[33\] la_data_out_core[33] _196_/X vssd vssd vccd vccd _016_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_2552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__613__A _613_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput500 _387_/X vssd vssd vccd vccd la_data_in_core[18] sky130_fd_sc_hd__buf_8
Xoutput511 wire1107/X vssd vssd vccd vccd la_data_in_core[28] sky130_fd_sc_hd__buf_8
XFILLER_9_3432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput522 wire1097/X vssd vssd vccd vccd la_data_in_core[38] sky130_fd_sc_hd__buf_8
XFILLER_5_4019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__332__B _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput533 wire1087/X vssd vssd vccd vccd la_data_in_core[48] sky130_fd_sc_hd__buf_8
Xoutput544 wire1077/X vssd vssd vccd vccd la_data_in_core[58] sky130_fd_sc_hd__buf_8
Xoutput555 wire1070/X vssd vssd vccd vccd la_data_in_core[68] sky130_fd_sc_hd__buf_8
Xoutput566 _447_/X vssd vssd vccd vccd la_data_in_core[78] sky130_fd_sc_hd__buf_8
XANTENNA_user_wb_dat_gates\[3\]_A mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput577 _457_/X vssd vssd vccd vccd la_data_in_core[88] sky130_fd_sc_hd__buf_8
XFILLER_29_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput588 wire1060/X vssd vssd vccd vccd la_data_in_core[98] sky130_fd_sc_hd__buf_8
Xoutput599 _090_/Y vssd vssd vccd vccd la_data_in_mprj[107] sky130_fd_sc_hd__buf_8
XFILLER_25_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1308 wire1309/X vssd vssd vccd vccd _361_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1319 wire1319/A vssd vssd vccd vccd wire1319/X sky130_fd_sc_hd__buf_6
XFILLER_3_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[3\]_A la_data_out_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__507__B _507_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_090_ _090_/A vssd vssd vccd vccd _090_/Y sky130_fd_sc_hd__inv_4
XFILLER_13_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__523__A _523_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__242__B _242_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input252_A la_iena_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_120 mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _197_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_142 _607_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_153 _329_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_164 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_426_ _554_/A _426_/B _426_/C vssd vssd vccd vccd _426_/X sky130_fd_sc_hd__and3b_4
XTAP_1762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__417__B _417_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_357_ _357_/A _357_/B vssd vssd vccd vccd _357_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_288_ _288_/A _288_/B vssd vssd vccd vccd _288_/X sky130_fd_sc_hd__and2_4
XANTENNA_output471_A _476_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output569_A _449_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output736_A _612_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1367_A wire1368/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output903_A wire984/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1534_A wire1534/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput4 la_data_out_mprj[0] vssd vssd vccd vccd _369_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_20_3176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1701_A wire1701/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__608__A _608_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__327__B _327_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__343__A _343_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3699 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1105 _399_/X vssd vssd vccd vccd wire1105/X sky130_fd_sc_hd__buf_6
Xwire1116 wire1117/X vssd vssd vccd vccd wire1116/X sky130_fd_sc_hd__buf_6
XFILLER_40_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1127 _361_/X vssd vssd vccd vccd wire1127/X sky130_fd_sc_hd__buf_6
XFILLER_25_2397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1138 wire1139/X vssd vssd vccd vccd wire1138/X sky130_fd_sc_hd__buf_6
Xwire1149 _350_/X vssd vssd vccd vccd wire1149/X sky130_fd_sc_hd__buf_6
XFILLER_21_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__518__A _518_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__237__B _237_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__416__A_N _544_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_211_ _211_/A _211_/B vssd vssd vccd vccd _211_/X sky130_fd_sc_hd__and2_2
XFILLER_36_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_142_ _142_/A vssd vssd vccd vccd _142_/Y sky130_fd_sc_hd__inv_4
XFILLER_32_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__253__A _253_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_073_ _073_/A vssd vssd vccd vccd _073_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_30_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input63_A la_data_out_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3671 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1650 wire1650/A vssd vssd vccd vccd _497_/B sky130_fd_sc_hd__buf_6
Xwire1661 wire1661/A vssd vssd vccd vccd wire1661/X sky130_fd_sc_hd__buf_6
XFILLER_24_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1672 wire1673/X vssd vssd vccd vccd _486_/B sky130_fd_sc_hd__buf_6
XFILLER_18_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1683 wire1683/A vssd vssd vccd vccd wire1683/X sky130_fd_sc_hd__buf_6
Xwire1694 wire1695/X vssd vssd vccd vccd _474_/B sky130_fd_sc_hd__buf_6
XFILLER_20_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1115_A _367_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output686_A _053_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_409_ _537_/A _409_/B _409_/C vssd vssd vccd vccd _409_/X sky130_fd_sc_hd__and3b_2
XFILLER_32_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output853_A wire1206/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire980 _120_/Y vssd vssd vccd vccd wire980/X sky130_fd_sc_hd__buf_6
XANTENNA_wire1484_A wire1485/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire991 _054_/Y vssd vssd vccd vccd wire991/X sky130_fd_sc_hd__buf_6
XFILLER_6_4103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1651_A wire1652/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__610__B _610_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_942 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[107\] la_data_out_core[107] wire1250/X vssd vssd vccd vccd
+ _090_/A sky130_fd_sc_hd__nand2_4
XANTENNA__439__A_N _567_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__338__A _338_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_330 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_20 _196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_31 _214_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_42 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_53 _375_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_64 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_75 _187_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3676 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__073__A _073_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_86 _168_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_97 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3463 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__520__B _520_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2150 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input215_A la_iena_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__248__A _248_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_125_ _125_/A vssd vssd vccd vccd _125_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_10_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_056_ _056_/A vssd vssd vccd vccd _056_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__430__B _430_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output601_A _092_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1480 wire1480/A vssd vssd vccd vccd wire1480/X sky130_fd_sc_hd__buf_6
XFILLER_1_3398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1491 wire1491/A vssd vssd vccd vccd _279_/A sky130_fd_sc_hd__buf_6
XFILLER_21_2581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1232_A _302_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__158__A _158_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[20\]_B split13/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1699_A wire1699/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__605__B _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput40 la_data_out_mprj[17] vssd vssd vccd vccd _386_/C sky130_fd_sc_hd__clkbuf_4
Xinput51 la_data_out_mprj[27] vssd vssd vccd vccd _396_/C sky130_fd_sc_hd__clkbuf_4
Xinput62 la_data_out_mprj[37] vssd vssd vccd vccd _406_/C sky130_fd_sc_hd__clkbuf_4
Xinput73 la_data_out_mprj[47] vssd vssd vccd vccd _416_/C sky130_fd_sc_hd__clkbuf_4
Xinput84 la_data_out_mprj[57] vssd vssd vccd vccd _426_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_7_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput95 la_data_out_mprj[67] vssd vssd vccd vccd _436_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__621__A _621_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__340__B _340_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2058 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2470 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3298 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_912 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_794 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__068__A _068_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__515__B _515_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__531__A _531_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input165_A la_iena_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__250__B _250_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput400 mprj_adr_o_core[20] vssd vssd vccd vccd wire1390/A sky130_fd_sc_hd__buf_6
XFILLER_27_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput411 mprj_adr_o_core[30] vssd vssd vccd vccd wire1366/A sky130_fd_sc_hd__buf_6
XFILLER_24_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput422 mprj_dat_o_core[10] vssd vssd vccd vccd wire1339/A sky130_fd_sc_hd__buf_6
Xinput433 mprj_dat_o_core[20] vssd vssd vccd vccd wire1317/A sky130_fd_sc_hd__buf_6
XANTENNA_input332_A la_oenb_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput444 mprj_dat_o_core[30] vssd vssd vccd vccd wire1295/A sky130_fd_sc_hd__buf_6
Xinput455 mprj_sel_o_core[1] vssd vssd vccd vccd wire1274/A sky130_fd_sc_hd__buf_6
XFILLER_0_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input26_A la_data_out_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_108_ _108_/A vssd vssd vccd vccd _108_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput907 wire982/X vssd vssd vccd vccd mprj_dat_i_core[4] sky130_fd_sc_hd__buf_8
XANTENNA_output551_A wire1072/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput918 wire1146/X vssd vssd vccd vccd mprj_dat_o_user[14] sky130_fd_sc_hd__buf_8
XFILLER_25_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput929 wire1126/X vssd vssd vccd vccd mprj_dat_o_user[24] sky130_fd_sc_hd__buf_8
XANTENNA_output649_A _020_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_039_ _039_/A vssd vssd vccd vccd _039_/Y sky130_fd_sc_hd__inv_2
XANTENNA_wire1182_A wire1183/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output816_A _569_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1076 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[63\] la_data_out_core[63] _226_/X vssd vssd vccd vccd _046_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_23_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__616__A _616_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__335__B _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_390_ _518_/A _390_/B _390_/C vssd vssd vccd vccd _390_/X sky130_fd_sc_hd__and3b_4
XFILLER_0_1270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__526__A _526_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__245__B _245_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input282_A la_oenb_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__261__A _261_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput230 la_iena_mprj[73] vssd vssd vccd vccd _236_/B sky130_fd_sc_hd__clkbuf_4
Xinput241 la_iena_mprj[83] vssd vssd vccd vccd _246_/B sky130_fd_sc_hd__clkbuf_4
Xinput252 la_iena_mprj[93] vssd vssd vccd vccd _256_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3460 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput263 la_oenb_mprj[102] vssd vssd vccd vccd _599_/A sky130_fd_sc_hd__clkbuf_4
Xinput274 la_oenb_mprj[112] vssd vssd vccd vccd _609_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput285 la_oenb_mprj[122] vssd vssd vccd vccd _619_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput296 la_oenb_mprj[17] vssd vssd vccd vccd _514_/A sky130_fd_sc_hd__buf_4
XFILLER_18_3424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3468 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_588_ _588_/A _588_/B vssd vssd vccd vccd _588_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1028_A wire1028/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output599_A _090_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output766_A _524_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1397_A wire1398/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output933_A wire1118/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput704 _070_/Y vssd vssd vccd vccd la_data_in_mprj[87] sky130_fd_sc_hd__buf_8
XFILLER_29_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput715 _080_/Y vssd vssd vccd vccd la_data_in_mprj[97] sky130_fd_sc_hd__buf_8
XANTENNA__171__A _171_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput726 _603_/X vssd vssd vccd vccd la_oenb_core[106] sky130_fd_sc_hd__buf_8
XFILLER_25_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput737 wire1040/X vssd vssd vccd vccd la_oenb_core[116] sky130_fd_sc_hd__buf_8
XANTENNA_wire1564_A wire1565/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput748 wire1033/X vssd vssd vccd vccd la_oenb_core[126] sky130_fd_sc_hd__buf_8
XFILLER_28_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput759 _517_/X vssd vssd vccd vccd la_oenb_core[20] sky130_fd_sc_hd__buf_8
XTAP_200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1731_A wire1732/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[93\]_A la_data_out_core[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3030 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input128_A la_data_out_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_511_ _511_/A _511_/B vssd vssd vccd vccd _511_/X sky130_fd_sc_hd__and2_4
XTAP_3368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_442_ _570_/A _442_/B _442_/C vssd vssd vccd vccd _442_/X sky130_fd_sc_hd__and3b_4
XTAP_1933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__256__A _256_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_373_ _501_/A _373_/B _373_/C vssd vssd vccd vccd _373_/X sky130_fd_sc_hd__and3b_4
XTAP_1988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input93_A la_data_out_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_A la_data_out_core[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[9\] mprj_dat_i_user[9] rebuffer2/X vssd vssd vccd vccd wire992/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_6_955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2832 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output514_A wire1105/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1145_A _352_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1312_A wire1313/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output883_A wire975/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__472__A_N _600_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__166__A _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3298 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[26\] la_data_out_core[26] _189_/X vssd vssd vccd vccd _009_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_36_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[75\]_A la_data_out_core[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__613__B _613_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput501 _388_/X vssd vssd vccd vccd la_data_in_core[19] sky130_fd_sc_hd__buf_8
Xoutput512 wire1106/X vssd vssd vccd vccd la_data_in_core[29] sky130_fd_sc_hd__buf_8
XFILLER_29_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput523 wire1096/X vssd vssd vccd vccd la_data_in_core[39] sky130_fd_sc_hd__buf_8
XFILLER_9_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput534 wire1086/X vssd vssd vccd vccd la_data_in_core[49] sky130_fd_sc_hd__buf_8
Xoutput545 wire1076/X vssd vssd vccd vccd la_data_in_core[59] sky130_fd_sc_hd__buf_8
Xoutput556 _438_/X vssd vssd vccd vccd la_data_in_core[69] sky130_fd_sc_hd__buf_8
XFILLER_5_3308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput567 _448_/X vssd vssd vccd vccd la_data_in_core[79] sky130_fd_sc_hd__buf_8
XFILLER_5_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput578 wire1067/X vssd vssd vccd vccd la_data_in_core[89] sky130_fd_sc_hd__buf_8
Xoutput589 _468_/X vssd vssd vccd vccd la_data_in_core[99] sky130_fd_sc_hd__buf_8
Xwire1309 wire1309/A vssd vssd vccd vccd wire1309/X sky130_fd_sc_hd__buf_6
XFILLER_25_1834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[3\]_B _166_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__076__A _076_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[66\]_A la_data_out_core[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__523__B _523_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_936 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input245_A la_iena_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2056 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input412_A mprj_adr_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__495__A_N _623_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_121 mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 _197_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_143 _565_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _329_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_165 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_425_ _553_/A _425_/B _425_/C vssd vssd vccd vccd _425_/X sky130_fd_sc_hd__and3b_4
XTAP_2497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_356_ _356_/A _356_/B vssd vssd vccd vccd _356_/X sky130_fd_sc_hd__and2_4
XFILLER_35_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[57\]_A la_data_out_core[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_287_ _287_/A _287_/B vssd vssd vccd vccd _287_/X sky130_fd_sc_hd__and2_4
XANTENNA__433__B _433_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output464_A wire1059/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output631_A _003_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output729_A _606_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput5 la_data_out_mprj[100] vssd vssd vccd vccd _469_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1527_A wire1527/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__608__B _608_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[48\]_A la_data_out_core[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__624__A _624_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__343__B _343_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_max_cap1247_A wire1248/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1106 _398_/X vssd vssd vccd vccd wire1106/X sky130_fd_sc_hd__buf_6
XFILLER_25_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1117 _366_/X vssd vssd vccd vccd wire1117/X sky130_fd_sc_hd__buf_6
Xwire1128 wire1129/X vssd vssd vccd vccd wire1128/X sky130_fd_sc_hd__buf_6
XFILLER_38_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1139 _355_/X vssd vssd vccd vccd wire1139/X sky130_fd_sc_hd__buf_6
XFILLER_19_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__518__B _518_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_210_ _210_/A _210_/B vssd vssd vccd vccd _210_/X sky130_fd_sc_hd__and2_2
XFILLER_14_3460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[39\]_A la_data_out_core[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[123\]_A la_data_out_core[123] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__534__A _534_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_141_ _141_/A vssd vssd vccd vccd _141_/Y sky130_fd_sc_hd__inv_4
XANTENNA_input195_A la_iena_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__253__B _253_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_072_ _072_/A vssd vssd vccd vccd _072_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_13_1056 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input362_A la_oenb_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2719 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input56_A la_data_out_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3683 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1640 wire1640/A vssd vssd vccd vccd _507_/B sky130_fd_sc_hd__buf_6
Xwire1651 wire1652/X vssd vssd vccd vccd _496_/B sky130_fd_sc_hd__buf_6
Xwire1662 wire1663/X vssd vssd vccd vccd _491_/B sky130_fd_sc_hd__buf_6
Xwire1673 wire1673/A vssd vssd vccd vccd wire1673/X sky130_fd_sc_hd__buf_6
XFILLER_19_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1684 wire1685/X vssd vssd vccd vccd _480_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1695 wire1695/A vssd vssd vccd vccd wire1695/X sky130_fd_sc_hd__buf_6
XFILLER_19_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__428__B _428_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_408_ _536_/A _408_/B _408_/C vssd vssd vccd vccd _408_/X sky130_fd_sc_hd__and3b_2
XFILLER_15_2534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1010_A wire1011/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output581_A wire1065/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output679_A _047_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[114\]_A la_data_out_core[114] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_32_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_339_ _339_/A _339_/B vssd vssd vccd vccd _339_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire970 _130_/Y vssd vssd vccd vccd wire970/X sky130_fd_sc_hd__buf_6
XANTENNA_output846_A _506_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire981 _119_/Y vssd vssd vccd vccd wire981/X sky130_fd_sc_hd__buf_6
Xwire992 wire992/A vssd vssd vccd vccd _123_/A sky130_fd_sc_hd__buf_8
XFILLER_31_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1477_A wire1478/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[93\] la_data_out_core[93] wire1261/X vssd vssd vccd vccd _076_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_41_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1644_A wire1644/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__619__A _619_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__338__B _338_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_10 _317_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_854 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_21 _196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_342 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[105\]_A la_data_out_core[105] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_32 _613_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__354__A _354_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_43 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_54 _270_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_65 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_76 _187_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_87 _168_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_98 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1218 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3475 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2162 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__529__A _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__248__B _248_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input110_A la_data_out_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input208_A la_iena_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__264__A _264_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_124_ _124_/A vssd vssd vccd vccd _124_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_32_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_055_ _055_/A vssd vssd vccd vccd _055_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__430__C _430_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1058_A _471_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1470 wire1471/X vssd vssd vccd vccd _293_/A sky130_fd_sc_hd__buf_6
XFILLER_39_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1481 wire1481/A vssd vssd vccd vccd _287_/A sky130_fd_sc_hd__buf_6
XFILLER_46_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1492 wire1492/A vssd vssd vccd vccd _278_/A sky130_fd_sc_hd__buf_6
XFILLER_21_2593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1225_A _306_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output796_A _551_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1310 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__174__A _174_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[21\] mprj_dat_i_user[21] split13/X vssd vssd vccd vccd wire1016/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_30_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1594_A wire1594/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput30 la_data_out_mprj[123] vssd vssd vccd vccd _492_/C sky130_fd_sc_hd__clkbuf_4
Xinput41 la_data_out_mprj[18] vssd vssd vccd vccd _387_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput52 la_data_out_mprj[28] vssd vssd vccd vccd _397_/C sky130_fd_sc_hd__clkbuf_4
Xinput63 la_data_out_mprj[38] vssd vssd vccd vccd _407_/C sky130_fd_sc_hd__clkbuf_4
Xinput74 la_data_out_mprj[48] vssd vssd vccd vccd _417_/C sky130_fd_sc_hd__clkbuf_4
Xinput85 la_data_out_mprj[58] vssd vssd vccd vccd _427_/C sky130_fd_sc_hd__clkbuf_4
Xinput96 la_data_out_mprj[68] vssd vssd vccd vccd _437_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_2725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__621__B _621_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2758 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__406__A_N _534_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__349__A _349_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__531__B _531_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input158_A la_iena_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput401 mprj_adr_o_core[21] vssd vssd vccd vccd wire1388/A sky130_fd_sc_hd__buf_6
Xinput412 mprj_adr_o_core[31] vssd vssd vccd vccd wire1364/A sky130_fd_sc_hd__buf_6
Xinput423 mprj_dat_o_core[11] vssd vssd vccd vccd wire1337/A sky130_fd_sc_hd__buf_6
Xinput434 mprj_dat_o_core[21] vssd vssd vccd vccd wire1315/A sky130_fd_sc_hd__buf_6
XFILLER_40_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput445 mprj_dat_o_core[31] vssd vssd vccd vccd wire1293/A sky130_fd_sc_hd__buf_6
XFILLER_40_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput456 mprj_sel_o_core[2] vssd vssd vccd vccd wire1272/A sky130_fd_sc_hd__buf_6
XFILLER_22_3592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input325_A la_oenb_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__259__A _259_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input19_A la_data_out_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__425__C _425_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_107_ _107_/A vssd vssd vccd vccd _107_/Y sky130_fd_sc_hd__inv_2
Xoutput908 wire981/X vssd vssd vccd vccd mprj_dat_i_core[5] sky130_fd_sc_hd__buf_8
XFILLER_45_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput919 wire1144/X vssd vssd vccd vccd mprj_dat_o_user[15] sky130_fd_sc_hd__buf_8
XANTENNA__429__A_N _557_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_038_ _038_/A vssd vssd vccd vccd _038_/Y sky130_fd_sc_hd__inv_2
XANTENNA__441__B _441_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output544_A wire1077/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1175_A _337_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output711_A _076_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output809_A _563_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1342_A wire1343/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__169__A _169_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[56\] la_data_out_core[56] _219_/X vssd vssd vccd vccd _039_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_1_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1607_A wire1607/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__616__B _616_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_3306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__351__B _351_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__079__A _079_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__526__B _526_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__542__A _542_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input275_A la_oenb_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_rebuffer11_A wire1245/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input442_A mprj_dat_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput220 la_iena_mprj[64] vssd vssd vccd vccd _227_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput231 la_iena_mprj[74] vssd vssd vccd vccd _237_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput242 la_iena_mprj[84] vssd vssd vccd vccd _247_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput253 la_iena_mprj[94] vssd vssd vccd vccd _257_/B sky130_fd_sc_hd__clkbuf_4
Xinput264 la_oenb_mprj[103] vssd vssd vccd vccd _600_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput275 la_oenb_mprj[113] vssd vssd vccd vccd _610_/A sky130_fd_sc_hd__buf_4
XFILLER_2_3483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput286 la_oenb_mprj[123] vssd vssd vccd vccd _620_/A sky130_fd_sc_hd__clkbuf_4
Xinput297 la_oenb_mprj[18] vssd vssd vccd vccd _515_/A sky130_fd_sc_hd__buf_4
XFILLER_40_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_587_ _587_/A _587_/B vssd vssd vccd vccd _587_/X sky130_fd_sc_hd__and2_4
XFILLER_32_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__436__B _436_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output494_A _381_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output661_A _031_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output759_A _517_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1292_A wire1293/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput705 _071_/Y vssd vssd vccd vccd la_data_in_mprj[88] sky130_fd_sc_hd__buf_8
XANTENNA__171__B _171_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput716 _081_/Y vssd vssd vccd vccd la_data_in_mprj[98] sky130_fd_sc_hd__buf_8
XFILLER_29_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput727 _604_/X vssd vssd vccd vccd la_oenb_core[107] sky130_fd_sc_hd__buf_8
Xoutput738 _614_/X vssd vssd vccd vccd la_oenb_core[117] sky130_fd_sc_hd__buf_8
XFILLER_7_4051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput749 wire1032/X vssd vssd vccd vccd la_oenb_core[127] sky130_fd_sc_hd__buf_8
XANTENNA_output926_A wire1132/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1557_A wire1557/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3236 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1724_A wire1724/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__346__B _346_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[93\]_B wire1261/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__362__A _362_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_510_ _510_/A _510_/B vssd vssd vccd vccd _510_/X sky130_fd_sc_hd__and2_4
XTAP_2602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_441_ _569_/A _441_/B _441_/C vssd vssd vccd vccd _441_/X sky130_fd_sc_hd__and3b_4
XANTENNA__537__A _537_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_372_ _500_/A _372_/B _372_/C vssd vssd vccd vccd _372_/X sky130_fd_sc_hd__and3b_4
XTAP_1967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input392_A mprj_adr_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_790 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_B _247_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_2654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input86_A la_data_out_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1699 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__272__A _272_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output507_A _393_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1138_A wire1139/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__166__B _166_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1305_A wire1305/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output876_A wire1219/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[19\] la_data_out_core[19] _182_/X vssd vssd vccd vccd _002_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_32_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[75\]_B _238_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__182__A _182_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1674_A wire1675/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput502 _370_/X vssd vssd vccd vccd la_data_in_core[1] sky130_fd_sc_hd__buf_8
Xoutput513 _371_/X vssd vssd vccd vccd la_data_in_core[2] sky130_fd_sc_hd__buf_8
XFILLER_44_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput524 _372_/X vssd vssd vccd vccd la_data_in_core[3] sky130_fd_sc_hd__buf_8
Xoutput535 _373_/X vssd vssd vccd vccd la_data_in_core[4] sky130_fd_sc_hd__buf_8
XFILLER_9_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput546 _374_/X vssd vssd vccd vccd la_data_in_core[5] sky130_fd_sc_hd__buf_8
Xoutput557 wire1111/X vssd vssd vccd vccd la_data_in_core[6] sky130_fd_sc_hd__buf_8
Xoutput568 _376_/X vssd vssd vccd vccd la_data_in_core[7] sky130_fd_sc_hd__buf_8
XFILLER_25_3259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput579 wire1110/X vssd vssd vccd vccd la_data_in_core[8] sky130_fd_sc_hd__buf_8
XFILLER_5_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__357__A _357_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1806 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[66\]_B _229_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_rebuffer9_A wire1245/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__092__A _092_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2182 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input140_A la_iena_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input238_A la_iena_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input405_A mprj_adr_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_100 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__267__A _267_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _295_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 _203_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _503_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_155 _268_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_166 _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_424_ _552_/A _424_/B _424_/C vssd vssd vccd vccd _424_/X sky130_fd_sc_hd__and3b_4
XFILLER_15_3428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_355_ _355_/A _355_/B vssd vssd vccd vccd _355_/X sky130_fd_sc_hd__and2_4
XFILLER_41_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[57\]_B _220_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_286_ _286_/A _286_/B vssd vssd vccd vccd _286_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__433__C _433_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output624_A _161_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput6 la_data_out_mprj[101] vssd vssd vccd vccd _470_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_20_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__177__A _177_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__624__B _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[0\] la_data_out_core[0] _625_/X vssd vssd vccd vccd _147_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_5_3139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_2563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1107 _397_/X vssd vssd vccd vccd wire1107/X sky130_fd_sc_hd__buf_6
Xwire1118 wire1119/X vssd vssd vccd vccd wire1118/X sky130_fd_sc_hd__buf_6
XFILLER_25_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1129 _360_/X vssd vssd vccd vccd wire1129/X sky130_fd_sc_hd__buf_6
XFILLER_38_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[39\]_B _202_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_140_ _140_/A vssd vssd vccd vccd _140_/Y sky130_fd_sc_hd__inv_4
XANTENNA_user_to_mprj_in_gates\[123\]_B _286_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__534__B _534_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1614 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_071_ _071_/A vssd vssd vccd vccd _071_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_32_1669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input188_A la_iena_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__550__A _550_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input355_A la_oenb_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__462__A_N _590_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input49_A la_data_out_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1630 wire1630/A vssd vssd vccd vccd _520_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1641 wire1641/A vssd vssd vccd vccd _506_/B sky130_fd_sc_hd__buf_6
Xwire1652 wire1652/A vssd vssd vccd vccd wire1652/X sky130_fd_sc_hd__buf_6
XFILLER_46_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1663 wire1663/A vssd vssd vccd vccd wire1663/X sky130_fd_sc_hd__buf_6
Xwire1674 wire1675/X vssd vssd vccd vccd _485_/B sky130_fd_sc_hd__buf_6
Xwire1685 wire1685/A vssd vssd vccd vccd wire1685/X sky130_fd_sc_hd__buf_6
XFILLER_19_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1696 wire1696/A vssd vssd vccd vccd _473_/B sky130_fd_sc_hd__buf_6
XFILLER_19_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__428__C _428_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_407_ _535_/A _407_/B _407_/C vssd vssd vccd vccd _407_/X sky130_fd_sc_hd__and3b_2
XTAP_1572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_338_ _338_/A _338_/B vssd vssd vccd vccd _338_/X sky130_fd_sc_hd__and2_2
XANTENNA__444__B _444_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[114\]_B _277_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1003_A wire1004/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output574_A _454_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_269_ _269_/A _269_/B vssd vssd vccd vccd _269_/X sky130_fd_sc_hd__and2_2
Xwire971 _129_/Y vssd vssd vccd vccd wire971/X sky130_fd_sc_hd__buf_6
XFILLER_10_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire982 _118_/Y vssd vssd vccd vccd wire982/X sky130_fd_sc_hd__buf_6
Xwire993 wire993/A vssd vssd vccd vccd _122_/A sky130_fd_sc_hd__buf_8
XANTENNA_output741_A _508_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output839_A _590_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1372_A wire1373/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[86\] la_data_out_core[86] _249_/X vssd vssd vccd vccd _069_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1637_A wire1637/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_966 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__619__B _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[23\]_A mprj_dat_i_user[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire992_A wire992/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_11 _317_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_22 _196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[105\]_B wire1252/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__354__B _354_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_33 _622_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_44 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_55 _270_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_66 _267_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_77 _186_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_88 _168_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_99 _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__485__A_N _613_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__529__B _529_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[14\]_A mprj_dat_i_user[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input103_A la_data_out_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__545__A _545_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_682 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_123_ _123_/A vssd vssd vccd vccd _123_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_10_3144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_054_ _054_/A vssd vssd vccd vccd _054_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_2454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__280__A _280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1460 wire1461/X vssd vssd vccd vccd _371_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1471 wire1471/A vssd vssd vccd vccd wire1471/X sky130_fd_sc_hd__buf_6
XANTENNA__439__B _439_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1482 wire1482/A vssd vssd vccd vccd _286_/A sky130_fd_sc_hd__buf_6
Xwire1493 wire1493/A vssd vssd vccd vccd _277_/A sky130_fd_sc_hd__buf_6
XFILLER_34_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1120_A wire1121/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1218_A _312_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output691_A _058_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1322 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output789_A _545_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__174__B _174_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output956_A wire1241/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[14\] mprj_dat_i_user[14] rebuffer12/X vssd vssd vccd vccd wire1025/A
+ sky130_fd_sc_hd__nand2_8
Xinput20 la_data_out_mprj[114] vssd vssd vccd vccd _483_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput31 la_data_out_mprj[124] vssd vssd vccd vccd _493_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1587_A wire1588/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput42 la_data_out_mprj[19] vssd vssd vccd vccd _388_/C sky130_fd_sc_hd__clkbuf_4
Xinput53 la_data_out_mprj[29] vssd vssd vccd vccd _398_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput64 la_data_out_mprj[39] vssd vssd vccd vccd _408_/C sky130_fd_sc_hd__clkbuf_4
Xinput75 la_data_out_mprj[49] vssd vssd vccd vccd _418_/C sky130_fd_sc_hd__clkbuf_4
Xinput86 la_data_out_mprj[59] vssd vssd vccd vccd _428_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__190__A _190_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput97 la_data_out_mprj[69] vssd vssd vccd vccd _438_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[112\] la_data_out_core[112] _275_/X vssd vssd vccd vccd _095_/A
+ sky130_fd_sc_hd__nand2_4
XANTENNA__349__B _349_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__365__A _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput402 mprj_adr_o_core[22] vssd vssd vccd vccd wire1385/A sky130_fd_sc_hd__buf_6
Xinput413 mprj_adr_o_core[3] vssd vssd vccd vccd wire1362/A sky130_fd_sc_hd__buf_6
Xinput424 mprj_dat_o_core[12] vssd vssd vccd vccd wire1335/A sky130_fd_sc_hd__buf_6
XFILLER_2_3632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput435 mprj_dat_o_core[22] vssd vssd vccd vccd wire1313/A sky130_fd_sc_hd__buf_6
Xinput446 mprj_dat_o_core[3] vssd vssd vccd vccd wire1291/A sky130_fd_sc_hd__buf_6
XFILLER_0_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput457 mprj_sel_o_core[3] vssd vssd vccd vccd wire1270/A sky130_fd_sc_hd__buf_6
XFILLER_29_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input220_A la_iena_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input318_A la_oenb_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__275__A _275_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_106_ _106_/A vssd vssd vccd vccd _106_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_9_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput909 wire980/X vssd vssd vccd vccd mprj_dat_i_core[6] sky130_fd_sc_hd__buf_8
X_037_ _037_/A vssd vssd vccd vccd _037_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__441__C _441_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output537_A wire1084/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1168_A wire1169/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output704_A _070_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__169__B _169_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1335_A wire1335/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1290 wire1291/X vssd vssd vccd vccd _340_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[49\] la_data_out_core[49] _212_/X vssd vssd vccd vccd _032_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_34_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_906 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1502_A wire1502/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__185__A _185_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2374 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__542__B _542_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input170_A la_iena_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input268_A la_oenb_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2044 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input435_A mprj_dat_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput210 la_iena_mprj[55] vssd vssd vccd vccd _218_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input31_A la_data_out_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput221 la_iena_mprj[65] vssd vssd vccd vccd _228_/B sky130_fd_sc_hd__clkbuf_4
Xinput232 la_iena_mprj[75] vssd vssd vccd vccd _238_/B sky130_fd_sc_hd__clkbuf_4
Xinput243 la_iena_mprj[85] vssd vssd vccd vccd _248_/B sky130_fd_sc_hd__clkbuf_4
Xinput254 la_iena_mprj[95] vssd vssd vccd vccd _258_/B sky130_fd_sc_hd__clkbuf_4
Xinput265 la_oenb_mprj[104] vssd vssd vccd vccd _601_/A sky130_fd_sc_hd__buf_4
XFILLER_40_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput276 la_oenb_mprj[114] vssd vssd vccd vccd _611_/A sky130_fd_sc_hd__clkbuf_4
Xinput287 la_oenb_mprj[124] vssd vssd vccd vccd _621_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput298 la_oenb_mprj[19] vssd vssd vccd vccd _516_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_586_ _586_/A _586_/B vssd vssd vccd vccd _586_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__436__C _436_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output487_A _490_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__452__B _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output654_A _024_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput706 _072_/Y vssd vssd vccd vccd la_data_in_mprj[89] sky130_fd_sc_hd__buf_8
Xoutput717 wire990/X vssd vssd vccd vccd la_data_in_mprj[99] sky130_fd_sc_hd__buf_8
XFILLER_9_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput728 wire1043/X vssd vssd vccd vccd la_oenb_core[108] sky130_fd_sc_hd__buf_8
XANTENNA_wire1285_A wire1285/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput739 wire1039/X vssd vssd vccd vccd la_oenb_core[118] sky130_fd_sc_hd__buf_8
XFILLER_7_4063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output821_A _574_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output919_A wire1144/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1452_A wire1453/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1717_A wire1717/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__362__B _362_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[6\]_A mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[6\]_A la_data_out_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_440_ _568_/A _440_/B _440_/C vssd vssd vccd vccd _440_/X sky130_fd_sc_hd__and3b_1
XANTENNA__537__B _537_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__419__A_N _547_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_371_ _499_/A _371_/B _371_/C vssd vssd vccd vccd _371_/X sky130_fd_sc_hd__and3b_4
XFILLER_18_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__553__A _553_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input385_A la_oenb_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input79_A la_data_out_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__447__B _447_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_569_ _569_/A _569_/B vssd vssd vccd vccd _569_/X sky130_fd_sc_hd__and2_4
XFILLER_18_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1200_A _324_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output771_A _528_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output869_A wire1180/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput503 _389_/X vssd vssd vccd vccd la_data_in_core[20] sky130_fd_sc_hd__buf_8
Xoutput514 wire1105/X vssd vssd vccd vccd la_data_in_core[30] sky130_fd_sc_hd__buf_8
Xoutput525 wire1095/X vssd vssd vccd vccd la_data_in_core[40] sky130_fd_sc_hd__buf_8
XFILLER_25_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput536 wire1085/X vssd vssd vccd vccd la_data_in_core[50] sky130_fd_sc_hd__buf_8
XFILLER_29_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput547 wire1075/X vssd vssd vccd vccd la_data_in_core[60] sky130_fd_sc_hd__buf_8
XFILLER_9_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput558 wire1069/X vssd vssd vccd vccd la_data_in_core[70] sky130_fd_sc_hd__buf_8
Xoutput569 _449_/X vssd vssd vccd vccd la_data_in_core[80] sky130_fd_sc_hd__buf_8
XFILLER_25_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__357__B _357_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2194 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input133_A la_iena_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__548__A _548_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_112 _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input300_A la_oenb_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_123 _295_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _203_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _589_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _268_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 _171_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_423_ _551_/A _423_/B _423_/C vssd vssd vccd vccd _423_/X sky130_fd_sc_hd__and3b_2
XFILLER_14_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__391__A_N _519_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_354_ _354_/A _354_/B vssd vssd vccd vccd _354_/X sky130_fd_sc_hd__and2_4
XFILLER_35_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__283__A _283_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_285_ _285_/A _285_/B vssd vssd vccd vccd _285_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output617_A _106_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1150_A wire1151/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput7 la_data_out_mprj[102] vssd vssd vccd vccd _471_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1248_A wire1249/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1415_A wire1416/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[31\] la_data_out_core[31] _194_/X vssd vssd vccd vccd _014_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_17_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__193__A _193_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1108 _396_/X vssd vssd vccd vccd wire1108/X sky130_fd_sc_hd__buf_6
Xwire1119 _365_/X vssd vssd vccd vccd wire1119/X sky130_fd_sc_hd__buf_6
XFILLER_25_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__368__A _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1626 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_070_ _070_/A vssd vssd vccd vccd _070_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_32_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input250_A la_iena_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input348_A la_oenb_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1620 wire1620/A vssd vssd vccd vccd _575_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1631 wire1631/A vssd vssd vccd vccd _518_/B sky130_fd_sc_hd__buf_6
Xwire1642 wire1642/A vssd vssd vccd vccd _505_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1653 wire1654/X vssd vssd vccd vccd _495_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__278__A _278_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1664 wire1665/X vssd vssd vccd vccd _490_/B sky130_fd_sc_hd__buf_6
Xwire1675 wire1675/A vssd vssd vccd vccd wire1675/X sky130_fd_sc_hd__buf_6
XFILLER_46_433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1686 wire1686/A vssd vssd vccd vccd _479_/B sky130_fd_sc_hd__buf_6
Xwire1697 wire1697/A vssd vssd vccd vccd _472_/B sky130_fd_sc_hd__buf_6
XFILLER_19_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_406_ _534_/A _406_/B _406_/C vssd vssd vccd vccd _406_/X sky130_fd_sc_hd__and3b_2
XFILLER_14_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_337_ _337_/A _337_/B vssd vssd vccd vccd _337_/X sky130_fd_sc_hd__and2_2
XANTENNA__444__C _444_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_268_ _268_/A _268_/B vssd vssd vccd vccd _268_/X sky130_fd_sc_hd__and2_1
XFILLER_10_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output567_A _448_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire961 _146_/Y vssd vssd vccd vccd wire961/X sky130_fd_sc_hd__buf_8
Xwire972 _128_/Y vssd vssd vccd vccd wire972/X sky130_fd_sc_hd__buf_6
Xwire983 _117_/Y vssd vssd vccd vccd wire983/X sky130_fd_sc_hd__buf_8
Xwire994 wire994/A vssd vssd vccd vccd _121_/A sky130_fd_sc_hd__buf_8
X_199_ _199_/A _199_/B vssd vssd vccd vccd _199_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1198_A _325_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__460__B _460_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output734_A _610_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1365_A wire1366/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output901_A _142_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[79\] la_data_out_core[79] _242_/X vssd vssd vccd vccd _062_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_26_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1532_A wire1532/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__188__A _188_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[23\]_B split13/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire985_A _115_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_12 _552_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_23 _196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_34 _499_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_45 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_56 _270_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_67 _267_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_78 _186_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_89 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__370__B _370_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__098__A _098_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__545__B _545_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input298_A la_oenb_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_366 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_122_ _122_/A vssd vssd vccd vccd _122_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_7_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__561__A _561_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_053_ _053_/A vssd vssd vccd vccd _053_/Y sky130_fd_sc_hd__inv_4
XFILLER_7_3703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input61_A la_data_out_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1450 wire1451/X vssd vssd vccd vccd _376_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1461 wire1461/A vssd vssd vccd vccd wire1461/X sky130_fd_sc_hd__buf_6
Xwire1472 wire1473/X vssd vssd vccd vccd _292_/A sky130_fd_sc_hd__buf_6
XANTENNA__439__C _439_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1483 wire1483/A vssd vssd vccd vccd _285_/A sky130_fd_sc_hd__buf_6
Xwire1494 wire1494/A vssd vssd vccd vccd _276_/A sky130_fd_sc_hd__buf_6
XFILLER_19_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_926 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__455__B _455_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1113_A _368_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output684_A _052_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput10 la_data_out_mprj[105] vssd vssd vccd vccd _474_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_output851_A wire1208/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput21 la_data_out_mprj[115] vssd vssd vccd vccd _484_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput32 la_data_out_mprj[125] vssd vssd vccd vccd _494_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_output949_A wire1237/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput43 la_data_out_mprj[1] vssd vssd vccd vccd _370_/C sky130_fd_sc_hd__clkbuf_4
Xinput54 la_data_out_mprj[2] vssd vssd vccd vccd _371_/C sky130_fd_sc_hd__clkbuf_4
Xinput65 la_data_out_mprj[3] vssd vssd vccd vccd _372_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1482_A wire1482/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput76 la_data_out_mprj[4] vssd vssd vccd vccd _373_/C sky130_fd_sc_hd__clkbuf_4
Xinput87 la_data_out_mprj[5] vssd vssd vccd vccd _374_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_2705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput98 la_data_out_mprj[6] vssd vssd vccd vccd _375_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_45_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[105\] la_data_out_core[105] wire1252/X vssd vssd vccd vccd
+ _088_/A sky130_fd_sc_hd__nand2_4
XFILLER_17_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj2_logic_high_inst wire1732/A vccd2_uq0 vssd2_uq0 mprj2_logic_high
XFILLER_11_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__365__B _365_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__452__A_N _580_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput403 mprj_adr_o_core[23] vssd vssd vccd vccd wire1383/A sky130_fd_sc_hd__buf_6
XFILLER_44_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput414 mprj_adr_o_core[4] vssd vssd vccd vccd wire1359/A sky130_fd_sc_hd__buf_6
XFILLER_2_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput425 mprj_dat_o_core[13] vssd vssd vccd vccd wire1333/A sky130_fd_sc_hd__buf_6
XFILLER_0_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput436 mprj_dat_o_core[23] vssd vssd vccd vccd wire1311/A sky130_fd_sc_hd__buf_6
Xinput447 mprj_dat_o_core[4] vssd vssd vccd vccd wire1289/A sky130_fd_sc_hd__buf_6
XFILLER_40_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput458 mprj_stb_o_core vssd vssd vccd vccd wire1268/A sky130_fd_sc_hd__buf_6
XFILLER_2_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_712 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input213_A la_iena_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__556__A _556_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__275__B _275_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__291__A _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_105_ _105_/A vssd vssd vccd vccd _105_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_036_ _036_/A vssd vssd vccd vccd _036_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2876 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_2646 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1280 wire1281/X vssd vssd vccd vccd _345_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1291 wire1291/A vssd vssd vccd vccd wire1291/X sky130_fd_sc_hd__buf_6
XANTENNA_wire1230_A _303_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1328_A wire1329/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__475__A_N _603_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output899_A _140_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_918 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__185__B _185_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1697_A wire1697/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xmprj_logic_high_inst _295_/B _395_/B _396_/B _397_/B _398_/B _399_/B _400_/B _401_/B
+ _402_/B _403_/B _404_/B _305_/A _405_/B _406_/B _407_/B _408_/B _409_/B _410_/B
+ _411_/B _412_/B _413_/B _414_/B _306_/A _415_/B _416_/B _417_/B _418_/B _419_/B
+ _420_/B _421_/B _422_/B _423_/B _424_/B _307_/A _425_/B _426_/B _427_/B _428_/B
+ _429_/B _430_/B _431_/B _432_/B _433_/B _434_/B _308_/A _435_/B _436_/B _437_/B
+ _438_/B _439_/B _440_/B wire1728/A wire1727/A wire1726/A wire1725/A _309_/A wire1724/A
+ wire1723/A wire1722/A wire1721/A wire1720/A wire1719/A wire1718/A wire1717/A wire1716/A
+ wire1715/A _310_/A wire1714/A wire1713/A wire1712/A wire1711/A wire1710/A wire1709/A
+ wire1708/A wire1707/A wire1706/A wire1705/A _311_/A wire1704/A wire1703/A wire1702/A
+ wire1701/A wire1700/A wire1699/A wire1698/A wire1697/A wire1696/A wire1695/A _312_/A
+ wire1693/A wire1692/A wire1690/A wire1688/A wire1686/A wire1685/A wire1683/A wire1681/A
+ wire1679/A wire1677/A _313_/A wire1675/A wire1673/A wire1671/A wire1669/A wire1667/A
+ wire1665/A wire1663/A wire1661/A wire1659/A wire1657/A _314_/A wire1655/A wire1654/A
+ wire1652/A wire1650/A wire1649/A wire1648/A wire1647/A wire1646/A wire1645/A wire1644/A
+ wire1643/A _315_/A wire1642/A wire1641/A wire1640/A wire1639/A wire1638/A wire1637/A
+ wire1636/A wire1635/A wire1634/A wire1633/A _316_/A wire1632/A _516_/B _517_/B wire1631/A
+ _519_/B wire1630/A wire1629/A _522_/B _523_/B wire1628/A _317_/A _525_/B _526_/B
+ _527_/B wire1627/A _529_/B _530_/B _531_/B _532_/B _533_/B _534_/B _318_/A _535_/B
+ _536_/B _537_/B _538_/B _539_/B _540_/B _541_/B _542_/B _543_/B _544_/B _319_/A
+ _545_/B _546_/B _547_/B _548_/B _549_/B _550_/B _551_/B _552_/B _553_/B _554_/B
+ _320_/A _555_/B _556_/B _557_/B _558_/B _559_/B _560_/B _561_/B _562_/B _563_/B
+ _564_/B _321_/A _565_/B wire1626/A _567_/B wire1625/A wire1624/A _570_/B _571_/B
+ wire1623/A wire1622/A wire1621/A _322_/A wire1620/A _576_/B wire1619/A wire1618/A
+ wire1617/A wire1616/A wire1615/A wire1614/A wire1613/A wire1612/A _323_/A wire1611/A
+ wire1610/A wire1609/A wire1608/A wire1607/A wire1606/A wire1605/A wire1604/A wire1603/A
+ wire1602/A _324_/A wire1601/A wire1598/A wire1597/A wire1596/A wire1595/A wire1594/A
+ wire1593/A wire1592/A wire1591/A wire1590/A wire1589/A _325_/A wire1588/A wire1586/A
+ wire1585/A wire1583/A wire1582/A wire1581/A wire1579/A wire1577/A wire1575/A wire1573/A
+ _326_/A wire1571/A wire1569/A wire1567/A wire1565/A wire1563/A wire1561/A wire1559/A
+ wire1557/A wire1555/A wire1553/A _327_/A wire1551/A wire1550/A wire1549/A wire1548/A
+ wire1547/A wire1546/A wire1545/A wire1544/A wire1543/A wire1542/A _328_/A wire1541/A
+ wire1540/A wire1539/A wire1538/A wire1537/A wire1536/A wire1535/A wire1534/A wire1533/A
+ wire1532/A _329_/A wire1531/A wire1530/A wire1529/A wire1528/A wire1527/A wire1526/A
+ wire1525/A wire1524/A wire1523/A wire1522/A _330_/A wire1521/A _194_/A _195_/A _196_/A
+ _197_/A _198_/A _199_/A _200_/A _201_/A _202_/A _331_/A _203_/A _204_/A _205_/A
+ _206_/A _207_/A _208_/A _209_/A _210_/A _211_/A _212_/A _332_/A _213_/A _214_/A
+ _215_/A _216_/A _217_/A _218_/A _219_/A _220_/A _221_/A _222_/A _333_/A _223_/A
+ _224_/A _225_/A _226_/A _227_/A _228_/A _229_/A _230_/A _231_/A _232_/A _334_/A
+ _298_/A _233_/A wire1520/A _235_/A _236_/A _237_/A _238_/A _239_/A _240_/A _241_/A
+ _242_/A _335_/A _243_/A wire1519/A _245_/A _246_/A _247_/A _248_/A wire1518/A wire1517/A
+ _251_/A wire1516/A _336_/A wire1515/A _254_/A _255_/A wire1514/A wire1513/A wire1512/A
+ wire1511/A wire1510/A wire1509/A wire1508/A _337_/A wire1507/A wire1506/A wire1505/A
+ wire1504/A wire1503/A wire1502/A wire1501/A wire1500/A wire1499/A wire1498/A _338_/A
+ wire1497/A wire1496/A wire1495/A wire1494/A wire1493/A wire1492/A wire1491/A wire1490/A
+ wire1489/A wire1488/A _339_/A wire1486/A wire1485/A wire1483/A wire1482/A wire1481/A
+ wire1480/A wire1478/A wire1476/A wire1475/A wire1473/A _340_/A wire1471/A wire1469/A
+ wire1466/A _341_/A _342_/A _343_/A _344_/A _299_/A _345_/A _346_/A _347_/A _348_/A
+ _349_/A _350_/A _351_/A _352_/A _353_/A _354_/A _300_/A _355_/A _356_/A _357_/A
+ _358_/A _359_/A _360_/A _361_/A _362_/A _363_/A _364_/A _301_/A _365_/A _366_/A
+ _367_/A _368_/A wire1465/A wire1463/A wire1461/A wire1459/A wire1457/A wire1455/A
+ _302_/A wire1453/A wire1451/A wire1449/A wire1447/A wire1445/A wire1443/A wire1441/A
+ wire1439/A wire1438/A wire1437/A _303_/A wire1436/A wire1435/A wire1434/A wire1433/A
+ wire1432/A wire1431/A wire1430/A wire1429/A wire1428/A wire1427/A _304_/A vccd1_uq1
+ vssd1_uq1 mprj_logic_high
XTAP_995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_A la_data_out_core[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input163_A la_iena_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[20\]_A la_data_out_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput200 la_iena_mprj[46] vssd vssd vccd vccd _209_/B sky130_fd_sc_hd__clkbuf_4
Xinput211 la_iena_mprj[56] vssd vssd vccd vccd _219_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput222 la_iena_mprj[66] vssd vssd vccd vccd _229_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput233 la_iena_mprj[76] vssd vssd vccd vccd _239_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_input330_A la_oenb_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input428_A mprj_dat_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput244 la_iena_mprj[86] vssd vssd vccd vccd _249_/B sky130_fd_sc_hd__clkbuf_4
Xinput255 la_iena_mprj[96] vssd vssd vccd vccd _259_/B sky130_fd_sc_hd__clkbuf_4
Xinput266 la_oenb_mprj[105] vssd vssd vccd vccd _602_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input24_A la_data_out_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput277 la_oenb_mprj[115] vssd vssd vccd vccd _612_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput288 la_oenb_mprj[125] vssd vssd vccd vccd _622_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput299 la_oenb_mprj[1] vssd vssd vccd vccd wire1424/A sky130_fd_sc_hd__buf_6
XFILLER_18_4128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__286__A _286_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_585_ _585_/A _585_/B vssd vssd vccd vccd _585_/X sky130_fd_sc_hd__and2_4
XFILLER_17_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[87\]_A la_data_out_core[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__452__C _452_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput707 _155_/Y vssd vssd vccd vccd la_data_in_mprj[8] sky130_fd_sc_hd__buf_8
Xoutput718 _156_/Y vssd vssd vccd vccd la_data_in_mprj[9] sky130_fd_sc_hd__buf_8
Xoutput729 _606_/X vssd vssd vccd vccd la_oenb_core[109] sky130_fd_sc_hd__buf_8
X_019_ _019_/A vssd vssd vccd vccd _019_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_2123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1180_A wire1181/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1278_A wire1279/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3280 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output814_A _567_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[11\]_A la_data_out_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[61\] la_data_out_core[61] _224_/X vssd vssd vccd vccd _044_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_23_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1612_A wire1612/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__196__A _196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[78\]_A la_data_out_core[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2218 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[6\]_B _169_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1296 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_370_ _498_/A _370_/B _370_/C vssd vssd vccd vccd _370_/X sky130_fd_sc_hd__and3b_4
XTAP_1947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[69\]_A la_data_out_core[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input280_A la_oenb_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input378_A la_oenb_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_958 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__447__C _447_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_568_ _568_/A _568_/B vssd vssd vccd vccd _568_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1026_A wire1026/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output597_A _088_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_499_ _499_/A _499_/B vssd vssd vccd vccd _499_/X sky130_fd_sc_hd__and2_4
XFILLER_31_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__463__B _463_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output764_A _522_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1395_A wire1395/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output931_A wire1122/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput504 _390_/X vssd vssd vccd vccd la_data_in_core[21] sky130_fd_sc_hd__buf_8
XFILLER_29_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput515 wire1104/X vssd vssd vccd vccd la_data_in_core[31] sky130_fd_sc_hd__buf_8
Xoutput526 wire1094/X vssd vssd vccd vccd la_data_in_core[41] sky130_fd_sc_hd__buf_8
Xoutput537 wire1084/X vssd vssd vccd vccd la_data_in_core[51] sky130_fd_sc_hd__buf_8
XFILLER_25_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput548 wire1074/X vssd vssd vccd vccd la_data_in_core[61] sky130_fd_sc_hd__buf_8
XFILLER_5_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1562_A wire1563/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput559 wire1068/X vssd vssd vccd vccd la_data_in_core[71] sky130_fd_sc_hd__buf_8
XFILLER_7_3171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__373__B _373_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1354 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__548__B _548_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input126_A la_data_out_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_113 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_124 _295_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _203_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 _590_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _268_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_422_ _550_/A _422_/B _422_/C vssd vssd vccd vccd _422_/X sky130_fd_sc_hd__and3b_4
XTAP_1722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _610_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[126\]_A la_data_out_core[126] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__564__A _564_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_353_ _353_/A _353_/B vssd vssd vccd vccd _353_/X sky130_fd_sc_hd__and2_4
XTAP_1788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input91_A la_data_out_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_284_ _284_/A _284_/B vssd vssd vccd vccd _284_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[7\] mprj_dat_i_user[7] rebuffer1/X vssd vssd vccd vccd wire994/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_3537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output512_A wire1106/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput8 la_data_out_mprj[103] vssd vssd vccd vccd _472_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__458__B _458_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1143_A _353_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1310_A wire1311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1408_A wire1409/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output881_A wire986/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_2342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[117\]_A la_data_out_core[117] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_33_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[24\] la_data_out_core[24] _187_/X vssd vssd vccd vccd _007_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_36_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__409__A_N _537_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2947 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1109 _395_/X vssd vssd vccd vccd wire1109/X sky130_fd_sc_hd__buf_6
XFILLER_45_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__368__B _368_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[108\]_A la_data_out_core[108] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_10_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2030 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2626 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput890 wire968/X vssd vssd vccd vccd mprj_dat_i_core[18] sky130_fd_sc_hd__buf_8
XFILLER_21_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input243_A la_iena_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1610 wire1610/A vssd vssd vccd vccd _586_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__559__A _559_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1621 wire1621/A vssd vssd vccd vccd _574_/B sky130_fd_sc_hd__buf_6
XFILLER_4_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1632 wire1632/A vssd vssd vccd vccd _515_/B sky130_fd_sc_hd__buf_6
XFILLER_19_604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1643 wire1643/A vssd vssd vccd vccd _504_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1654 wire1654/A vssd vssd vccd vccd wire1654/X sky130_fd_sc_hd__buf_6
XANTENNA_input410_A mprj_adr_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1665 wire1665/A vssd vssd vccd vccd wire1665/X sky130_fd_sc_hd__buf_6
XFILLER_24_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1676 wire1677/X vssd vssd vccd vccd _484_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1687 wire1688/X vssd vssd vccd vccd _478_/B sky130_fd_sc_hd__buf_6
Xwire1698 wire1698/A vssd vssd vccd vccd _471_/B sky130_fd_sc_hd__buf_6
XTAP_2220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__294__A _294_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_405_ _533_/A _405_/B _405_/C vssd vssd vccd vccd _405_/X sky130_fd_sc_hd__and3b_2
XTAP_1552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_336_ _336_/A _336_/B vssd vssd vccd vccd _336_/X sky130_fd_sc_hd__and2_2
XFILLER_15_2559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_267_ _267_/A _267_/B vssd vssd vccd vccd _267_/X sky130_fd_sc_hd__and2_1
Xwire962 _138_/Y vssd vssd vccd vccd wire962/X sky130_fd_sc_hd__buf_6
XFILLER_10_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire973 _127_/Y vssd vssd vccd vccd wire973/X sky130_fd_sc_hd__buf_6
Xwire984 _116_/Y vssd vssd vccd vccd wire984/X sky130_fd_sc_hd__buf_8
X_198_ _198_/A _198_/B vssd vssd vccd vccd _198_/X sky130_fd_sc_hd__and2_2
Xwire995 wire995/A vssd vssd vccd vccd _120_/A sky130_fd_sc_hd__buf_8
XFILLER_26_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__460__C _460_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1093_A _411_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output727_A _604_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1358_A wire1359/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1525_A wire1525/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_13 _552_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire978_A _122_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_24 _198_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_35 _367_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_46 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_57 _270_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_68 _267_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_378 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_79 _186_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__370__C _370_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__381__A_N _509_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_121_ _121_/A vssd vssd vccd vccd _121_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_36_1582 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input193_A la_iena_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_052_ _052_/A vssd vssd vccd vccd _052_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__561__B _561_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input360_A la_oenb_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input458_A mprj_stb_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input54_A la_data_out_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__289__A _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1440 wire1441/X vssd vssd vccd vccd _381_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1451 wire1451/A vssd vssd vccd vccd wire1451/X sky130_fd_sc_hd__buf_6
XFILLER_4_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1462 wire1463/X vssd vssd vccd vccd _370_/B sky130_fd_sc_hd__buf_6
XFILLER_19_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1473 wire1473/A vssd vssd vccd vccd wire1473/X sky130_fd_sc_hd__buf_6
Xwire1484 wire1485/X vssd vssd vccd vccd _284_/A sky130_fd_sc_hd__buf_6
XFILLER_46_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1495 wire1495/A vssd vssd vccd vccd _275_/A sky130_fd_sc_hd__buf_6
Xpowergood_check vccd vssd vdda1_uq0 vssa1_uq0 vdda2_uq0 vssa2_uq0 output954/A output952/A
+ mgmt_protect_hv
XFILLER_19_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_938 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__455__C _455_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output677_A _045_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_319_ _319_/A _319_/B vssd vssd vccd vccd _319_/X sky130_fd_sc_hd__and2_4
Xinput11 la_data_out_mprj[106] vssd vssd vccd vccd _475_/C sky130_fd_sc_hd__buf_4
Xinput22 la_data_out_mprj[116] vssd vssd vccd vccd _485_/C sky130_fd_sc_hd__clkbuf_4
Xinput33 la_data_out_mprj[126] vssd vssd vccd vccd _495_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__471__B _471_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput44 la_data_out_mprj[20] vssd vssd vccd vccd _389_/C sky130_fd_sc_hd__clkbuf_4
Xinput55 la_data_out_mprj[30] vssd vssd vccd vccd _399_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output844_A _595_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput66 la_data_out_mprj[40] vssd vssd vccd vccd _409_/C sky130_fd_sc_hd__clkbuf_4
Xinput77 la_data_out_mprj[50] vssd vssd vccd vccd _419_/C sky130_fd_sc_hd__clkbuf_4
Xinput88 la_data_out_mprj[60] vssd vssd vccd vccd _429_/C sky130_fd_sc_hd__clkbuf_4
Xinput99 la_data_out_mprj[70] vssd vssd vccd vccd _439_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_2717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1475_A wire1475/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[91\] la_data_out_core[91] _254_/X vssd vssd vccd vccd _074_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_26_2430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__199__A _199_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__381__B _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput404 mprj_adr_o_core[24] vssd vssd vccd vccd wire1381/A sky130_fd_sc_hd__buf_6
Xinput415 mprj_adr_o_core[5] vssd vssd vccd vccd wire1356/A sky130_fd_sc_hd__buf_6
XFILLER_0_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput426 mprj_dat_o_core[14] vssd vssd vccd vccd wire1331/A sky130_fd_sc_hd__buf_6
Xinput437 mprj_dat_o_core[24] vssd vssd vccd vccd wire1309/A sky130_fd_sc_hd__buf_6
Xinput448 mprj_dat_o_core[5] vssd vssd vccd vccd wire1287/A sky130_fd_sc_hd__buf_6
XFILLER_25_1250 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput459 mprj_we_o_core vssd vssd vccd vccd wire1266/A sky130_fd_sc_hd__buf_6
XFILLER_2_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__556__B _556_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input206_A la_iena_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2654 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__572__A _572_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_104_ _104_/A vssd vssd vccd vccd _104_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__291__B _291_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_035_ _035_/A vssd vssd vccd vccd _035_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1298 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1270 wire1270/A vssd vssd vccd vccd wire1270/X sky130_fd_sc_hd__buf_6
XFILLER_21_2371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1281 wire1281/A vssd vssd vccd vccd wire1281/X sky130_fd_sc_hd__buf_6
XFILLER_19_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1292 wire1293/X vssd vssd vccd vccd _368_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__466__B _466_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1223_A _308_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output794_A _549_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1592_A wire1592/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__376__B _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3664 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_B wire1259/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2540 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input156_A la_iena_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput201 la_iena_mprj[47] vssd vssd vccd vccd _210_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_gates\[20\]_B _183_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput212 la_iena_mprj[57] vssd vssd vccd vccd _220_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput223 la_iena_mprj[67] vssd vssd vccd vccd _230_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput234 la_iena_mprj[77] vssd vssd vccd vccd _240_/B sky130_fd_sc_hd__clkbuf_4
Xinput245 la_iena_mprj[87] vssd vssd vccd vccd _250_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput256 la_iena_mprj[97] vssd vssd vccd vccd _260_/B sky130_fd_sc_hd__clkbuf_4
Xinput267 la_oenb_mprj[106] vssd vssd vccd vccd _603_/A sky130_fd_sc_hd__buf_4
XANTENNA_input323_A la_oenb_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput278 la_oenb_mprj[116] vssd vssd vccd vccd _613_/A sky130_fd_sc_hd__clkbuf_4
Xinput289 la_oenb_mprj[126] vssd vssd vccd vccd _623_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_2741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__567__A _567_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input17_A la_data_out_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_584_ _584_/A _584_/B vssd vssd vccd vccd _584_/X sky130_fd_sc_hd__and2_4
XFILLER_16_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[87\]_B _250_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput708 _073_/Y vssd vssd vccd vccd la_data_in_mprj[90] sky130_fd_sc_hd__buf_8
XFILLER_29_2812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput719 _497_/X vssd vssd vccd vccd la_oenb_core[0] sky130_fd_sc_hd__buf_8
X_018_ _018_/A vssd vssd vccd vccd _018_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_2845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output542_A wire1079/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1173_A _338_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[11\]_B _174_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__442__A_N _570_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output807_A _561_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1340_A wire1341/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1438_A wire1438/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[54\] la_data_out_core[54] _217_/X vssd vssd vccd vccd _037_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_1_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1605_A wire1605/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[78\]_B _241_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input9_A la_data_out_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[69\]_B _232_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input273_A la_oenb_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__465__A_N _593_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input440_A mprj_dat_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__297__A _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_567_ _567_/A _567_/B vssd vssd vccd vccd _567_/X sky130_fd_sc_hd__and2_4
XFILLER_31_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_498_ _498_/A _498_/B vssd vssd vccd vccd _498_/X sky130_fd_sc_hd__and2_4
XANTENNA_output492_A wire1055/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1019_A wire1019/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output757_A _516_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1290_A wire1291/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput505 _391_/X vssd vssd vccd vccd la_data_in_core[22] sky130_fd_sc_hd__buf_8
XANTENNA_wire1388_A wire1388/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput516 wire1103/X vssd vssd vccd vccd la_data_in_core[32] sky130_fd_sc_hd__buf_8
Xoutput527 wire1093/X vssd vssd vccd vccd la_data_in_core[42] sky130_fd_sc_hd__buf_8
XFILLER_9_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput538 wire1083/X vssd vssd vccd vccd la_data_in_core[52] sky130_fd_sc_hd__buf_8
XANTENNA_output924_A wire1172/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput549 wire1073/X vssd vssd vccd vccd la_data_in_core[62] sky130_fd_sc_hd__buf_8
XFILLER_10_1190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1555_A wire1555/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__373__C _373_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1366 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__488__A_N _616_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 _600_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 wire1685/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input119_A la_data_out_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_136 _207_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_421_ _549_/A _421_/B _421_/C vssd vssd vccd vccd _421_/X sky130_fd_sc_hd__and3b_2
XTAP_1712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _368_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 _256_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_169 _599_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[126\]_B _289_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_352_ _352_/A _352_/B vssd vssd vccd vccd _352_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__564__B _564_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ _283_/A _283_/B vssd vssd vccd vccd _283_/X sky130_fd_sc_hd__and2_4
XANTENNA_input390_A mprj_adr_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input84_A la_data_out_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__580__A _580_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput9 la_data_out_mprj[104] vssd vssd vccd vccd _473_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_24_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__458__C _458_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output505_A _391_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1136_A wire1137/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_619_ _619_/A _619_/B vssd vssd vccd vccd _619_/X sky130_fd_sc_hd__and2_1
XFILLER_33_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__474__B _474_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[117\]_B _280_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output874_A wire1222/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[17\] la_data_out_core[17] _180_/X vssd vssd vccd vccd _000_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_20_549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1672_A wire1673/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2959 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[26\]_A mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__384__B _384_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[108\]_B _271_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_rebuffer7_A wire1248/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_3497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2638 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput880 wire1239/X vssd vssd vccd vccd mprj_cyc_o_user sky130_fd_sc_hd__buf_8
XFILLER_5_3632 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput891 wire967/X vssd vssd vccd vccd mprj_dat_i_core[19] sky130_fd_sc_hd__buf_8
XFILLER_8_1320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1600 wire1601/X vssd vssd vccd vccd wire1600/X sky130_fd_sc_hd__buf_6
Xwire1611 wire1611/A vssd vssd vccd vccd _585_/B sky130_fd_sc_hd__buf_6
XANTENNA__559__B _559_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input236_A la_iena_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1622 wire1622/A vssd vssd vccd vccd _573_/B sky130_fd_sc_hd__buf_6
XANTENNA_user_wb_dat_gates\[17\]_A mprj_dat_i_user[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1633 wire1633/A vssd vssd vccd vccd _514_/B sky130_fd_sc_hd__buf_6
XFILLER_4_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1644 wire1644/A vssd vssd vccd vccd _503_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1655 wire1655/A vssd vssd vccd vccd _296_/A sky130_fd_sc_hd__buf_6
Xwire1666 wire1667/X vssd vssd vccd vccd _489_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1677 wire1677/A vssd vssd vccd vccd wire1677/X sky130_fd_sc_hd__buf_6
XFILLER_24_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1688 wire1688/A vssd vssd vccd vccd wire1688/X sky130_fd_sc_hd__buf_6
XFILLER_41_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1699 wire1699/A vssd vssd vccd vccd _470_/B sky130_fd_sc_hd__buf_6
XANTENNA_input403_A mprj_adr_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__575__A _575_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__294__B _294_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_404_ _532_/A _404_/B _404_/C vssd vssd vccd vccd _404_/X sky130_fd_sc_hd__and3b_2
XPHY_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_2516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_335_ _335_/A _335_/B vssd vssd vccd vccd _335_/X sky130_fd_sc_hd__and2_2
XFILLER_30_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_266_ _266_/A _266_/B vssd vssd vccd vccd _266_/X sky130_fd_sc_hd__and2_1
XFILLER_32_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire963 _137_/Y vssd vssd vccd vccd wire963/X sky130_fd_sc_hd__buf_6
XFILLER_26_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire974 _126_/Y vssd vssd vccd vccd wire974/X sky130_fd_sc_hd__buf_6
X_197_ _197_/A _197_/B vssd vssd vccd vccd _197_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire985 _115_/Y vssd vssd vccd vccd wire985/X sky130_fd_sc_hd__buf_6
Xwire996 wire996/A vssd vssd vccd vccd _119_/A sky130_fd_sc_hd__buf_8
XFILLER_6_3407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__469__B _469_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1420_A wire1420/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_14 _553_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_25 _198_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_36 _314_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_47 _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_58 _270_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_69 _267_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__379__B _379_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_120_ _120_/A vssd vssd vccd vccd _120_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_36_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_051_ _051_/A vssd vssd vccd vccd _051_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input186_A la_iena_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input353_A la_oenb_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input47_A la_data_out_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1430 wire1430/A vssd vssd vccd vccd _391_/B sky130_fd_sc_hd__buf_6
Xwire1441 wire1441/A vssd vssd vccd vccd wire1441/X sky130_fd_sc_hd__buf_6
XFILLER_21_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1452 wire1453/X vssd vssd vccd vccd _375_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1463 wire1463/A vssd vssd vccd vccd wire1463/X sky130_fd_sc_hd__buf_6
Xwire1474 wire1475/X vssd vssd vccd vccd _291_/A sky130_fd_sc_hd__buf_6
XFILLER_1_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1485 wire1485/A vssd vssd vccd vccd wire1485/X sky130_fd_sc_hd__buf_6
Xwire1496 wire1496/A vssd vssd vccd vccd _274_/A sky130_fd_sc_hd__buf_6
XFILLER_46_265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_318_ _318_/A _318_/B vssd vssd vccd vccd _318_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1001_A wire1001/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output572_A _452_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput12 la_data_out_mprj[107] vssd vssd vccd vccd _476_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_30_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput23 la_data_out_mprj[117] vssd vssd vccd vccd _486_/C sky130_fd_sc_hd__clkbuf_4
Xinput34 la_data_out_mprj[127] vssd vssd vccd vccd _496_/C sky130_fd_sc_hd__clkbuf_4
X_249_ _249_/A _249_/B vssd vssd vccd vccd _249_/X sky130_fd_sc_hd__and2_4
Xinput45 la_data_out_mprj[21] vssd vssd vccd vccd _390_/C sky130_fd_sc_hd__clkbuf_4
Xinput56 la_data_out_mprj[31] vssd vssd vccd vccd _400_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput67 la_data_out_mprj[41] vssd vssd vccd vccd _410_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput78 la_data_out_mprj[51] vssd vssd vccd vccd _420_/C sky130_fd_sc_hd__clkbuf_4
Xinput89 la_data_out_mprj[61] vssd vssd vccd vccd _430_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_output837_A _588_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1370_A wire1371/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1468_A wire1469/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[84\] la_data_out_core[84] _247_/X vssd vssd vccd vccd _067_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_6_3259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_3893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__381__C _381_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput405 mprj_adr_o_core[25] vssd vssd vccd vccd wire1379/A sky130_fd_sc_hd__buf_6
XFILLER_2_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput416 mprj_adr_o_core[6] vssd vssd vccd vccd wire1353/A sky130_fd_sc_hd__buf_6
XFILLER_40_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput427 mprj_dat_o_core[15] vssd vssd vccd vccd wire1329/A sky130_fd_sc_hd__buf_6
XFILLER_2_3624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput438 mprj_dat_o_core[25] vssd vssd vccd vccd wire1307/A sky130_fd_sc_hd__buf_6
Xinput449 mprj_dat_o_core[6] vssd vssd vccd vccd wire1285/A sky130_fd_sc_hd__buf_6
XFILLER_29_711 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input101_A la_data_out_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__572__B _572_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_103_ _103_/A vssd vssd vccd vccd _103_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_034_ _034_/A vssd vssd vccd vccd _034_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3270 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1260 _258_/X vssd vssd vccd vccd wire1260/X sky130_fd_sc_hd__buf_6
XFILLER_23_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1271 wire1272/X vssd vssd vccd vccd _303_/B sky130_fd_sc_hd__buf_6
Xwire1282 wire1283/X vssd vssd vccd vccd _344_/B sky130_fd_sc_hd__buf_6
Xwire1293 wire1293/A vssd vssd vccd vccd wire1293/X sky130_fd_sc_hd__buf_6
XFILLER_19_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__466__C _466_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output787_A _543_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__371__A_N _499_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__482__B _482_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output954_A output954/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[12\] mprj_dat_i_user[12] wire1245/A vssd vssd vccd vccd wire1027/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_8_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__003__A _003_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[110\] la_data_out_core[110] _273_/X vssd vssd vccd vccd _093_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_27_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__376__C _376_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3676 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__392__B _392_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[9\]_A mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput202 la_iena_mprj[48] vssd vssd vccd vccd _211_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput213 la_iena_mprj[58] vssd vssd vccd vccd _221_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[9\]_A la_data_out_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput224 la_iena_mprj[68] vssd vssd vccd vccd _231_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_input149_A la_iena_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput235 la_iena_mprj[78] vssd vssd vccd vccd _241_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput246 la_iena_mprj[88] vssd vssd vccd vccd _251_/B sky130_fd_sc_hd__clkbuf_4
Xinput257 la_iena_mprj[98] vssd vssd vccd vccd _261_/B sky130_fd_sc_hd__clkbuf_4
Xinput268 la_oenb_mprj[107] vssd vssd vccd vccd _604_/A sky130_fd_sc_hd__clkbuf_4
Xinput279 la_oenb_mprj[117] vssd vssd vccd vccd _614_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__567__B _567_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input316_A la_oenb_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_583_ _583_/A _583_/B vssd vssd vccd vccd _583_/X sky130_fd_sc_hd__and2_4
XFILLER_44_544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__394__A_N _522_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__583__A _583_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput709 _074_/Y vssd vssd vccd vccd la_data_in_mprj[91] sky130_fd_sc_hd__buf_8
X_017_ _017_/A vssd vssd vccd vccd _017_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output535_A _373_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1166_A wire1167/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output702_A _068_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__477__B _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1333_A wire1333/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1090 _414_/X vssd vssd vccd vccd wire1090/X sky130_fd_sc_hd__buf_6
Xuser_to_mprj_in_gates\[47\] la_data_out_core[47] _210_/X vssd vssd vccd vccd _030_/A
+ sky130_fd_sc_hd__nand2_2
XANTENNA_wire1500_A wire1500/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[9\] la_data_out_core[9] _172_/X vssd vssd vccd vccd _156_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_25_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2080 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__387__B _387_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3440 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input266_A la_oenb_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input433_A mprj_dat_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__578__A _578_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__297__B _297_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_566_ _566_/A _566_/B vssd vssd vccd vccd _566_/X sky130_fd_sc_hd__and2_4
XFILLER_18_2536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_497_ _497_/A _497_/B vssd vssd vccd vccd _497_/X sky130_fd_sc_hd__and2_4
XFILLER_38_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output485_A _380_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput506 _392_/X vssd vssd vccd vccd la_data_in_core[23] sky130_fd_sc_hd__buf_8
Xoutput517 wire1102/X vssd vssd vccd vccd la_data_in_core[33] sky130_fd_sc_hd__buf_8
Xoutput528 wire1092/X vssd vssd vccd vccd la_data_in_core[43] sky130_fd_sc_hd__buf_8
XANTENNA_wire1283_A wire1283/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput539 wire1082/X vssd vssd vccd vccd la_data_in_core[53] sky130_fd_sc_hd__buf_8
XFILLER_46_3691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output917_A wire1148/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1450_A wire1451/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1548_A wire1548/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1715_A wire1715/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1036 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1378 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_104 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_115 _598_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 wire1685/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_420_ _548_/A _420_/B _420_/C vssd vssd vccd vccd _420_/X sky130_fd_sc_hd__and3b_4
XANTENNA_137 _207_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_148 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_159 _256_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_351_ _351_/A _351_/B vssd vssd vccd vccd _351_/X sky130_fd_sc_hd__and2_4
XFILLER_42_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_282_ _282_/A _282_/B vssd vssd vccd vccd _282_/X sky130_fd_sc_hd__and2_4
XFILLER_17_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__432__A_N _560_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input383_A la_oenb_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__580__B _580_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input77_A la_data_out_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__101__A _101_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_618_ _618_/A _618_/B vssd vssd vccd vccd _618_/X sky130_fd_sc_hd__and2_4
XTAP_3693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1031_A wire1031/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1129_A _360_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_549_ _549_/A _549_/B vssd vssd vccd vccd _549_/X sky130_fd_sc_hd__and2_4
XANTENNA__474__C _474_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output867_A wire1184/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1498_A wire1498/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__490__B _490_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1665_A wire1665/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__011__A _011_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3650 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[26\]_B wire1248/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__455__A_N _583_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__384__C _384_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput870 wire1224/X vssd vssd vccd vccd mprj_adr_o_user[2] sky130_fd_sc_hd__buf_8
Xoutput881 wire986/X vssd vssd vccd vccd mprj_dat_i_core[0] sky130_fd_sc_hd__buf_8
XFILLER_5_3644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput892 wire985/X vssd vssd vccd vccd mprj_dat_i_core[1] sky130_fd_sc_hd__buf_8
XFILLER_25_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1601 wire1601/A vssd vssd vccd vccd wire1601/X sky130_fd_sc_hd__buf_6
XFILLER_5_2943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1612 wire1612/A vssd vssd vccd vccd _584_/B sky130_fd_sc_hd__buf_6
Xwire1623 wire1623/A vssd vssd vccd vccd _572_/B sky130_fd_sc_hd__buf_6
Xwire1634 wire1634/A vssd vssd vccd vccd _513_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1645 wire1645/A vssd vssd vccd vccd _502_/B sky130_fd_sc_hd__buf_6
XFILLER_41_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1656 wire1657/X vssd vssd vccd vccd _494_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input131_A la_data_out_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_628 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1667 wire1667/A vssd vssd vccd vccd wire1667/X sky130_fd_sc_hd__buf_6
Xwire1678 wire1679/X vssd vssd vccd vccd _483_/B sky130_fd_sc_hd__buf_6
XANTENNA_input229_A la_iena_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1689 wire1690/X vssd vssd vccd vccd _477_/B sky130_fd_sc_hd__buf_6
XFILLER_19_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__575__B _575_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_403_ _531_/A _403_/B _403_/C vssd vssd vccd vccd _403_/X sky130_fd_sc_hd__and3b_2
XTAP_1532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_50 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_334_ _334_/A _334_/B vssd vssd vccd vccd _334_/X sky130_fd_sc_hd__and2_2
XTAP_1587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__591__A _591_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_265_ _265_/A _265_/B vssd vssd vccd vccd _265_/X sky130_fd_sc_hd__and2_2
XFILLER_31_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_196_ _196_/A _196_/B vssd vssd vccd vccd _196_/X sky130_fd_sc_hd__and2_2
XFILLER_13_2296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire964 _136_/Y vssd vssd vccd vccd wire964/X sky130_fd_sc_hd__buf_6
Xwire975 _125_/Y vssd vssd vccd vccd wire975/X sky130_fd_sc_hd__buf_6
XFILLER_41_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire986 _114_/Y vssd vssd vccd vccd wire986/X sky130_fd_sc_hd__buf_6
XFILLER_45_3915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire997 wire997/A vssd vssd vccd vccd _118_/A sky130_fd_sc_hd__buf_8
XFILLER_6_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1079_A _425_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_irq_gates\[2\]_A user_irq_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output615_A _104_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__478__A_N _606_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2486 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__485__B _485_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1413_A wire1414/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_15 _553_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_26 _198_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_37 _314_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_48 _375_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2330 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_59 _270_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__006__A _006_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2779 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__379__C _379_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__395__B _395_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3538 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_050_ _050_/A vssd vssd vccd vccd _050_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_30_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input179_A la_iena_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_4131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[50\]_A la_data_out_core[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input346_A la_oenb_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1420 wire1420/A vssd vssd vccd vccd wire1420/X sky130_fd_sc_hd__buf_6
XFILLER_21_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1431 wire1431/A vssd vssd vccd vccd _390_/B sky130_fd_sc_hd__buf_6
Xwire1442 wire1443/X vssd vssd vccd vccd _380_/B sky130_fd_sc_hd__buf_6
Xwire1453 wire1453/A vssd vssd vccd vccd wire1453/X sky130_fd_sc_hd__buf_6
XFILLER_4_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1464 wire1465/X vssd vssd vccd vccd _369_/B sky130_fd_sc_hd__buf_6
XANTENNA__586__A _586_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1475 wire1475/A vssd vssd vccd vccd wire1475/X sky130_fd_sc_hd__buf_6
XFILLER_1_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1486 wire1486/A vssd vssd vccd vccd _283_/A sky130_fd_sc_hd__buf_6
Xwire1497 wire1497/A vssd vssd vccd vccd _273_/A sky130_fd_sc_hd__buf_6
XFILLER_28_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_317_ _317_/A _317_/B vssd vssd vccd vccd _317_/X sky130_fd_sc_hd__and2_2
XFILLER_32_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput13 la_data_out_mprj[108] vssd vssd vccd vccd _477_/C sky130_fd_sc_hd__clkbuf_4
Xinput24 la_data_out_mprj[118] vssd vssd vccd vccd _487_/C sky130_fd_sc_hd__clkbuf_4
X_248_ _248_/A _248_/B vssd vssd vccd vccd _248_/X sky130_fd_sc_hd__and2_4
XFILLER_7_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput35 la_data_out_mprj[12] vssd vssd vccd vccd _381_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput46 la_data_out_mprj[22] vssd vssd vccd vccd _391_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_output565_A _446_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput57 la_data_out_mprj[32] vssd vssd vccd vccd _401_/C sky130_fd_sc_hd__clkbuf_4
Xinput68 la_data_out_mprj[42] vssd vssd vccd vccd _411_/C sky130_fd_sc_hd__clkbuf_4
Xinput79 la_data_out_mprj[52] vssd vssd vccd vccd _421_/C sky130_fd_sc_hd__clkbuf_4
X_179_ _179_/A _179_/B vssd vssd vccd vccd _179_/X sky130_fd_sc_hd__and2_1
XANTENNA_wire1196_A _326_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output732_A _608_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[41\]_A la_data_out_core[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1363_A wire1364/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[77\] la_data_out_core[77] _240_/X vssd vssd vccd vccd _060_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_38_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1530_A wire1530/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire983_A _117_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[32\]_A la_data_out_core[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput406 mprj_adr_o_core[26] vssd vssd vccd vccd wire1377/A sky130_fd_sc_hd__buf_6
Xinput417 mprj_adr_o_core[7] vssd vssd vccd vccd wire1351/A sky130_fd_sc_hd__buf_6
Xinput428 mprj_dat_o_core[16] vssd vssd vccd vccd wire1327/A sky130_fd_sc_hd__buf_6
XFILLER_40_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput439 mprj_dat_o_core[26] vssd vssd vccd vccd wire1305/A sky130_fd_sc_hd__buf_6
XFILLER_5_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[99\]_A la_data_out_core[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input296_A la_oenb_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_102_ _102_/A vssd vssd vccd vccd _102_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_33_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_033_ _033_/A vssd vssd vccd vccd _033_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[23\]_A la_data_out_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3282 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1250 _270_/X vssd vssd vccd vccd wire1250/X sky130_fd_sc_hd__buf_6
Xwire1261 _256_/X vssd vssd vccd vccd wire1261/X sky130_fd_sc_hd__buf_6
Xwire1272 wire1272/A vssd vssd vccd vccd wire1272/X sky130_fd_sc_hd__buf_6
Xwire1283 wire1283/A vssd vssd vccd vccd wire1283/X sky130_fd_sc_hd__buf_6
Xwire1294 wire1295/X vssd vssd vccd vccd _367_/B sky130_fd_sc_hd__buf_6
XFILLER_21_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output682_A _050_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__482__C _482_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1307 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output947_A wire1229/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1578_A wire1579/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[14\]_A la_data_out_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[103\] la_data_out_core[103] wire1254/X vssd vssd vccd vccd
+ _086_/A sky130_fd_sc_hd__nand2_4
XFILLER_26_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__392__C _392_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput203 la_iena_mprj[49] vssd vssd vccd vccd _212_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[9\]_B _172_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput214 la_iena_mprj[59] vssd vssd vccd vccd _222_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput225 la_iena_mprj[69] vssd vssd vccd vccd _232_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput236 la_iena_mprj[79] vssd vssd vccd vccd _242_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput247 la_iena_mprj[89] vssd vssd vccd vccd _252_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput258 la_iena_mprj[99] vssd vssd vccd vccd _262_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput269 la_oenb_mprj[108] vssd vssd vccd vccd _605_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_1071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input211_A la_iena_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_582_ _582_/A _582_/B vssd vssd vccd vccd _582_/X sky130_fd_sc_hd__and2_4
XFILLER_17_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input309_A la_oenb_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__583__B _583_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_2306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_016_ _016_/A vssd vssd vccd vccd _016_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_4023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3322 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__104__A _104_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2560 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output528_A wire1092/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1159_A _345_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__477__C _477_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1080 _424_/X vssd vssd vccd vccd wire1080/X sky130_fd_sc_hd__buf_6
Xwire1091 _413_/X vssd vssd vccd vccd wire1091/X sky130_fd_sc_hd__buf_6
XANTENNA_wire1326_A wire1327/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output897_A wire962/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__493__B _493_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__014__A _014_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__387__C _387_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input161_A la_iena_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input259_A la_iena_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__578__B _578_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input426_A mprj_dat_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input22_A la_data_out_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1322 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__594__A _594_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_565_ _565_/A _565_/B vssd vssd vccd vccd _565_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_496_ _624_/A _496_/B _496_/C vssd vssd vccd vccd _496_/X sky130_fd_sc_hd__and3b_1
XFILLER_35_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output478_A _482_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput507 _393_/X vssd vssd vccd vccd la_data_in_core[24] sky130_fd_sc_hd__buf_8
Xoutput518 wire1101/X vssd vssd vccd vccd la_data_in_core[34] sky130_fd_sc_hd__buf_8
XFILLER_29_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput529 wire1091/X vssd vssd vccd vccd la_data_in_core[44] sky130_fd_sc_hd__buf_8
XANTENNA_output645_A _016_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1276_A wire1276/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output812_A _566_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__488__B _488_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1610_A wire1610/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1708_A wire1708/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1048 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__009__A _009_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__384__A_N _512_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__398__B _398_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _589_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _197_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _207_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_149 _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ _350_/A _350_/B vssd vssd vccd vccd _350_/X sky130_fd_sc_hd__and2_4
XTAP_1758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_281_ _281_/A _281_/B vssd vssd vccd vccd _281_/X sky130_fd_sc_hd__and2_4
XFILLER_39_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input376_A la_oenb_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__589__A _589_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_617_ _617_/A _617_/B vssd vssd vccd vccd _617_/X sky130_fd_sc_hd__and2_4
XFILLER_37_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_548_ _548_/A _548_/B vssd vssd vccd vccd _548_/X sky130_fd_sc_hd__and2_4
XTAP_2982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1024_A wire1024/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output595_A _086_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_479_ _607_/A _479_/B _479_/C vssd vssd vccd vccd _479_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output762_A _520_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__490__C _490_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1393_A wire1393/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1560_A wire1561/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1658_A wire1659/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__499__A _499_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3422 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3190 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput860 wire1197/X vssd vssd vccd vccd mprj_adr_o_user[20] sky130_fd_sc_hd__buf_8
Xoutput871 wire1178/X vssd vssd vccd vccd mprj_adr_o_user[30] sky130_fd_sc_hd__buf_8
XFILLER_25_3551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput882 wire976/X vssd vssd vccd vccd mprj_dat_i_core[10] sky130_fd_sc_hd__buf_8
XFILLER_8_1311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput893 wire966/X vssd vssd vccd vccd mprj_dat_i_core[20] sky130_fd_sc_hd__buf_8
XANTENNA__202__A _202_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1602 wire1602/A vssd vssd vccd vccd _594_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1613 wire1613/A vssd vssd vccd vccd _583_/B sky130_fd_sc_hd__buf_6
Xwire1624 wire1624/A vssd vssd vccd vccd _569_/B sky130_fd_sc_hd__buf_6
XFILLER_25_2894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1635 wire1635/A vssd vssd vccd vccd _512_/B sky130_fd_sc_hd__buf_6
Xwire1646 wire1646/A vssd vssd vccd vccd _501_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1657 wire1657/A vssd vssd vccd vccd wire1657/X sky130_fd_sc_hd__buf_6
XFILLER_5_2999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1668 wire1669/X vssd vssd vccd vccd _488_/B sky130_fd_sc_hd__buf_6
Xwire1679 wire1679/A vssd vssd vccd vccd wire1679/X sky130_fd_sc_hd__buf_6
XFILLER_18_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input124_A la_data_out_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_684 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_402_ _530_/A _402_/B _402_/C vssd vssd vccd vccd _402_/X sky130_fd_sc_hd__and3b_2
XFILLER_19_2632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_333_ _333_/A _333_/B vssd vssd vccd vccd _333_/X sky130_fd_sc_hd__and2_2
XTAP_1577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__591__B _591_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_264_ _264_/A _264_/B vssd vssd vccd vccd _264_/X sky130_fd_sc_hd__and2_1
XFILLER_32_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_195_ _195_/A _195_/B vssd vssd vccd vccd _195_/X sky130_fd_sc_hd__and2_2
XFILLER_6_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire965 _135_/Y vssd vssd vccd vccd wire965/X sky130_fd_sc_hd__buf_6
XFILLER_26_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire976 _124_/Y vssd vssd vccd vccd wire976/X sky130_fd_sc_hd__buf_6
Xuser_wb_dat_gates\[5\] mprj_dat_i_user[5] rebuffer2/X vssd vssd vccd vccd wire996/A
+ sky130_fd_sc_hd__nand2_8
Xwire987 _085_/Y vssd vssd vccd vccd wire987/X sky130_fd_sc_hd__buf_6
Xwire998 wire998/A vssd vssd vccd vccd _117_/A sky130_fd_sc_hd__buf_8
XFILLER_26_3315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_irq_gates\[2\]_B _293_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output510_A wire1108/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output608_A _098_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1141_A _354_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1239_A wire1240/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__485__C _485_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1406_A wire1406/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[22\] la_data_out_core[22] _185_/X vssd vssd vccd vccd _005_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_36_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_16 _554_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_27 _201_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_38 _314_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_49 _375_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__422__A_N _550_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_938 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput690 _057_/Y vssd vssd vccd vccd la_data_in_mprj[74] sky130_fd_sc_hd__buf_8
XFILLER_40_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input241_A la_iena_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input339_A la_oenb_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1080 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1410 wire1411/X vssd vssd vccd vccd _318_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1421 wire1421/A vssd vssd vccd vccd _506_/A sky130_fd_sc_hd__buf_6
XFILLER_8_1174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1432 wire1432/A vssd vssd vccd vccd _389_/B sky130_fd_sc_hd__buf_6
XFILLER_46_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1443 wire1443/A vssd vssd vccd vccd wire1443/X sky130_fd_sc_hd__buf_6
XFILLER_5_2785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1454 wire1455/X vssd vssd vccd vccd _374_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1465 wire1465/A vssd vssd vccd vccd wire1465/X sky130_fd_sc_hd__buf_6
XFILLER_21_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1476 wire1476/A vssd vssd vccd vccd _290_/A sky130_fd_sc_hd__buf_6
XANTENNA__586__B _586_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1487 wire1488/X vssd vssd vccd vccd _282_/A sky130_fd_sc_hd__buf_6
Xwire1498 wire1498/A vssd vssd vccd vccd _272_/A sky130_fd_sc_hd__buf_6
XFILLER_46_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_316_ _316_/A _316_/B vssd vssd vccd vccd _316_/X sky130_fd_sc_hd__and2_4
XFILLER_30_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__107__A _107_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput14 la_data_out_mprj[109] vssd vssd vccd vccd _478_/C sky130_fd_sc_hd__clkbuf_4
X_247_ _247_/A _247_/B vssd vssd vccd vccd _247_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput25 la_data_out_mprj[119] vssd vssd vccd vccd _488_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_7_831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput36 la_data_out_mprj[13] vssd vssd vccd vccd _382_/C sky130_fd_sc_hd__clkbuf_4
Xinput47 la_data_out_mprj[23] vssd vssd vccd vccd _392_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_7_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput58 la_data_out_mprj[33] vssd vssd vccd vccd _402_/C sky130_fd_sc_hd__clkbuf_4
Xinput69 la_data_out_mprj[43] vssd vssd vccd vccd _412_/C sky130_fd_sc_hd__clkbuf_4
X_178_ _178_/A _178_/B vssd vssd vccd vccd _178_/X sky130_fd_sc_hd__and2_2
XFILLER_7_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output558_A wire1069/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1091_A _413_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__445__A_N _573_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output725_A _602_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__496__B _496_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire976_A _124_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__017__A _017_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[32\]_B _195_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput407 mprj_adr_o_core[27] vssd vssd vccd vccd wire1375/A sky130_fd_sc_hd__buf_6
Xinput418 mprj_adr_o_core[8] vssd vssd vccd vccd wire1348/A sky130_fd_sc_hd__buf_6
Xinput429 mprj_dat_o_core[17] vssd vssd vccd vccd wire1325/A sky130_fd_sc_hd__buf_6
XFILLER_22_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[99\]_B wire1258/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_996 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_101_ _101_/A vssd vssd vccd vccd _101_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_36_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input191_A la_iena_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input289_A la_oenb_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_032_ _032_/A vssd vssd vccd vccd _032_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__468__A_N _596_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input456_A mprj_sel_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input52_A la_data_out_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__597__A _597_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1240 _298_/X vssd vssd vccd vccd wire1240/X sky130_fd_sc_hd__buf_6
Xwire1251 _269_/X vssd vssd vccd vccd wire1251/X sky130_fd_sc_hd__buf_8
XFILLER_21_3086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1262 wire1262/A vssd vssd vccd vccd _293_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1273 wire1274/X vssd vssd vccd vccd _302_/B sky130_fd_sc_hd__buf_6
Xwire1284 wire1285/X vssd vssd vccd vccd _343_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1295 wire1295/A vssd vssd vccd vccd wire1295/X sky130_fd_sc_hd__buf_6
XFILLER_34_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_462 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output842_A _593_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1190 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1473_A wire1473/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1640_A wire1640/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1562 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__300__A _300_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3266 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput204 la_iena_mprj[4] vssd vssd vccd vccd _167_/B sky130_fd_sc_hd__clkbuf_4
Xinput215 la_iena_mprj[5] vssd vssd vccd vccd _168_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput226 la_iena_mprj[6] vssd vssd vccd vccd _169_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput237 la_iena_mprj[7] vssd vssd vccd vccd _170_/B sky130_fd_sc_hd__buf_4
XFILLER_2_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput248 la_iena_mprj[8] vssd vssd vccd vccd _171_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_2711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput259 la_iena_mprj[9] vssd vssd vccd vccd _172_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__210__A _210_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_581_ _581_/A _581_/B vssd vssd vccd vccd _581_/X sky130_fd_sc_hd__and2_4
XFILLER_38_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input204_A la_iena_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_015_ _015_/A vssd vssd vccd vccd _015_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_2826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__120__A _120_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1768 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1070 _437_/X vssd vssd vccd vccd wire1070/X sky130_fd_sc_hd__buf_6
Xwire1081 _423_/X vssd vssd vccd vccd wire1081/X sky130_fd_sc_hd__buf_6
Xwire1092 _412_/X vssd vssd vccd vccd wire1092/X sky130_fd_sc_hd__buf_6
XFILLER_21_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1221_A _310_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output792_A wire1051/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1319_A wire1319/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__493__C _493_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1590_A wire1590/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1688_A wire1688/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_992 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3682 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__205__A _205_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input154_A la_iena_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input321_A la_oenb_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input419_A mprj_adr_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1334 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input15_A la_data_out_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__594__B _594_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_564_ _564_/A _564_/B vssd vssd vccd vccd _564_/X sky130_fd_sc_hd__and2_4
XFILLER_17_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_495_ _623_/A _495_/B _495_/C vssd vssd vccd vccd _495_/X sky130_fd_sc_hd__and3b_1
XFILLER_31_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__115__A _115_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput508 _394_/X vssd vssd vccd vccd la_data_in_core[25] sky130_fd_sc_hd__buf_8
XFILLER_5_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput519 wire1100/X vssd vssd vccd vccd la_data_in_core[35] sky130_fd_sc_hd__buf_8
XFILLER_29_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output540_A wire1081/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output638_A _010_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3092 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1171_A _339_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1269_A wire1270/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_ack_gate mprj_ack_i_user max_cap1244/X vssd vssd vccd vccd wire1031/A sky130_fd_sc_hd__nand2_8
XFILLER_7_3197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__488__C _488_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output805_A _559_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1532 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1436_A wire1436/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[52\] la_data_out_core[52] _215_/X vssd vssd vccd vccd _035_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1603_A wire1603/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[29\]_A mprj_dat_i_user[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A la_data_out_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__398__C _398_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1643 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 _513_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_128 _197_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _213_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_280_ _280_/A _280_/B vssd vssd vccd vccd _280_/X sky130_fd_sc_hd__and2_4
XFILLER_13_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input271_A la_oenb_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input369_A la_oenb_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__589__B _589_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_616_ _616_/A _616_/B vssd vssd vccd vccd _616_/X sky130_fd_sc_hd__and2_2
XTAP_3673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_547_ _547_/A _547_/B vssd vssd vccd vccd _547_/X sky130_fd_sc_hd__and2_1
XTAP_2983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_478_ _606_/A _478_/B _478_/C vssd vssd vccd vccd _478_/X sky130_fd_sc_hd__and3b_4
XANTENNA_output490_A _493_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1017_A wire1018/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output588_A wire1060/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output755_A _514_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1386_A wire1387/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output922_A wire1138/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__499__B _499_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1553_A wire1553/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1720_A wire1720/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput850 wire1210/X vssd vssd vccd vccd mprj_adr_o_user[11] sky130_fd_sc_hd__buf_8
XFILLER_5_3602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput861 wire1196/X vssd vssd vccd vccd mprj_adr_o_user[21] sky130_fd_sc_hd__buf_8
XFILLER_21_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput872 wire1176/X vssd vssd vccd vccd mprj_adr_o_user[31] sky130_fd_sc_hd__buf_8
Xoutput883 wire975/X vssd vssd vccd vccd mprj_dat_i_core[11] sky130_fd_sc_hd__buf_8
XFILLER_25_3563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput894 wire965/X vssd vssd vccd vccd mprj_dat_i_core[21] sky130_fd_sc_hd__buf_8
XFILLER_5_2901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1603 wire1603/A vssd vssd vccd vccd _593_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1614 wire1614/A vssd vssd vccd vccd _582_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1625 wire1625/A vssd vssd vccd vccd _568_/B sky130_fd_sc_hd__buf_6
XTAP_390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1636 wire1636/A vssd vssd vccd vccd _511_/B sky130_fd_sc_hd__buf_6
XFILLER_46_405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1647 wire1647/A vssd vssd vccd vccd _500_/B sky130_fd_sc_hd__buf_6
XFILLER_41_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1658 wire1659/X vssd vssd vccd vccd _493_/B sky130_fd_sc_hd__buf_6
Xwire1669 wire1669/A vssd vssd vccd vccd wire1669/X sky130_fd_sc_hd__buf_6
XFILLER_46_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input117_A la_data_out_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_401_ _529_/A _401_/B _401_/C vssd vssd vccd vccd _401_/X sky130_fd_sc_hd__and3b_2
XTAP_2257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_332_ _332_/A _332_/B vssd vssd vccd vccd _332_/X sky130_fd_sc_hd__and2_2
XTAP_1578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_263_ _263_/A _263_/B vssd vssd vccd vccd _263_/X sky130_fd_sc_hd__and2_2
XFILLER_6_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input82_A la_data_out_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_194_ _194_/A _194_/B vssd vssd vccd vccd _194_/X sky130_fd_sc_hd__and2_2
Xwire966 _134_/Y vssd vssd vccd vccd wire966/X sky130_fd_sc_hd__buf_6
Xwire977 _123_/Y vssd vssd vccd vccd wire977/X sky130_fd_sc_hd__buf_6
XFILLER_6_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire988 _084_/Y vssd vssd vccd vccd wire988/X sky130_fd_sc_hd__buf_6
XFILLER_30_2590 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire999 wire999/A vssd vssd vccd vccd _145_/A sky130_fd_sc_hd__buf_6
XFILLER_6_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output503_A _389_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1134_A wire1135/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__374__A_N _502_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_828 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output872_A wire1176/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_17 _554_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_28 _201_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[15\] la_data_out_core[15] _178_/X vssd vssd vccd vccd _162_/A
+ sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_gates\[28\] mprj_dat_i_user[28] split13/X vssd vssd vccd vccd wire1004/A
+ sky130_fd_sc_hd__nand2_2
XANTENNA_39 _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1670_A wire1671/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__303__A _303_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[126\] la_data_out_core[126] _289_/X vssd vssd vccd vccd _109_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_25_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_rebuffer5_A split13/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__213__A _213_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput680 _048_/Y vssd vssd vccd vccd la_data_in_mprj[65] sky130_fd_sc_hd__buf_8
Xoutput691 _058_/Y vssd vssd vccd vccd la_data_in_mprj[75] sky130_fd_sc_hd__buf_8
XFILLER_43_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3476 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1400 wire1400/A vssd vssd vccd vccd wire1400/X sky130_fd_sc_hd__buf_6
XFILLER_21_2501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1411 wire1412/X vssd vssd vccd vccd wire1411/X sky130_fd_sc_hd__buf_6
Xwire1422 wire1422/A vssd vssd vccd vccd _502_/A sky130_fd_sc_hd__buf_6
XANTENNA_input234_A la_iena_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1433 wire1433/A vssd vssd vccd vccd _388_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1444 wire1445/X vssd vssd vccd vccd _379_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1455 wire1455/A vssd vssd vccd vccd wire1455/X sky130_fd_sc_hd__buf_6
Xwire1466 wire1466/A vssd vssd vccd vccd _294_/A sky130_fd_sc_hd__buf_6
Xwire1477 wire1478/X vssd vssd vccd vccd _289_/A sky130_fd_sc_hd__buf_6
XFILLER_1_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__397__A_N _525_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1488 wire1488/A vssd vssd vccd vccd wire1488/X sky130_fd_sc_hd__buf_6
XFILLER_35_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1499 wire1499/A vssd vssd vccd vccd _271_/A sky130_fd_sc_hd__buf_6
XFILLER_46_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input401_A mprj_adr_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_315_ _315_/A _315_/B vssd vssd vccd vccd _315_/X sky130_fd_sc_hd__and2_2
XTAP_1397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_246_ _246_/A _246_/B vssd vssd vccd vccd _246_/X sky130_fd_sc_hd__and2_4
XFILLER_7_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput15 la_data_out_mprj[10] vssd vssd vccd vccd _379_/C sky130_fd_sc_hd__clkbuf_4
Xinput26 la_data_out_mprj[11] vssd vssd vccd vccd _380_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_32_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput37 la_data_out_mprj[14] vssd vssd vccd vccd _383_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_32_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput48 la_data_out_mprj[24] vssd vssd vccd vccd _393_/C sky130_fd_sc_hd__clkbuf_4
Xinput59 la_data_out_mprj[34] vssd vssd vccd vccd _403_/C sky130_fd_sc_hd__clkbuf_4
X_177_ _177_/A _177_/B vssd vssd vccd vccd _177_/X sky130_fd_sc_hd__and2_2
XFILLER_26_3102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__123__A _123_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1084_A _420_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output620_A _109_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1349_A wire1350/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__496__C _496_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1354 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire969_A _131_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__033__A _033_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput408 mprj_adr_o_core[28] vssd vssd vccd vccd wire1373/A sky130_fd_sc_hd__buf_6
XFILLER_44_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput419 mprj_adr_o_core[9] vssd vssd vccd vccd wire1345/A sky130_fd_sc_hd__buf_6
XFILLER_6_3785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__208__A _208_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_100_ _100_/A vssd vssd vccd vccd _100_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_031_ _031_/A vssd vssd vccd vccd _031_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input184_A la_iena_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input351_A la_oenb_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input449_A mprj_dat_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input45_A la_data_out_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__597__B _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1230 _303_/X vssd vssd vccd vccd wire1230/X sky130_fd_sc_hd__buf_6
Xwire1241 _297_/X vssd vssd vccd vccd wire1241/X sky130_fd_sc_hd__buf_6
XFILLER_40_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1252 _268_/X vssd vssd vccd vccd wire1252/X sky130_fd_sc_hd__buf_6
XFILLER_5_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1263 wire1263/A vssd vssd vccd vccd _292_/B sky130_fd_sc_hd__buf_6
Xwire1274 wire1274/A vssd vssd vccd vccd wire1274/X sky130_fd_sc_hd__buf_6
Xwire1285 wire1285/A vssd vssd vccd vccd wire1285/X sky130_fd_sc_hd__buf_6
XFILLER_1_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1296 wire1297/X vssd vssd vccd vccd _339_/B sky130_fd_sc_hd__buf_6
XFILLER_1_1746 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__118__A _118_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__412__A_N _540_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output570_A _450_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_229_ _229_/A _229_/B vssd vssd vccd vccd _229_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1299_A wire1299/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_684 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output835_A _505_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1466_A wire1466/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[82\] la_data_out_core[82] _245_/X vssd vssd vccd vccd _065_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_6_3059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2887 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__300__B _300_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__028__A _028_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3278 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput205 la_iena_mprj[50] vssd vssd vccd vccd _213_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput216 la_iena_mprj[60] vssd vssd vccd vccd _223_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput227 la_iena_mprj[70] vssd vssd vccd vccd _233_/B sky130_fd_sc_hd__clkbuf_4
Xinput238 la_iena_mprj[80] vssd vssd vccd vccd _243_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput249 la_iena_mprj[90] vssd vssd vccd vccd _253_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__210__B _210_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_580_ _580_/A _580_/B vssd vssd vccd vccd _580_/X sky130_fd_sc_hd__and2_4
XFILLER_44_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__435__A_N _563_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input399_A mprj_adr_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_014_ _014_/A vssd vssd vccd vccd _014_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_3831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1060 _467_/X vssd vssd vccd vccd wire1060/X sky130_fd_sc_hd__buf_6
XFILLER_1_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1071 _434_/X vssd vssd vccd vccd wire1071/X sky130_fd_sc_hd__buf_6
Xwire1082 _422_/X vssd vssd vccd vccd wire1082/X sky130_fd_sc_hd__buf_6
XFILLER_35_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1093 _411_/X vssd vssd vccd vccd wire1093/X sky130_fd_sc_hd__buf_6
XFILLER_21_1471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output785_A _541_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output952_A output952/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[10\] mprj_dat_i_user[10] rebuffer10/X vssd vssd vccd vccd wire1029/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_11_1106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1583_A wire1583/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__311__A _311_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__458__A_N _586_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_908 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__221__A _221_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input147_A la_iena_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1346 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input314_A la_oenb_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_563_ _563_/A _563_/B vssd vssd vccd vccd _563_/X sky130_fd_sc_hd__and2_4
XFILLER_2_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_494_ _622_/A _494_/B _494_/C vssd vssd vccd vccd _494_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput509 wire1109/X vssd vssd vccd vccd la_data_in_core[26] sky130_fd_sc_hd__buf_8
XFILLER_10_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output533_A wire1087/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__131__A _131_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2234 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1164_A wire1165/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_2267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output700_A _066_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1331_A wire1331/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1429_A wire1429/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[45\] la_data_out_core[45] _208_/X vssd vssd vccd vccd _028_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_39_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__306__A _306_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[7\] la_data_out_core[7] _170_/X vssd vssd vccd vccd _154_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_25_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3839 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__041__A _041_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[29\]_B wire1248/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_107 _613_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 la_iena_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _197_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__216__A _216_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[80\]_A la_data_out_core[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input264_A la_oenb_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3474 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input431_A mprj_dat_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_615_ _615_/A _615_/B vssd vssd vccd vccd _615_/X sky130_fd_sc_hd__and2_1
XTAP_3663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_546_ _546_/A _546_/B vssd vssd vccd vccd _546_/X sky130_fd_sc_hd__and2_4
XTAP_2962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_477_ _605_/A _477_/B _477_/C vssd vssd vccd vccd _477_/X sky130_fd_sc_hd__and3b_4
XFILLER_38_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output483_A _487_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__126__A _126_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output650_A _021_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[71\]_A la_data_out_core[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output748_A wire1033/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1281_A wire1281/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1379_A wire1379/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output915_A wire1152/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1546_A wire1546/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1713_A wire1713/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire999_A wire999/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__036__A _036_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[62\]_A la_data_out_core[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput840 _591_/X vssd vssd vccd vccd la_oenb_core[94] sky130_fd_sc_hd__buf_8
XFILLER_43_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput851 wire1208/X vssd vssd vccd vccd mprj_adr_o_user[12] sky130_fd_sc_hd__buf_8
Xoutput862 wire1194/X vssd vssd vccd vccd mprj_adr_o_user[22] sky130_fd_sc_hd__buf_8
XFILLER_5_3614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput873 wire1223/X vssd vssd vccd vccd mprj_adr_o_user[3] sky130_fd_sc_hd__buf_8
Xoutput884 wire974/X vssd vssd vccd vccd mprj_dat_i_core[12] sky130_fd_sc_hd__buf_8
XFILLER_25_3575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput895 wire964/X vssd vssd vccd vccd mprj_dat_i_core[22] sky130_fd_sc_hd__buf_8
XFILLER_25_2841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1604 wire1604/A vssd vssd vccd vccd _592_/B sky130_fd_sc_hd__buf_6
XFILLER_28_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1615 wire1615/A vssd vssd vccd vccd _581_/B sky130_fd_sc_hd__buf_6
XFILLER_41_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1626 wire1626/A vssd vssd vccd vccd _566_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1637 wire1637/A vssd vssd vccd vccd _510_/B sky130_fd_sc_hd__buf_6
XTAP_391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1648 wire1648/A vssd vssd vccd vccd _499_/B sky130_fd_sc_hd__buf_6
XFILLER_3_3393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1659 wire1659/A vssd vssd vccd vccd wire1659/X sky130_fd_sc_hd__buf_6
XFILLER_41_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_400_ _528_/A _400_/B _400_/C vssd vssd vccd vccd _400_/X sky130_fd_sc_hd__and3b_2
XTAP_1502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_331_ _331_/A _331_/B vssd vssd vccd vccd _331_/X sky130_fd_sc_hd__and2_2
XFILLER_32_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_262_ _262_/A _262_/B vssd vssd vccd vccd _262_/X sky130_fd_sc_hd__and2_2
XFILLER_23_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input381_A la_oenb_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_193_ _193_/A _193_/B vssd vssd vccd vccd _193_/X sky130_fd_sc_hd__and2_2
XFILLER_6_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire967 _133_/Y vssd vssd vccd vccd wire967/X sky130_fd_sc_hd__buf_6
Xwire978 _122_/Y vssd vssd vccd vccd wire978/X sky130_fd_sc_hd__buf_6
XANTENNA_input75_A la_data_out_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire989 _083_/Y vssd vssd vccd vccd wire989/X sky130_fd_sc_hd__buf_6
XFILLER_6_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[53\]_A la_data_out_core[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1127_A _361_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output698_A _064_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_529_ _529_/A _529_/B vssd vssd vccd vccd _529_/X sky130_fd_sc_hd__and2_4
XTAP_2792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_18 _196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_29 _201_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output865_A wire1188/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1496_A wire1496/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[44\]_A la_data_out_core[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1663_A wire1663/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__303__B _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3923 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1550 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[119\] la_data_out_core[119] _282_/X vssd vssd vccd vccd _102_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_0_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[35\]_A la_data_out_core[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__213__B _213_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput670 _039_/Y vssd vssd vccd vccd la_data_in_mprj[56] sky130_fd_sc_hd__buf_8
Xoutput681 _049_/Y vssd vssd vccd vccd la_data_in_mprj[66] sky130_fd_sc_hd__buf_8
XFILLER_27_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput692 _059_/Y vssd vssd vccd vccd la_data_in_mprj[76] sky130_fd_sc_hd__buf_8
XFILLER_40_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1401 wire1402/X vssd vssd vccd vccd _321_/B sky130_fd_sc_hd__buf_6
Xwire1412 wire1412/A vssd vssd vccd vccd wire1412/X sky130_fd_sc_hd__buf_6
XFILLER_28_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1423 input3/X vssd vssd vccd vccd _295_/A_N sky130_fd_sc_hd__buf_6
XFILLER_43_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1434 wire1434/A vssd vssd vccd vccd _387_/B sky130_fd_sc_hd__buf_6
XFILLER_4_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1445 wire1445/A vssd vssd vccd vccd wire1445/X sky130_fd_sc_hd__buf_6
Xwire1456 wire1457/X vssd vssd vccd vccd _373_/B sky130_fd_sc_hd__buf_6
Xwire1467 wire1468/X vssd vssd vccd vccd wire1467/X sky130_fd_sc_hd__buf_6
XFILLER_46_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input227_A la_iena_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1478 wire1478/A vssd vssd vccd vccd wire1478/X sky130_fd_sc_hd__buf_6
Xwire1489 wire1489/A vssd vssd vccd vccd _281_/A sky130_fd_sc_hd__buf_6
XTAP_2000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_314_ _314_/A _314_/B vssd vssd vccd vccd _314_/X sky130_fd_sc_hd__and2_2
XFILLER_12_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_800 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_245_ _245_/A _245_/B vssd vssd vccd vccd _245_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput16 la_data_out_mprj[110] vssd vssd vccd vccd _479_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_32_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput27 la_data_out_mprj[120] vssd vssd vccd vccd _489_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_35_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput38 la_data_out_mprj[15] vssd vssd vccd vccd _384_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_6_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_176_ _176_/A _176_/B vssd vssd vccd vccd _176_/X sky130_fd_sc_hd__and2_4
Xinput49 la_data_out_mprj[25] vssd vssd vccd vccd _394_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_gates\[26\]_A la_data_out_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[110\]_A la_data_out_core[110] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_13_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2446 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1077_A _427_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1411_A wire1412/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__491__A_N _619_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1509_A wire1509/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1716 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[17\]_A la_data_out_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_A la_data_out_core[101] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_6_3731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2092 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput409 mprj_adr_o_core[29] vssd vssd vccd vccd wire1371/A sky130_fd_sc_hd__buf_6
XFILLER_44_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_030_ _030_/A vssd vssd vccd vccd _030_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input177_A la_iena_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input344_A la_oenb_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input38_A la_data_out_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1220 _311_/X vssd vssd vccd vccd wire1220/X sky130_fd_sc_hd__buf_6
XFILLER_21_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1231 wire1232/X vssd vssd vccd vccd wire1231/X sky130_fd_sc_hd__buf_6
Xwire1242 _296_/X vssd vssd vccd vccd wire1242/X sky130_fd_sc_hd__buf_6
Xwire1253 _267_/X vssd vssd vccd vccd wire1253/X sky130_fd_sc_hd__buf_6
XFILLER_19_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1264 wire1264/A vssd vssd vccd vccd _291_/B sky130_fd_sc_hd__buf_4
Xwire1275 wire1276/X vssd vssd vccd vccd _301_/B sky130_fd_sc_hd__buf_6
Xwire1286 wire1287/X vssd vssd vccd vccd _342_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1297 wire1297/A vssd vssd vccd vccd wire1297/X sky130_fd_sc_hd__buf_6
XFILLER_21_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_228_ _228_/A _228_/B vssd vssd vccd vccd _228_/X sky130_fd_sc_hd__and2_4
XFILLER_7_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output563_A _444_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__134__A _134_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_159_ _159_/A vssd vssd vccd vccd _159_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_3523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1194_A wire1195/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output730_A _507_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output828_A _580_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1361_A wire1362/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1459_A wire1459/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[75\] la_data_out_core[75] _238_/X vssd vssd vccd vccd _058_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire981_A _119_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_3393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__044__A _044_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__387__A_N _515_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput206 la_iena_mprj[51] vssd vssd vccd vccd _214_/B sky130_fd_sc_hd__clkbuf_4
Xinput217 la_iena_mprj[61] vssd vssd vccd vccd _224_/B sky130_fd_sc_hd__clkbuf_4
Xinput228 la_iena_mprj[71] vssd vssd vccd vccd _234_/B sky130_fd_sc_hd__buf_4
XFILLER_44_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput239 la_iena_mprj[81] vssd vssd vccd vccd _244_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__219__A _219_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input294_A la_oenb_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_013_ _013_/A vssd vssd vccd vccd _013_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1078 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input461_A user_irq_ena[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__401__B _401_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1050 _553_/X vssd vssd vccd vccd wire1050/X sky130_fd_sc_hd__buf_6
XFILLER_1_2223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1061 _466_/X vssd vssd vccd vccd wire1061/X sky130_fd_sc_hd__buf_6
XFILLER_40_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1072 _433_/X vssd vssd vccd vccd wire1072/X sky130_fd_sc_hd__buf_6
XFILLER_38_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1083 _421_/X vssd vssd vccd vccd wire1083/X sky130_fd_sc_hd__buf_6
Xwire1094 _410_/X vssd vssd vccd vccd wire1094/X sky130_fd_sc_hd__buf_6
XFILLER_21_1461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__129__A _129_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_710 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1207_A _318_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1800 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output778_A _535_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output945_A wire1233/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_482 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1576_A wire1577/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__311__B _311_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[101\] la_data_out_core[101] wire1256/X vssd vssd vccd vccd
+ _084_/A sky130_fd_sc_hd__nand2_2
XFILLER_17_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__039__A _039_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__502__A _502_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__221__B _221_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__402__A_N _530_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1358 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_562_ _562_/A _562_/B vssd vssd vccd vccd _562_/X sky130_fd_sc_hd__and2_4
XANTENNA_input307_A la_oenb_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_493_ _621_/A _493_/B _493_/C vssd vssd vccd vccd _493_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_931 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output526_A wire1094/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1157_A _346_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1324_A wire1325/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output895_A wire964/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[38\] la_data_out_core[38] _201_/X vssd vssd vccd vccd _021_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_36_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1693_A wire1693/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3374 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__306__B _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__322__A _322_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__425__A_N _553_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_108 _613_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_119 mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1438 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__216__B _216_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1162 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[80\]_B _243_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__232__A _232_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3464 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input257_A la_iena_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3486 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input424_A mprj_dat_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input20_A la_data_out_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_614_ _614_/A _614_/B vssd vssd vccd vccd _614_/X sky130_fd_sc_hd__and2_4
XTAP_3653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_545_ _545_/A _545_/B vssd vssd vccd vccd _545_/X sky130_fd_sc_hd__and2_4
XFILLER_33_827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_2348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_476_ _604_/A _476_/B _476_/C vssd vssd vccd vccd _476_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output476_A _480_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[71\]_B _234_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__448__A_N _576_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output643_A _014_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__142__A _142_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1274_A wire1274/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output810_A _564_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output908_A wire981/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1539_A wire1539/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1706_A wire1706/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[62\]_B _225_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput830 _582_/X vssd vssd vccd vccd la_oenb_core[85] sky130_fd_sc_hd__buf_8
XANTENNA__052__A _052_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput841 wire1047/X vssd vssd vccd vccd la_oenb_core[95] sky130_fd_sc_hd__buf_8
Xoutput852 wire1207/X vssd vssd vccd vccd mprj_adr_o_user[13] sky130_fd_sc_hd__buf_8
Xoutput863 wire1192/X vssd vssd vccd vccd mprj_adr_o_user[23] sky130_fd_sc_hd__buf_8
Xoutput874 wire1222/X vssd vssd vccd vccd mprj_adr_o_user[4] sky130_fd_sc_hd__buf_8
Xoutput885 wire973/X vssd vssd vccd vccd mprj_dat_i_core[13] sky130_fd_sc_hd__buf_8
Xoutput896 wire963/X vssd vssd vccd vccd mprj_dat_i_core[23] sky130_fd_sc_hd__buf_8
XFILLER_5_2914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1605 wire1605/A vssd vssd vccd vccd _591_/B sky130_fd_sc_hd__buf_6
Xwire1616 wire1616/A vssd vssd vccd vccd _580_/B sky130_fd_sc_hd__buf_6
XTAP_370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1627 wire1627/A vssd vssd vccd vccd _528_/B sky130_fd_sc_hd__buf_6
XFILLER_41_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1638 wire1638/A vssd vssd vccd vccd _509_/B sky130_fd_sc_hd__buf_4
XFILLER_3_3372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1649 wire1649/A vssd vssd vccd vccd _498_/B sky130_fd_sc_hd__buf_6
XFILLER_19_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_643 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_43 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_330_ _330_/A _330_/B vssd vssd vccd vccd _330_/X sky130_fd_sc_hd__and2_1
XFILLER_26_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__227__A _227_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_261_ _261_/A _261_/B vssd vssd vccd vccd _261_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_192_ _192_/A _192_/B vssd vssd vccd vccd _192_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire968 _132_/Y vssd vssd vccd vccd wire968/X sky130_fd_sc_hd__buf_6
Xwire979 _121_/Y vssd vssd vccd vccd wire979/X sky130_fd_sc_hd__buf_6
XANTENNA_input374_A la_oenb_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input68_A la_data_out_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_528_ _528_/A _528_/B vssd vssd vccd vccd _528_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1022_A wire1022/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output593_A wire988/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__137__A _137_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_19 _196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_459_ _587_/A _459_/B _459_/C vssd vssd vccd vccd _459_/X sky130_fd_sc_hd__and3b_2
XFILLER_32_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output760_A _518_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output858_A wire1199/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1391_A wire1392/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1489_A wire1489/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1656_A wire1657/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__600__A _600_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__047__A _047_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1110 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput660 _030_/Y vssd vssd vccd vccd la_data_in_mprj[47] sky130_fd_sc_hd__buf_8
XFILLER_40_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput671 _040_/Y vssd vssd vccd vccd la_data_in_mprj[57] sky130_fd_sc_hd__buf_8
Xoutput682 _050_/Y vssd vssd vccd vccd la_data_in_mprj[67] sky130_fd_sc_hd__buf_8
XFILLER_21_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput693 _060_/Y vssd vssd vccd vccd la_data_in_mprj[77] sky130_fd_sc_hd__buf_8
XFILLER_8_1111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__510__A _510_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1402 wire1403/X vssd vssd vccd vccd wire1402/X sky130_fd_sc_hd__buf_6
XFILLER_8_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1413 wire1414/X vssd vssd vccd vccd _317_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1424 wire1424/A vssd vssd vccd vccd _498_/A sky130_fd_sc_hd__buf_6
XFILLER_5_2766 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1435 wire1435/A vssd vssd vccd vccd _386_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1446 wire1447/X vssd vssd vccd vccd _378_/B sky130_fd_sc_hd__buf_6
Xwire1457 wire1457/A vssd vssd vccd vccd wire1457/X sky130_fd_sc_hd__buf_6
Xwire1468 wire1469/X vssd vssd vccd vccd wire1468/X sky130_fd_sc_hd__buf_6
XFILLER_46_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1479 wire1480/X vssd vssd vccd vccd _288_/A sky130_fd_sc_hd__buf_6
XFILLER_38_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input122_A la_data_out_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_313_ _313_/A _313_/B vssd vssd vccd vccd _313_/X sky130_fd_sc_hd__and2_4
XTAP_1388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_244_ _244_/A _244_/B vssd vssd vccd vccd _244_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput17 la_data_out_mprj[111] vssd vssd vccd vccd _480_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput28 la_data_out_mprj[121] vssd vssd vccd vccd _490_/C sky130_fd_sc_hd__clkbuf_4
Xinput39 la_data_out_mprj[16] vssd vssd vccd vccd _385_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_175_ _175_/A _175_/B vssd vssd vccd vccd _175_/X sky130_fd_sc_hd__and2_4
XFILLER_6_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[3\] mprj_dat_i_user[3] max_cap1244/X vssd vssd vccd vccd wire998/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_7_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__404__B _404_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[110\]_B _273_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3727 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2458 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output606_A _096_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1237_A wire1238/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1404_A wire1405/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[20\] la_data_out_core[20] _183_/X vssd vssd vccd vccd _003_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_15_3564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__314__B _314_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_B wire1256/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3743 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__330__A _330_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[10\]_A mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__505__A _505_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__224__B _224_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__240__A _240_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput490 _493_/X vssd vssd vccd vccd la_data_in_core[124] sky130_fd_sc_hd__buf_8
XFILLER_43_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input337_A la_oenb_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1210 wire1211/X vssd vssd vccd vccd wire1210/X sky130_fd_sc_hd__buf_6
XFILLER_43_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1221 _310_/X vssd vssd vccd vccd wire1221/X sky130_fd_sc_hd__buf_6
Xwire1232 _302_/X vssd vssd vccd vccd wire1232/X sky130_fd_sc_hd__buf_6
Xwire1243 _295_/X vssd vssd vccd vccd wire1243/X sky130_fd_sc_hd__buf_6
Xwire1254 _266_/X vssd vssd vccd vccd wire1254/X sky130_fd_sc_hd__buf_6
XFILLER_19_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1265 wire1266/X vssd vssd vccd vccd _300_/B sky130_fd_sc_hd__buf_6
XFILLER_25_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1276 wire1276/A vssd vssd vccd vccd wire1276/X sky130_fd_sc_hd__buf_6
XFILLER_1_2449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1287 wire1287/A vssd vssd vccd vccd wire1287/X sky130_fd_sc_hd__buf_6
Xwire1298 wire1299/X vssd vssd vccd vccd _366_/B sky130_fd_sc_hd__buf_6
XFILLER_34_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_227_ _227_/A _227_/B vssd vssd vccd vccd _227_/X sky130_fd_sc_hd__and2_4
XFILLER_6_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_158_ _158_/A vssd vssd vccd vccd _158_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_13_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1794 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output556_A _438_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_089_ _089_/A vssd vssd vccd vccd _089_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_3579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output723_A wire1044/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__150__A _150_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1354_A wire1355/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[68\] la_data_out_core[68] _231_/X vssd vssd vccd vccd _051_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_22_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1619_A wire1619/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__309__B _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire974_A _126_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__325__A _325_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__060__A _060_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput207 la_iena_mprj[52] vssd vssd vccd vccd _215_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput218 la_iena_mprj[62] vssd vssd vccd vccd _225_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_41_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput229 la_iena_mprj[72] vssd vssd vccd vccd _235_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__219__B _219_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__235__A _235_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input287_A la_oenb_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_012_ _012_/A vssd vssd vccd vccd _012_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input454_A mprj_sel_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input50_A la_data_out_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__481__A_N _609_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__401__C _401_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1040 _613_/X vssd vssd vccd vccd wire1040/X sky130_fd_sc_hd__buf_6
Xwire1051 _547_/X vssd vssd vccd vccd wire1051/X sky130_fd_sc_hd__buf_6
Xwire1062 _464_/X vssd vssd vccd vccd wire1062/X sky130_fd_sc_hd__buf_6
Xwire1073 _431_/X vssd vssd vccd vccd wire1073/X sky130_fd_sc_hd__buf_6
XFILLER_35_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1084 _420_/X vssd vssd vccd vccd wire1084/X sky130_fd_sc_hd__buf_6
XFILLER_40_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1095 _409_/X vssd vssd vccd vccd wire1095/X sky130_fd_sc_hd__buf_6
XFILLER_1_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1856 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__145__A _145_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output840_A _591_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output938_A wire1168/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1569_A wire1569/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__055__A _055_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__502__B _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_561_ _561_/A _561_/B vssd vssd vccd vccd _561_/X sky130_fd_sc_hd__and2_4
XFILLER_2_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input202_A la_iena_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_492_ _620_/A _492_/B _492_/C vssd vssd vccd vccd _492_/X sky130_fd_sc_hd__and3b_4
XFILLER_44_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input98_A la_data_out_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__412__B _412_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output519_A wire1100/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__377__A_N _505_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output790_A _546_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1317_A wire1317/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_880 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output888_A wire970/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1686_A wire1686/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__603__A _603_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__322__B _322_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[2\]_A mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1446 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 _613_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[2\]_A la_data_out_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__513__A _513_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__232__B _232_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input152_A la_iena_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input417_A mprj_adr_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_613_ _613_/A _613_/B vssd vssd vccd vccd _613_/X sky130_fd_sc_hd__and2_2
XTAP_3643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input13_A la_data_out_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_544_ _544_/A _544_/B vssd vssd vccd vccd _544_/X sky130_fd_sc_hd__and2_4
XTAP_2942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_475_ _603_/A _475_/B _475_/C vssd vssd vccd vccd _475_/X sky130_fd_sc_hd__and3b_4
XTAP_2997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__407__B _407_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1940 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output469_A wire1056/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output636_A _008_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1267_A wire1268/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output803_A wire1048/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1434_A wire1434/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput390 mprj_adr_o_core[11] vssd vssd vccd vccd wire1416/A sky130_fd_sc_hd__buf_6
Xuser_to_mprj_in_gates\[50\] la_data_out_core[50] _213_/X vssd vssd vccd vccd _033_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_3_1448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__317__B _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__333__A _333_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput820 _573_/X vssd vssd vccd vccd la_oenb_core[76] sky130_fd_sc_hd__buf_8
Xoutput831 _583_/X vssd vssd vccd vccd la_oenb_core[86] sky130_fd_sc_hd__buf_8
XFILLER_9_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput842 _593_/X vssd vssd vccd vccd la_oenb_core[96] sky130_fd_sc_hd__buf_8
Xoutput853 wire1206/X vssd vssd vccd vccd mprj_adr_o_user[14] sky130_fd_sc_hd__buf_8
XFILLER_25_3533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput864 wire1190/X vssd vssd vccd vccd mprj_adr_o_user[24] sky130_fd_sc_hd__buf_8
Xoutput875 wire1221/X vssd vssd vccd vccd mprj_adr_o_user[5] sky130_fd_sc_hd__buf_8
XFILLER_8_1304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput886 wire972/X vssd vssd vccd vccd mprj_dat_i_core[14] sky130_fd_sc_hd__buf_8
Xoutput897 wire962/X vssd vssd vccd vccd mprj_dat_i_core[24] sky130_fd_sc_hd__buf_8
XFILLER_25_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input5_A la_data_out_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1606 wire1606/A vssd vssd vccd vccd _590_/B sky130_fd_sc_hd__buf_6
XTAP_371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1617 wire1617/A vssd vssd vccd vccd _579_/B sky130_fd_sc_hd__buf_6
Xwire1628 wire1628/A vssd vssd vccd vccd _524_/B sky130_fd_sc_hd__buf_6
XTAP_382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1639 wire1639/A vssd vssd vccd vccd _508_/B sky130_fd_sc_hd__buf_6
XTAP_393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__508__A _508_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_260_ _260_/A _260_/B vssd vssd vccd vccd _260_/X sky130_fd_sc_hd__and2_4
XANTENNA__227__B _227_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_191_ _191_/A _191_/B vssd vssd vccd vccd _191_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire969 _131_/Y vssd vssd vccd vccd wire969/X sky130_fd_sc_hd__buf_6
XANTENNA__243__A _243_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input367_A la_oenb_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_irq_gates\[2\] user_irq_core[2] _293_/X vssd vssd vccd vccd _113_/A sky130_fd_sc_hd__nand2_2
XFILLER_43_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_527_ _527_/A _527_/B vssd vssd vccd vccd _527_/X sky130_fd_sc_hd__and2_4
XTAP_2772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_458_ _586_/A _458_/B _458_/C vssd vssd vccd vccd _458_/X sky130_fd_sc_hd__and3b_2
XANTENNA__415__A_N _543_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1015_A wire1016/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output586_A _465_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_389_ _517_/A _389_/B _389_/C vssd vssd vccd vccd _389_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_1601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output753_A _512_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1384_A wire1385/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output920_A wire1142/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[98\] la_data_out_core[98] _261_/X vssd vssd vccd vccd _081_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_42_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1551_A wire1551/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1649_A wire1649/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__600__B _600_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__328__A _328_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1122 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__063__A _063_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput650 _021_/Y vssd vssd vccd vccd la_data_in_mprj[38] sky130_fd_sc_hd__buf_8
XFILLER_25_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput661 _031_/Y vssd vssd vccd vccd la_data_in_mprj[48] sky130_fd_sc_hd__buf_8
Xoutput672 _041_/Y vssd vssd vccd vccd la_data_in_mprj[58] sky130_fd_sc_hd__buf_8
XFILLER_40_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput683 _051_/Y vssd vssd vccd vccd la_data_in_mprj[68] sky130_fd_sc_hd__buf_8
XFILLER_43_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput694 _061_/Y vssd vssd vccd vccd la_data_in_mprj[78] sky130_fd_sc_hd__buf_8
XFILLER_8_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__510__B _510_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1403 wire1403/A vssd vssd vccd vccd wire1403/X sky130_fd_sc_hd__buf_6
XFILLER_5_2734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1414 wire1414/A vssd vssd vccd vccd wire1414/X sky130_fd_sc_hd__buf_6
Xwire1425 input2/X vssd vssd vccd vccd _297_/B sky130_fd_sc_hd__buf_6
XTAP_190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1436 wire1436/A vssd vssd vccd vccd _385_/B sky130_fd_sc_hd__buf_6
XFILLER_25_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1447 wire1447/A vssd vssd vccd vccd wire1447/X sky130_fd_sc_hd__buf_6
XFILLER_5_2789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1458 wire1459/X vssd vssd vccd vccd _372_/B sky130_fd_sc_hd__buf_6
Xwire1469 wire1469/A vssd vssd vccd vccd wire1469/X sky130_fd_sc_hd__buf_6
XFILLER_28_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input115_A la_data_out_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__438__A_N _566_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__238__A _238_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_312_ _312_/A _312_/B vssd vssd vccd vccd _312_/X sky130_fd_sc_hd__and2_4
XFILLER_42_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_243_ _243_/A _243_/B vssd vssd vccd vccd _243_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput18 la_data_out_mprj[112] vssd vssd vccd vccd _481_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_input80_A la_data_out_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput29 la_data_out_mprj[122] vssd vssd vccd vccd _491_/C sky130_fd_sc_hd__clkbuf_4
X_174_ _174_/A _174_/B vssd vssd vccd vccd _174_/X sky130_fd_sc_hd__and2_4
XFILLER_10_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__404__C _404_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__420__B _420_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1758 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output501_A _388_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1132_A wire1133/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__148__A _148_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output870_A wire1224/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[13\] la_data_out_core[13] _176_/X vssd vssd vccd vccd _160_/A
+ sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_gates\[26\] mprj_dat_i_user[26] wire1248/X vssd vssd vccd vccd wire1008/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_18_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1599_A wire1600/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2198 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3711 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__611__A _611_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3755 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__330__B _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[124\] la_data_out_core[124] _287_/X vssd vssd vccd vccd _107_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_42_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__058__A _058_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_rebuffer3_A split13/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__505__B _505_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__521__A _521_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput480 _484_/X vssd vssd vccd vccd la_data_in_core[115] sky130_fd_sc_hd__buf_8
Xoutput491 _494_/X vssd vssd vccd vccd la_data_in_core[125] sky130_fd_sc_hd__buf_8
XFILLER_40_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__240__B _240_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1200 _324_/X vssd vssd vccd vccd wire1200/X sky130_fd_sc_hd__buf_6
Xwire1211 _316_/X vssd vssd vccd vccd wire1211/X sky130_fd_sc_hd__buf_6
XFILLER_43_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1222 _309_/X vssd vssd vccd vccd wire1222/X sky130_fd_sc_hd__buf_6
XANTENNA_input232_A la_iena_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1233 wire1234/X vssd vssd vccd vccd wire1233/X sky130_fd_sc_hd__buf_6
XFILLER_1_2417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1255 _265_/X vssd vssd vccd vccd wire1255/X sky130_fd_sc_hd__buf_6
Xwire1266 wire1266/A vssd vssd vccd vccd wire1266/X sky130_fd_sc_hd__buf_6
XFILLER_21_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1277 wire1277/A vssd vssd vccd vccd _294_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1288 wire1289/X vssd vssd vccd vccd _341_/B sky130_fd_sc_hd__buf_6
Xwire1299 wire1299/A vssd vssd vccd vccd wire1299/X sky130_fd_sc_hd__buf_6
XFILLER_21_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_226_ _226_/A _226_/B vssd vssd vccd vccd _226_/X sky130_fd_sc_hd__and2_4
XFILLER_7_621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__415__B _415_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_157_ _157_/A vssd vssd vccd vccd _157_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_3503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_088_ _088_/A vssd vssd vccd vccd _088_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_6_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output549_A wire1073/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1082_A _422_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output716_A _081_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1347_A wire1348/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__606__A _606_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__325__B _325_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire967_A _133_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__341__A _341_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput208 la_iena_mprj[53] vssd vssd vccd vccd _216_/B sky130_fd_sc_hd__clkbuf_4
Xinput219 la_iena_mprj[63] vssd vssd vccd vccd _226_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__516__A _516_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__235__B _235_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_011_ _011_/A vssd vssd vccd vccd _011_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input182_A la_iena_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__251__A _251_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input447_A mprj_dat_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input43_A la_data_out_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1030 wire1030/A vssd vssd vccd vccd _114_/A sky130_fd_sc_hd__buf_8
XFILLER_40_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1041 _611_/X vssd vssd vccd vccd wire1041/X sky130_fd_sc_hd__buf_6
XFILLER_5_2383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1052 _542_/X vssd vssd vccd vccd wire1052/X sky130_fd_sc_hd__buf_6
XFILLER_40_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1063 _463_/X vssd vssd vccd vccd wire1063/X sky130_fd_sc_hd__buf_6
Xwire1074 _430_/X vssd vssd vccd vccd wire1074/X sky130_fd_sc_hd__buf_6
XFILLER_21_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1085 _419_/X vssd vssd vccd vccd wire1085/X sky130_fd_sc_hd__buf_6
XFILLER_1_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1096 _408_/X vssd vssd vccd vccd wire1096/X sky130_fd_sc_hd__buf_6
XFILLER_35_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output499_A _386_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output666_A _035_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_209_ _209_/A _209_/B vssd vssd vccd vccd _209_/X sky130_fd_sc_hd__and2_2
XFILLER_45_4023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1297_A wire1297/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output833_A _585_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1464_A wire1465/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[80\] la_data_out_core[80] _243_/X vssd vssd vccd vccd _063_/A
+ sky130_fd_sc_hd__nand2_8
XTAP_734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1729_A wire1730/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__336__A _336_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[92\]_A la_data_out_core[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__071__A _071_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2863 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_560_ _560_/A _560_/B vssd vssd vccd vccd _560_/X sky130_fd_sc_hd__and2_4
XFILLER_45_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_491_ _619_/A _491_/B _491_/C vssd vssd vccd vccd _491_/X sky130_fd_sc_hd__and3b_4
XFILLER_0_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__246__A _246_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input397_A mprj_adr_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[83\]_A la_data_out_core[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1212_A wire1213/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output783_A _539_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output950_A wire1235/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[74\]_A la_data_out_core[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1518 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1679_A wire1679/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__603__B _603_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1458 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[2\]_B _165_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__471__A_N _599_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__066__A _066_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[65\]_A la_data_out_core[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__513__B _513_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input145_A la_iena_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_612_ _612_/A _612_/B vssd vssd vccd vccd _612_/X sky130_fd_sc_hd__and2_4
XANTENNA_input312_A la_oenb_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_543_ _543_/A _543_/B vssd vssd vccd vccd _543_/X sky130_fd_sc_hd__and2_4
XTAP_2932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_2339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_474_ _602_/A _474_/B _474_/C vssd vssd vccd vccd _474_/X sky130_fd_sc_hd__and3b_2
XTAP_2987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[56\]_A la_data_out_core[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output531_A wire1089/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output629_A _002_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1162_A wire1163/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3875 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput380 la_oenb_mprj[93] vssd vssd vccd vccd _590_/A sky130_fd_sc_hd__buf_4
XFILLER_20_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput391 mprj_adr_o_core[12] vssd vssd vccd vccd wire1414/A sky130_fd_sc_hd__buf_6
XANTENNA__494__A_N _622_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1427_A wire1427/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[43\] la_data_out_core[43] _206_/X vssd vssd vccd vccd _026_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_14_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[47\]_A la_data_out_core[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__614__A _614_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__333__B _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput810 _564_/X vssd vssd vccd vccd la_oenb_core[67] sky130_fd_sc_hd__buf_8
Xoutput821 _574_/X vssd vssd vccd vccd la_oenb_core[77] sky130_fd_sc_hd__buf_8
Xoutput832 _584_/X vssd vssd vccd vccd la_oenb_core[87] sky130_fd_sc_hd__buf_8
XFILLER_25_3523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput843 _594_/X vssd vssd vccd vccd la_oenb_core[97] sky130_fd_sc_hd__buf_8
XFILLER_9_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput854 wire1205/X vssd vssd vccd vccd mprj_adr_o_user[15] sky130_fd_sc_hd__buf_8
Xoutput865 wire1188/X vssd vssd vccd vccd mprj_adr_o_user[25] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[5\] la_data_out_core[5] _168_/X vssd vssd vccd vccd _152_/A
+ sky130_fd_sc_hd__nand2_1
Xoutput876 wire1219/X vssd vssd vccd vccd mprj_adr_o_user[6] sky130_fd_sc_hd__buf_8
Xoutput887 wire971/X vssd vssd vccd vccd mprj_dat_i_core[15] sky130_fd_sc_hd__buf_8
XFILLER_25_2822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput898 _139_/Y vssd vssd vccd vccd mprj_dat_i_core[25] sky130_fd_sc_hd__buf_8
XTAP_350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1607 wire1607/A vssd vssd vccd vccd _589_/B sky130_fd_sc_hd__buf_6
XFILLER_3_3341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1618 wire1618/A vssd vssd vccd vccd _578_/B sky130_fd_sc_hd__buf_6
XTAP_383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1629 wire1629/A vssd vssd vccd vccd _521_/B sky130_fd_sc_hd__buf_4
XFILLER_45_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__508__B _508_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_190_ _190_/A _190_/B vssd vssd vccd vccd _190_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[38\]_A la_data_out_core[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__524__A _524_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[122\]_A la_data_out_core[122] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_41_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__243__B _243_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input262_A la_oenb_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_526_ _526_/A _526_/B vssd vssd vccd vccd _526_/X sky130_fd_sc_hd__and2_4
XTAP_2773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1402 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_457_ _585_/A _457_/B _457_/C vssd vssd vccd vccd _457_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_388_ _516_/A _388_/B _388_/C vssd vssd vccd vccd _388_/X sky130_fd_sc_hd__and3b_4
XANTENNA_output481_A _485_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[29\]_A la_data_out_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output579_A wire1110/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_A la_data_out_core[113] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_35_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output746_A wire1035/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1377_A wire1377/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3707 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output913_A wire1174/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1544_A wire1544/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1711_A wire1711/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__609__A _609_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__328__B _328_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire997_A wire997/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[104\]_A la_data_out_core[104] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1134 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput640 _012_/Y vssd vssd vccd vccd la_data_in_mprj[29] sky130_fd_sc_hd__buf_8
Xoutput651 _022_/Y vssd vssd vccd vccd la_data_in_mprj[39] sky130_fd_sc_hd__buf_8
XFILLER_25_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput662 _032_/Y vssd vssd vccd vccd la_data_in_mprj[49] sky130_fd_sc_hd__buf_8
XFILLER_25_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput673 _042_/Y vssd vssd vccd vccd la_data_in_mprj[59] sky130_fd_sc_hd__buf_8
Xoutput684 _052_/Y vssd vssd vccd vccd la_data_in_mprj[69] sky130_fd_sc_hd__buf_8
XFILLER_40_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput695 _062_/Y vssd vssd vccd vccd la_data_in_mprj[79] sky130_fd_sc_hd__buf_8
XFILLER_5_2724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1404 wire1405/X vssd vssd vccd vccd _320_/B sky130_fd_sc_hd__buf_6
Xwire1415 wire1416/X vssd vssd vccd vccd _316_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1426 input1/X vssd vssd vccd vccd _296_/B sky130_fd_sc_hd__buf_6
XFILLER_25_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1437 wire1437/A vssd vssd vccd vccd _384_/B sky130_fd_sc_hd__buf_6
Xwire1448 wire1449/X vssd vssd vccd vccd _377_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1459 wire1459/A vssd vssd vccd vccd wire1459/X sky130_fd_sc_hd__buf_6
XFILLER_28_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__519__A _519_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__238__B _238_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input108_A la_data_out_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_311_ _311_/A _311_/B vssd vssd vccd vccd _311_/X sky130_fd_sc_hd__and2_2
XFILLER_35_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_242_ _242_/A _242_/B vssd vssd vccd vccd _242_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__254__A _254_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput19 la_data_out_mprj[113] vssd vssd vccd vccd _482_/C sky130_fd_sc_hd__clkbuf_4
X_173_ _173_/A _173_/B vssd vssd vccd vccd _173_/X sky130_fd_sc_hd__and2_4
XFILLER_32_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input73_A la_data_out_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__420__C _420_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1125_A _362_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_509_ _509_/A _509_/B vssd vssd vccd vccd _509_/X sky130_fd_sc_hd__and2_4
XFILLER_33_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output863_A wire1192/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__164__A _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[19\] mprj_dat_i_user[19] rebuffer5/X vssd vssd vccd vccd wire1020/A
+ sky130_fd_sc_hd__nand2_4
XANTENNA_wire1494_A wire1494/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1476 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1661_A wire1661/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__611__B _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[117\] la_data_out_core[117] _280_/X vssd vssd vccd vccd _100_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_0_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__339__A _339_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__074__A _074_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__521__B _521_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput470 _475_/X vssd vssd vccd vccd la_data_in_core[106] sky130_fd_sc_hd__buf_8
XFILLER_43_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput481 _485_/X vssd vssd vccd vccd la_data_in_core[116] sky130_fd_sc_hd__buf_8
Xoutput492 wire1055/X vssd vssd vccd vccd la_data_in_core[126] sky130_fd_sc_hd__buf_8
XFILLER_40_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__405__A_N _533_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1201 _323_/X vssd vssd vccd vccd wire1201/X sky130_fd_sc_hd__buf_6
Xwire1212 wire1213/X vssd vssd vccd vccd wire1212/X sky130_fd_sc_hd__buf_6
Xwire1223 _308_/X vssd vssd vccd vccd wire1223/X sky130_fd_sc_hd__buf_6
XFILLER_43_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1234 _301_/X vssd vssd vccd vccd wire1234/X sky130_fd_sc_hd__buf_6
XFILLER_1_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1245 wire1245/A vssd vssd vccd vccd wire1245/X sky130_fd_sc_hd__buf_8
XFILLER_5_2587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1256 _264_/X vssd vssd vccd vccd wire1256/X sky130_fd_sc_hd__buf_6
XFILLER_1_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1267 wire1268/X vssd vssd vccd vccd _299_/B sky130_fd_sc_hd__buf_6
XANTENNA_input225_A la_iena_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1278 wire1279/X vssd vssd vccd vccd _346_/B sky130_fd_sc_hd__buf_6
Xwire1289 wire1289/A vssd vssd vccd vccd wire1289/X sky130_fd_sc_hd__buf_6
XFILLER_34_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__249__A _249_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_225_ _225_/A _225_/B vssd vssd vccd vccd _225_/X sky130_fd_sc_hd__and2_4
XFILLER_7_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_156_ _156_/A vssd vssd vccd vccd _156_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_087_ _087_/A vssd vssd vccd vccd _087_/Y sky130_fd_sc_hd__inv_4
XFILLER_45_3559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__431__B _431_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output611_A _101_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output709_A _074_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1242_A _296_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__159__A _159_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1507_A wire1507/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__606__B _606_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__622__A _622_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__428__A_N _556_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__341__B _341_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput209 la_iena_mprj[54] vssd vssd vccd vccd _217_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1022 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__069__A _069_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_710 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__516__B _516_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_010_ _010_/A vssd vssd vccd vccd _010_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_4007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__532__A _532_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input175_A la_iena_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input342_A la_oenb_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input36_A la_data_out_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1718 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1020 wire1020/A vssd vssd vccd vccd _133_/A sky130_fd_sc_hd__buf_6
XFILLER_0_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1031 wire1031/A vssd vssd vccd vccd _146_/A sky130_fd_sc_hd__buf_8
XFILLER_22_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1042 _607_/X vssd vssd vccd vccd wire1042/X sky130_fd_sc_hd__buf_6
XFILLER_2_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1053 _523_/X vssd vssd vccd vccd wire1053/X sky130_fd_sc_hd__buf_6
XFILLER_5_2395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1064 _461_/X vssd vssd vccd vccd wire1064/X sky130_fd_sc_hd__buf_6
XFILLER_38_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1075 _429_/X vssd vssd vccd vccd wire1075/X sky130_fd_sc_hd__buf_6
Xwire1086 _418_/X vssd vssd vccd vccd wire1086/X sky130_fd_sc_hd__buf_6
Xwire1097 _407_/X vssd vssd vccd vccd wire1097/X sky130_fd_sc_hd__buf_6
XFILLER_21_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_208_ _208_/A _208_/B vssd vssd vccd vccd _208_/X sky130_fd_sc_hd__and2_2
XFILLER_32_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output561_A _442_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output659_A _029_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_139_ _139_/A vssd vssd vccd vccd _139_/Y sky130_fd_sc_hd__inv_4
XANTENNA_wire1192_A wire1193/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output826_A _578_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1457_A wire1457/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[73\] la_data_out_core[73] _236_/X vssd vssd vccd vccd _056_/A
+ sky130_fd_sc_hd__nand2_8
XTAP_779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__617__A _617_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__336__B _336_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[92\]_B _255_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_490_ _618_/A _490_/B _490_/C vssd vssd vccd vccd _490_/X sky130_fd_sc_hd__and3b_4
Xsplit13 split13/A vssd vssd vccd vccd split13/X sky130_fd_sc_hd__buf_4
XANTENNA__527__A _527_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__246__B _246_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input292_A la_oenb_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[83\]_B _246_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__262__A _262_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1891 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1038_A _616_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1205_A _320_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output776_A _533_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[74\]_B _237_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output943_A wire1158/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__172__A _172_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1574_A wire1575/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[65\]_B _228_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__082__A _082_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4030 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input138_A la_iena_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_611_ _611_/A _611_/B vssd vssd vccd vccd _611_/X sky130_fd_sc_hd__and2_2
XTAP_3623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_542_ _542_/A _542_/B vssd vssd vccd vccd _542_/X sky130_fd_sc_hd__and2_1
XTAP_3678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input305_A la_oenb_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__257__A _257_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_473_ _601_/A _473_/B _473_/C vssd vssd vccd vccd _473_/X sky130_fd_sc_hd__and3b_4
XFILLER_44_189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3664 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[56\]_B _219_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__423__C _423_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output524_A _372_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1155_A _347_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput370 la_oenb_mprj[84] vssd vssd vccd vccd _581_/A sky130_fd_sc_hd__buf_4
Xinput381 la_oenb_mprj[94] vssd vssd vccd vccd _591_/A sky130_fd_sc_hd__clkbuf_4
Xinput392 mprj_adr_o_core[13] vssd vssd vccd vccd wire1412/A sky130_fd_sc_hd__buf_6
XFILLER_36_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1322_A wire1323/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output893_A wire966/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__167__A _167_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[36\] la_data_out_core[36] _199_/X vssd vssd vccd vccd _019_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_3564 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2006 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1691_A wire1692/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__614__B _614_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput800 wire1049/X vssd vssd vccd vccd la_oenb_core[58] sky130_fd_sc_hd__buf_8
Xoutput811 _565_/X vssd vssd vccd vccd la_oenb_core[68] sky130_fd_sc_hd__buf_8
XFILLER_9_3732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput822 _575_/X vssd vssd vccd vccd la_oenb_core[78] sky130_fd_sc_hd__buf_8
Xoutput833 _585_/X vssd vssd vccd vccd la_oenb_core[88] sky130_fd_sc_hd__buf_8
XFILLER_25_3513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput844 _595_/X vssd vssd vccd vccd la_oenb_core[98] sky130_fd_sc_hd__buf_8
Xoutput855 wire1204/X vssd vssd vccd vccd mprj_adr_o_user[16] sky130_fd_sc_hd__buf_8
XFILLER_9_3776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput866 wire1186/X vssd vssd vccd vccd mprj_adr_o_user[26] sky130_fd_sc_hd__buf_8
Xoutput877 wire1218/X vssd vssd vccd vccd mprj_adr_o_user[7] sky130_fd_sc_hd__buf_8
Xoutput888 wire970/X vssd vssd vccd vccd mprj_dat_i_core[16] sky130_fd_sc_hd__buf_8
Xoutput899 _140_/Y vssd vssd vccd vccd mprj_dat_i_core[26] sky130_fd_sc_hd__buf_8
XFILLER_45_2271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1608 wire1608/A vssd vssd vccd vccd _588_/B sky130_fd_sc_hd__buf_6
XFILLER_42_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1619 wire1619/A vssd vssd vccd vccd _577_/B sky130_fd_sc_hd__buf_6
XTAP_373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__077__A _077_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__524__B _524_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[122\]_B _285_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__540__A _540_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input255_A la_iena_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input422_A mprj_dat_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[31\]_A mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_525_ _525_/A _525_/B vssd vssd vccd vccd _525_/X sky130_fd_sc_hd__and2_4
XTAP_2763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_456_ _584_/A _456_/B _456_/C vssd vssd vccd vccd _456_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_387_ _515_/A _387_/B _387_/C vssd vssd vccd vccd _387_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__434__B _434_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_B _276_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output474_A _379_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output739_A wire1039/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1272_A wire1272/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__461__A_N _589_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output906_A wire983/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1537_A wire1537/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__609__B _609_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1704_A wire1704/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[22\]_A mprj_dat_i_user[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__625__A _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1558 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__344__B _344_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_B wire1253/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput630 _148_/Y vssd vssd vccd vccd la_data_in_mprj[1] sky130_fd_sc_hd__buf_8
XANTENNA__360__A _360_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput641 _149_/Y vssd vssd vccd vccd la_data_in_mprj[2] sky130_fd_sc_hd__buf_8
XFILLER_44_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput652 _150_/Y vssd vssd vccd vccd la_data_in_mprj[3] sky130_fd_sc_hd__buf_8
Xoutput663 _151_/Y vssd vssd vccd vccd la_data_in_mprj[4] sky130_fd_sc_hd__buf_8
XFILLER_9_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput674 _152_/Y vssd vssd vccd vccd la_data_in_mprj[5] sky130_fd_sc_hd__buf_8
Xoutput685 _153_/Y vssd vssd vccd vccd la_data_in_mprj[6] sky130_fd_sc_hd__buf_8
Xoutput696 _154_/Y vssd vssd vccd vccd la_data_in_mprj[7] sky130_fd_sc_hd__buf_8
XFILLER_5_2714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1405 wire1406/X vssd vssd vccd vccd wire1405/X sky130_fd_sc_hd__buf_6
Xwire1416 wire1416/A vssd vssd vccd vccd wire1416/X sky130_fd_sc_hd__buf_6
Xwire1427 wire1427/A vssd vssd vccd vccd _394_/B sky130_fd_sc_hd__buf_6
Xwire1438 wire1438/A vssd vssd vccd vccd _383_/B sky130_fd_sc_hd__buf_6
XFILLER_41_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1449 wire1449/A vssd vssd vccd vccd wire1449/X sky130_fd_sc_hd__buf_6
XFILLER_46_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__519__B _519_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[13\]_A mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ _310_/A _310_/B vssd vssd vccd vccd _310_/X sky130_fd_sc_hd__and2_4
XFILLER_42_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__535__A _535_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_241_ _241_/A _241_/B vssd vssd vccd vccd _241_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_172_ _172_/A _172_/B vssd vssd vccd vccd _172_/X sky130_fd_sc_hd__and2_4
XFILLER_10_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input372_A la_oenb_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__484__A_N _612_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input66_A la_data_out_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__270__A _270_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1462 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_508_ _508_/A _508_/B vssd vssd vccd vccd _508_/X sky130_fd_sc_hd__and2_4
XTAP_2582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1020_A wire1020/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1118_A wire1119/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output689_A _056_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_439_ _567_/A _439_/B _439_/C vssd vssd vccd vccd _439_/X sky130_fd_sc_hd__and3b_2
XFILLER_18_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__164__B _164_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output856_A wire1202/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1487_A wire1488/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__180__A _180_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1654_A wire1654/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__339__B _339_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__355__A _355_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__090__A _090_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput471 _476_/X vssd vssd vccd vccd la_data_in_core[107] sky130_fd_sc_hd__buf_8
Xoutput482 _486_/X vssd vssd vccd vccd la_data_in_core[117] sky130_fd_sc_hd__buf_8
Xoutput493 wire1054/X vssd vssd vccd vccd la_data_in_core[127] sky130_fd_sc_hd__buf_8
XFILLER_40_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1202 wire1203/X vssd vssd vccd vccd wire1202/X sky130_fd_sc_hd__buf_6
Xwire1213 wire1214/X vssd vssd vccd vccd wire1213/X sky130_fd_sc_hd__buf_6
XFILLER_21_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1224 _307_/X vssd vssd vccd vccd wire1224/X sky130_fd_sc_hd__buf_6
Xwire1235 wire1236/X vssd vssd vccd vccd wire1235/X sky130_fd_sc_hd__buf_6
Xwire1257 _263_/X vssd vssd vccd vccd wire1257/X sky130_fd_sc_hd__buf_6
XFILLER_38_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1268 wire1268/A vssd vssd vccd vccd wire1268/X sky130_fd_sc_hd__buf_6
XFILLER_25_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1279 wire1279/A vssd vssd vccd vccd wire1279/X sky130_fd_sc_hd__buf_6
XFILLER_28_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__249__B _249_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input120_A la_data_out_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input218_A la_iena_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__265__A _265_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_224_ _224_/A _224_/B vssd vssd vccd vccd _224_/X sky130_fd_sc_hd__and2_4
XFILLER_11_652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_155_ _155_/A vssd vssd vccd vccd _155_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[1\] mprj_dat_i_user[1] max_cap1244/X vssd vssd vccd vccd wire1019/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_7_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_086_ _086_/A vssd vssd vccd vccd _086_/Y sky130_fd_sc_hd__inv_4
XFILLER_45_2815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__431__C _431_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3908 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output604_A _094_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1235_A wire1236/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1402_A wire1403/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__175__A _175_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_980 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[31\] mprj_dat_i_user[31] wire1248/X vssd vssd vccd vccd wire999/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_30_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__622__B _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1034 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3092 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__085__A _085_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__532__B _532_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input168_A la_iena_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input335_A la_oenb_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1010 wire1011/X vssd vssd vccd vccd _138_/A sky130_fd_sc_hd__buf_6
Xwire1021 wire1021/A vssd vssd vccd vccd _132_/A sky130_fd_sc_hd__buf_6
Xwire1032 _624_/X vssd vssd vccd vccd wire1032/X sky130_fd_sc_hd__buf_6
Xwire1043 _605_/X vssd vssd vccd vccd wire1043/X sky130_fd_sc_hd__buf_6
XANTENNA_input29_A la_data_out_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1054 _496_/X vssd vssd vccd vccd wire1054/X sky130_fd_sc_hd__buf_6
XFILLER_2_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1065 _460_/X vssd vssd vccd vccd wire1065/X sky130_fd_sc_hd__buf_6
Xwire1076 _428_/X vssd vssd vccd vccd wire1076/X sky130_fd_sc_hd__buf_6
XFILLER_1_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1087 _417_/X vssd vssd vccd vccd wire1087/X sky130_fd_sc_hd__buf_6
XFILLER_38_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1098 _406_/X vssd vssd vccd vccd wire1098/X sky130_fd_sc_hd__buf_6
XFILLER_21_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__426__C _426_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_207_ _207_/A _207_/B vssd vssd vccd vccd _207_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3250 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__442__B _442_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_138_ _138_/A vssd vssd vccd vccd _138_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_32_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output554_A _436_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_069_ _069_/A vssd vssd vccd vccd _069_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output721_A wire1045/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output819_A _572_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1352_A wire1353/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[66\] la_data_out_core[66] _229_/X vssd vssd vccd vccd _049_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_39_858 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1617_A wire1617/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__617__B _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire972_A _128_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__352__B _352_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[5\]_A mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1410 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[5\]_A la_data_out_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__527__B _527_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__543__A _543_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input285_A la_oenb_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input452_A mprj_dat_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__437__B _437_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__418__A_N _546_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output671_A _040_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output769_A _499_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__172__B _172_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output936_A wire1114/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__347__B _347_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__363__A _363_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_610_ _610_/A _610_/B vssd vssd vccd vccd _610_/X sky130_fd_sc_hd__and2_4
XTAP_3613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__538__A _538_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_541_ _541_/A _541_/B vssd vssd vccd vccd _541_/X sky130_fd_sc_hd__and2_4
XTAP_2912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input200_A la_iena_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_472_ _600_/A _472_/B _472_/C vssd vssd vccd vccd _472_/X sky130_fd_sc_hd__and3b_4
XTAP_2978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input96_A la_data_out_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__273__A _273_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3676 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output517_A wire1102/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput360 la_oenb_mprj[75] vssd vssd vccd vccd _572_/A sky130_fd_sc_hd__buf_4
XFILLER_42_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput371 la_oenb_mprj[85] vssd vssd vccd vccd _582_/A sky130_fd_sc_hd__buf_4
XFILLER_40_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput382 la_oenb_mprj[95] vssd vssd vccd vccd _592_/A sky130_fd_sc_hd__clkbuf_4
Xinput393 mprj_adr_o_core[14] vssd vssd vccd vccd wire1409/A sky130_fd_sc_hd__buf_6
XANTENNA_wire1148_A wire1149/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__167__B _167_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1315_A wire1315/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output886_A wire972/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[29\] la_data_out_core[29] _192_/X vssd vssd vccd vccd _012_/A
+ sky130_fd_sc_hd__nand2_2
XANTENNA__390__A_N _518_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__183__A _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1684_A wire1685/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput801 _556_/X vssd vssd vccd vccd la_oenb_core[59] sky130_fd_sc_hd__buf_8
Xoutput812 _566_/X vssd vssd vccd vccd la_oenb_core[69] sky130_fd_sc_hd__buf_8
Xoutput823 _576_/X vssd vssd vccd vccd la_oenb_core[79] sky130_fd_sc_hd__buf_8
XFILLER_9_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput834 _586_/X vssd vssd vccd vccd la_oenb_core[89] sky130_fd_sc_hd__buf_8
Xoutput845 _596_/X vssd vssd vccd vccd la_oenb_core[99] sky130_fd_sc_hd__buf_8
Xoutput856 wire1202/X vssd vssd vccd vccd mprj_adr_o_user[17] sky130_fd_sc_hd__buf_8
XFILLER_5_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput867 wire1184/X vssd vssd vccd vccd mprj_adr_o_user[27] sky130_fd_sc_hd__buf_8
XFILLER_9_3788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput878 wire1217/X vssd vssd vccd vccd mprj_adr_o_user[8] sky130_fd_sc_hd__buf_8
XFILLER_29_2982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput889 wire969/X vssd vssd vccd vccd mprj_dat_i_core[17] sky130_fd_sc_hd__buf_8
XFILLER_3_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1609 wire1609/A vssd vssd vccd vccd _587_/B sky130_fd_sc_hd__buf_6
XTAP_374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xrebuffer10 wire1245/A vssd vssd vccd vccd rebuffer10/X sky130_fd_sc_hd__bufbuf_8
XANTENNA__358__A _358_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_2330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__093__A _093_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__540__B _540_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input150_A la_iena_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2564 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input248_A la_iena_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input415_A mprj_adr_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__268__A _268_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input11_A la_data_out_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[31\]_B wire1248/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_524_ _524_/A _524_/B vssd vssd vccd vccd _524_/X sky130_fd_sc_hd__and2_4
XTAP_2742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_455_ _583_/A _455_/B _455_/C vssd vssd vccd vccd _455_/X sky130_fd_sc_hd__and3b_4
XTAP_2797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_386_ _514_/A _386_/B _386_/C vssd vssd vccd vccd _386_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_3451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__434__C _434_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output467_A wire1057/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__450__B _450_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output634_A _006_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1265_A wire1266/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output801_A _556_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1432_A wire1432/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput190 la_iena_mprj[37] vssd vssd vccd vccd _200_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__178__A _178_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1198 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__625__B _625_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput620 _109_/Y vssd vssd vccd vccd la_data_in_mprj[126] sky130_fd_sc_hd__buf_8
XFILLER_27_2908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput631 _003_/Y vssd vssd vccd vccd la_data_in_mprj[20] sky130_fd_sc_hd__buf_8
XANTENNA__360__B _360_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput642 _013_/Y vssd vssd vccd vccd la_data_in_mprj[30] sky130_fd_sc_hd__buf_8
XFILLER_44_3967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput653 _023_/Y vssd vssd vccd vccd la_data_in_mprj[40] sky130_fd_sc_hd__buf_8
Xoutput664 _033_/Y vssd vssd vccd vccd la_data_in_mprj[50] sky130_fd_sc_hd__buf_8
XFILLER_25_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput675 _043_/Y vssd vssd vccd vccd la_data_in_mprj[60] sky130_fd_sc_hd__buf_8
XFILLER_9_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput686 _053_/Y vssd vssd vccd vccd la_data_in_mprj[70] sky130_fd_sc_hd__buf_8
Xoutput697 _063_/Y vssd vssd vccd vccd la_data_in_mprj[80] sky130_fd_sc_hd__buf_8
XFILLER_28_1043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1406 wire1406/A vssd vssd vccd vccd wire1406/X sky130_fd_sc_hd__buf_6
XANTENNA_input3_A caravel_rstn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1417 wire1417/A vssd vssd vccd vccd _315_/B sky130_fd_sc_hd__buf_6
XTAP_182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1428 wire1428/A vssd vssd vccd vccd _393_/B sky130_fd_sc_hd__buf_6
XFILLER_25_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1439 wire1439/A vssd vssd vccd vccd _382_/B sky130_fd_sc_hd__buf_6
XFILLER_25_1975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__088__A _088_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_240_ _240_/A _240_/B vssd vssd vccd vccd _240_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__535__B _535_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_171_ _171_/A _171_/B vssd vssd vccd vccd _171_/X sky130_fd_sc_hd__and2_4
XFILLER_10_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input198_A la_iena_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__551__A _551_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input365_A la_oenb_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_irq_gates\[0\] user_irq_core[0] _291_/X vssd vssd vccd vccd _111_/A sky130_fd_sc_hd__nand2_2
XANTENNA_input59_A la_data_out_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3502 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_507_ _507_/A _507_/B vssd vssd vccd vccd _507_/X sky130_fd_sc_hd__and2_4
XTAP_2583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__445__B _445_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_438_ _566_/A _438_/B _438_/C vssd vssd vccd vccd _438_/X sky130_fd_sc_hd__and3b_4
XANTENNA_output584_A wire1063/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_369_ _497_/A _369_/B _369_/C vssd vssd vccd vccd _369_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output751_A _510_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xrebuffer1 wire1245/X vssd vssd vccd vccd rebuffer1/X sky130_fd_sc_hd__buf_8
XANTENNA_output849_A wire1212/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1382_A wire1383/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__180__B _180_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[96\] la_data_out_core[96] wire1259/X vssd vssd vccd vccd _079_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_26_3653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1647_A wire1647/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__355__B _355_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput472 _477_/X vssd vssd vccd vccd la_data_in_core[108] sky130_fd_sc_hd__buf_8
Xoutput483 _487_/X vssd vssd vccd vccd la_data_in_core[118] sky130_fd_sc_hd__buf_8
Xoutput494 _381_/X vssd vssd vccd vccd la_data_in_core[12] sky130_fd_sc_hd__buf_8
XFILLER_9_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1203 _322_/X vssd vssd vccd vccd wire1203/X sky130_fd_sc_hd__buf_6
Xwire1214 _315_/X vssd vssd vccd vccd wire1214/X sky130_fd_sc_hd__buf_6
Xwire1225 _306_/X vssd vssd vccd vccd wire1225/X sky130_fd_sc_hd__buf_6
Xwire1236 _300_/X vssd vssd vccd vccd wire1236/X sky130_fd_sc_hd__buf_6
XFILLER_5_2578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1258 _262_/X vssd vssd vccd vccd wire1258/X sky130_fd_sc_hd__buf_6
Xwire1269 wire1270/X vssd vssd vccd vccd _304_/B sky130_fd_sc_hd__buf_6
XFILLER_21_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input113_A la_data_out_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__546__A _546_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__451__A_N _579_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_223_ _223_/A _223_/B vssd vssd vccd vccd _223_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2466 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_154_ _154_/A vssd vssd vccd vccd _154_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__281__A _281_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_085_ _085_/A vssd vssd vccd vccd _085_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_6_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1130_A wire1131/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1228_A _304_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output799_A _554_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1610 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__175__B _175_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[11\] la_data_out_core[11] _174_/X vssd vssd vccd vccd _158_/A
+ sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_gates\[24\] mprj_dat_i_user[24] split13/X vssd vssd vccd vccd wire1011/A
+ sky130_fd_sc_hd__nand2_2
XANTENNA_wire1597_A wire1597/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__191__A _191_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3314 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2832 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[122\] la_data_out_core[122] _285_/X vssd vssd vccd vccd _105_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_25_1046 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__474__A_N _602_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__366__A _366_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[95\]_A la_data_out_core[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1000 wire1000/A vssd vssd vccd vccd _144_/A sky130_fd_sc_hd__buf_6
XFILLER_27_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1011 wire1011/A vssd vssd vccd vccd wire1011/X sky130_fd_sc_hd__buf_6
XFILLER_21_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1022 wire1022/A vssd vssd vccd vccd _131_/A sky130_fd_sc_hd__buf_8
XANTENNA_input230_A la_iena_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1033 _623_/X vssd vssd vccd vccd wire1033/X sky130_fd_sc_hd__buf_6
XANTENNA_input328_A la_oenb_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1044 _600_/X vssd vssd vccd vccd wire1044/X sky130_fd_sc_hd__buf_6
XFILLER_22_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1055 _495_/X vssd vssd vccd vccd wire1055/X sky130_fd_sc_hd__buf_6
XFILLER_1_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1066 _459_/X vssd vssd vccd vccd wire1066/X sky130_fd_sc_hd__buf_6
XFILLER_2_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1077 _427_/X vssd vssd vccd vccd wire1077/X sky130_fd_sc_hd__buf_6
XFILLER_21_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1088 _416_/X vssd vssd vccd vccd wire1088/X sky130_fd_sc_hd__buf_6
Xwire1099 _405_/X vssd vssd vccd vccd wire1099/X sky130_fd_sc_hd__buf_6
XFILLER_18_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__276__A _276_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[86\]_A la_data_out_core[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_206_ _206_/A _206_/B vssd vssd vccd vccd _206_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_137_ _137_/A vssd vssd vccd vccd _137_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_3295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__442__C _442_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_068_ _068_/A vssd vssd vccd vccd _068_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_2594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output547_A wire1075/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1080_A _424_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1178_A wire1179/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output714_A _079_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[10\]_A la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1345_A wire1345/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[59\] la_data_out_core[59] _222_/X vssd vssd vccd vccd _042_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_19_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__186__A _186_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_A la_data_out_core[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[5\]_B _168_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__096__A _096_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[68\]_A la_data_out_core[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__543__B _543_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input180_A la_iena_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input278_A la_oenb_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input445_A mprj_dat_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input41_A la_data_out_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__437__C _437_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_A la_data_out_core[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output497_A _384_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__453__B _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output664_A _033_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output831_A _583_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output929_A wire1126/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1462_A wire1463/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__363__B _363_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1230 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__538__B _538_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_540_ _540_/A _540_/B vssd vssd vccd vccd _540_/X sky130_fd_sc_hd__and2_4
XTAP_2913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_471_ _599_/A _471_/B _471_/C vssd vssd vccd vccd _471_/X sky130_fd_sc_hd__and3b_2
XFILLER_32_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[125\]_A la_data_out_core[125] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__554__A _554_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input395_A mprj_adr_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input89_A la_data_out_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput350 la_oenb_mprj[66] vssd vssd vccd vccd _563_/A sky130_fd_sc_hd__clkbuf_8
Xinput361 la_oenb_mprj[76] vssd vssd vccd vccd _573_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_1408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput372 la_oenb_mprj[86] vssd vssd vccd vccd _583_/A sky130_fd_sc_hd__clkbuf_4
Xinput383 la_oenb_mprj[96] vssd vssd vccd vccd _593_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput394 mprj_adr_o_core[15] vssd vssd vccd vccd wire1406/A sky130_fd_sc_hd__buf_6
XFILLER_36_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__448__B _448_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1210_A wire1211/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output781_A _537_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1308_A wire1309/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output879_A wire1215/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_A la_data_out_core[116] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__183__B _183_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1677_A wire1677/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput802 _502_/X vssd vssd vccd vccd la_oenb_core[5] sky130_fd_sc_hd__buf_8
Xoutput813 _503_/X vssd vssd vccd vccd la_oenb_core[6] sky130_fd_sc_hd__buf_8
Xoutput824 _504_/X vssd vssd vccd vccd la_oenb_core[7] sky130_fd_sc_hd__buf_8
Xoutput835 _505_/X vssd vssd vccd vccd la_oenb_core[8] sky130_fd_sc_hd__buf_8
XFILLER_6_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput846 _506_/X vssd vssd vccd vccd la_oenb_core[9] sky130_fd_sc_hd__buf_8
XFILLER_25_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput857 wire1201/X vssd vssd vccd vccd mprj_adr_o_user[18] sky130_fd_sc_hd__buf_8
XFILLER_3_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput868 wire1182/X vssd vssd vccd vccd mprj_adr_o_user[28] sky130_fd_sc_hd__buf_8
XFILLER_28_1225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput879 wire1215/X vssd vssd vccd vccd mprj_adr_o_user[9] sky130_fd_sc_hd__buf_8
XFILLER_8_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_604 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xrebuffer11 wire1245/A vssd vssd vccd vccd rebuffer11/X sky130_fd_sc_hd__bufbuf_8
XANTENNA__358__B _358_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[107\]_A la_data_out_core[107] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_17_2375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1251 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__408__A_N _536_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input143_A la_iena_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__549__A _549_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input310_A la_oenb_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input408_A mprj_adr_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3842 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_523_ _523_/A _523_/B vssd vssd vccd vccd _523_/X sky130_fd_sc_hd__and2_1
XTAP_3488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_454_ _582_/A _454_/B _454_/C vssd vssd vccd vccd _454_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__284__A _284_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_385_ _513_/A _385_/B _385_/C vssd vssd vccd vccd _385_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_2306 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__450__C _450_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output627_A _000_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1160_A wire1161/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput180 la_iena_mprj[28] vssd vssd vccd vccd _191_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput191 la_iena_mprj[38] vssd vssd vccd vccd _201_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[41\] la_data_out_core[41] _204_/X vssd vssd vccd vccd _024_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_24_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__194__A _194_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput610 _100_/Y vssd vssd vccd vccd la_data_in_mprj[117] sky130_fd_sc_hd__buf_8
XFILLER_5_4107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput621 _110_/Y vssd vssd vccd vccd la_data_in_mprj[127] sky130_fd_sc_hd__buf_8
XFILLER_25_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput632 _004_/Y vssd vssd vccd vccd la_data_in_mprj[21] sky130_fd_sc_hd__buf_8
Xoutput643 _014_/Y vssd vssd vccd vccd la_data_in_mprj[31] sky130_fd_sc_hd__buf_8
Xoutput654 _024_/Y vssd vssd vccd vccd la_data_in_mprj[41] sky130_fd_sc_hd__buf_8
XFILLER_5_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput665 _034_/Y vssd vssd vccd vccd la_data_in_mprj[51] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[3\] la_data_out_core[3] _166_/X vssd vssd vccd vccd _150_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_44_3979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput676 _044_/Y vssd vssd vccd vccd la_data_in_mprj[61] sky130_fd_sc_hd__buf_8
Xoutput687 wire991/X vssd vssd vccd vccd la_data_in_mprj[71] sky130_fd_sc_hd__buf_8
XFILLER_25_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput698 _064_/Y vssd vssd vccd vccd la_data_in_mprj[81] sky130_fd_sc_hd__buf_8
XFILLER_45_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1407 wire1408/X vssd vssd vccd vccd _319_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1418 wire1419/X vssd vssd vccd vccd _305_/B sky130_fd_sc_hd__buf_6
XFILLER_25_1943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1429 wire1429/A vssd vssd vccd vccd _392_/B sky130_fd_sc_hd__buf_6
XTAP_183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_170_ _170_/A _170_/B vssd vssd vccd vccd _170_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input260_A la_oenb_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input358_A la_oenb_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__380__A_N _508_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__279__A _279_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_506_ _506_/A _506_/B vssd vssd vccd vccd _506_/X sky130_fd_sc_hd__and2_4
XTAP_2562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_437_ _565_/A _437_/B _437_/C vssd vssd vccd vccd _437_/X sky130_fd_sc_hd__and3b_2
XANTENNA__445__C _445_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_368_ _368_/A _368_/B vssd vssd vccd vccd _368_/X sky130_fd_sc_hd__and2_4
XFILLER_13_3282 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output577_A _457_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_299_ _299_/A _299_/B vssd vssd vccd vccd _299_/X sky130_fd_sc_hd__and2_4
Xrebuffer2 wire1245/X vssd vssd vccd vccd rebuffer2/X sky130_fd_sc_hd__buf_4
XFILLER_31_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__461__B _461_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output744_A wire1037/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1375_A wire1375/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1807 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output911_A wire978/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[89\] la_data_out_core[89] _252_/X vssd vssd vccd vccd _072_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1542_A wire1542/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__189__A _189_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire995_A wire995/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__371__B _371_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput473 _478_/X vssd vssd vccd vccd la_data_in_core[109] sky130_fd_sc_hd__buf_8
Xoutput484 _488_/X vssd vssd vccd vccd la_data_in_core[119] sky130_fd_sc_hd__buf_8
XFILLER_44_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput495 _382_/X vssd vssd vccd vccd la_data_in_core[13] sky130_fd_sc_hd__buf_8
Xwire1204 _321_/X vssd vssd vccd vccd wire1204/X sky130_fd_sc_hd__buf_6
XFILLER_25_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__099__A _099_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1215 wire1216/X vssd vssd vccd vccd wire1215/X sky130_fd_sc_hd__buf_6
XFILLER_40_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1226 _305_/X vssd vssd vccd vccd wire1226/X sky130_fd_sc_hd__buf_6
XFILLER_19_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1237 wire1238/X vssd vssd vccd vccd wire1237/X sky130_fd_sc_hd__buf_6
XFILLER_21_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1248 wire1249/X vssd vssd vccd vccd wire1248/X sky130_fd_sc_hd__buf_8
Xwire1259 _259_/X vssd vssd vccd vccd wire1259/X sky130_fd_sc_hd__buf_6
XFILLER_41_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__546__B _546_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input106_A la_data_out_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_222_ _222_/A _222_/B vssd vssd vccd vccd _222_/X sky130_fd_sc_hd__and2_4
XFILLER_8_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__562__A _562_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2478 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_153_ _153_/A vssd vssd vccd vccd _153_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__281__B _281_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input71_A la_data_out_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_084_ _084_/A vssd vssd vccd vccd _084_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__456__B _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1123_A _363_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output694_A _061_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output861_A wire1196/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1210 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[17\] mprj_dat_i_user[17] rebuffer3/X vssd vssd vccd vccd wire1022/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA_wire1492_A wire1492/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[115\] la_data_out_core[115] _278_/X vssd vssd vccd vccd _098_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_39_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__366__B _366_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[95\]_B wire1260/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1001 wire1001/A vssd vssd vccd vccd _116_/A sky130_fd_sc_hd__buf_8
XFILLER_25_2271 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1012 wire1013/X vssd vssd vccd vccd _137_/A sky130_fd_sc_hd__buf_6
XFILLER_22_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1023 wire1023/A vssd vssd vccd vccd _130_/A sky130_fd_sc_hd__buf_8
Xwire1034 _622_/X vssd vssd vccd vccd wire1034/X sky130_fd_sc_hd__buf_6
XFILLER_43_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1045 _598_/X vssd vssd vccd vccd wire1045/X sky130_fd_sc_hd__buf_6
XFILLER_21_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1056 _474_/X vssd vssd vccd vccd wire1056/X sky130_fd_sc_hd__buf_6
XFILLER_25_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1067 _458_/X vssd vssd vccd vccd wire1067/X sky130_fd_sc_hd__buf_6
XANTENNA_input223_A la_iena_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1078 _426_/X vssd vssd vccd vccd wire1078/X sky130_fd_sc_hd__buf_6
XFILLER_38_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1089 _415_/X vssd vssd vccd vccd wire1089/X sky130_fd_sc_hd__buf_6
XANTENNA__557__A _557_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[86\]_B _249_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__292__A _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_205_ _205_/A _205_/B vssd vssd vccd vccd _205_/X sky130_fd_sc_hd__and2_2
XFILLER_7_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_136_ _136_/A vssd vssd vccd vccd _136_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_7_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_067_ _067_/A vssd vssd vccd vccd _067_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_7_3843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[10\]_B _173_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1338_A wire1339/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1590 wire1590/A vssd vssd vccd vccd _603_/B sky130_fd_sc_hd__buf_6
XFILLER_4_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__186__B _186_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1505_A wire1505/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_B _240_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_2451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__441__A_N _569_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[68\]_B _231_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input173_A la_iena_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input340_A la_oenb_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input438_A mprj_dat_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input34_A la_data_out_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__287__A _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_B _222_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__453__C _453_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output657_A _027_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_119_ _119_/A vssd vssd vccd vccd _119_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_32_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1190_A wire1191/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1288_A wire1289/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__464__A_N _592_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output824_A _504_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1455_A wire1455/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[71\] la_data_out_core[71] _234_/X vssd vssd vccd vccd _054_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_7_2972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__197__A _197_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2502 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1242 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_470_ _598_/A _470_/B _470_/C vssd vssd vccd vccd _470_/X sky130_fd_sc_hd__and3b_4
XTAP_2947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[125\]_B _288_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input290_A la_oenb_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input388_A mprj_adr_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__487__A_N _615_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__570__A _570_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3638 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput340 la_oenb_mprj[57] vssd vssd vccd vccd _554_/A sky130_fd_sc_hd__buf_4
Xinput351 la_oenb_mprj[67] vssd vssd vccd vccd _564_/A sky130_fd_sc_hd__clkbuf_8
Xinput362 la_oenb_mprj[77] vssd vssd vccd vccd _574_/A sky130_fd_sc_hd__buf_4
Xinput373 la_oenb_mprj[87] vssd vssd vccd vccd _584_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput384 la_oenb_mprj[97] vssd vssd vccd vccd _594_/A sky130_fd_sc_hd__clkbuf_4
Xinput395 mprj_adr_o_core[16] vssd vssd vccd vccd wire1403/A sky130_fd_sc_hd__buf_6
XFILLER_40_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__448__C _448_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_599_ _599_/A _599_/B vssd vssd vccd vccd _599_/X sky130_fd_sc_hd__and2_4
XFILLER_38_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__464__B _464_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_B _279_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1203_A _322_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output774_A _531_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output941_A wire1162/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput803 wire1048/X vssd vssd vccd vccd la_oenb_core[60] sky130_fd_sc_hd__buf_8
XANTENNA_wire1572_A wire1573/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput814 _567_/X vssd vssd vccd vccd la_oenb_core[70] sky130_fd_sc_hd__buf_8
Xoutput825 _577_/X vssd vssd vccd vccd la_oenb_core[80] sky130_fd_sc_hd__buf_8
Xoutput836 _587_/X vssd vssd vccd vccd la_oenb_core[90] sky130_fd_sc_hd__buf_8
Xoutput847 wire961/X vssd vssd vccd vccd mprj_ack_i_core sky130_fd_sc_hd__buf_8
Xoutput858 wire1199/X vssd vssd vccd vccd mprj_adr_o_user[19] sky130_fd_sc_hd__buf_8
XFILLER_45_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput869 wire1180/X vssd vssd vccd vccd mprj_adr_o_user[29] sky130_fd_sc_hd__buf_8
XTAP_310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[25\]_A mprj_dat_i_user[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xrebuffer12 wire1245/A vssd vssd vccd vccd rebuffer12/X sky130_fd_sc_hd__bufbuf_8
XFILLER_3_1943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_822 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__374__B _374_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[107\]_B wire1250/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_516 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1050 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[16\]_A mprj_dat_i_user[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input136_A la_iena_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_522_ _522_/A _522_/B vssd vssd vccd vccd _522_/X sky130_fd_sc_hd__and2_4
XTAP_2722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input303_A la_oenb_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__565__A _565_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_453_ _581_/A _453_/B _453_/C vssd vssd vccd vccd _453_/X sky130_fd_sc_hd__and3b_4
XTAP_2777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__284__B _284_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_384_ _512_/A _384_/B _384_/C vssd vssd vccd vccd _384_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2318 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output522_A wire1097/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__459__B _459_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1153_A _348_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3468 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput170 la_iena_mprj[19] vssd vssd vccd vccd _182_/B sky130_fd_sc_hd__clkbuf_4
Xinput181 la_iena_mprj[29] vssd vssd vccd vccd _192_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_36_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput192 la_iena_mprj[39] vssd vssd vccd vccd _202_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1320_A wire1321/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1418_A wire1419/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output891_A wire967/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[34\] la_data_out_core[34] _197_/X vssd vssd vccd vccd _017_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_36_1506 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput600 _091_/Y vssd vssd vccd vccd la_data_in_mprj[108] sky130_fd_sc_hd__buf_8
Xoutput611 _101_/Y vssd vssd vccd vccd la_data_in_mprj[118] sky130_fd_sc_hd__buf_8
Xoutput622 _159_/Y vssd vssd vccd vccd la_data_in_mprj[12] sky130_fd_sc_hd__buf_8
XFILLER_5_4119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput633 _005_/Y vssd vssd vccd vccd la_data_in_mprj[22] sky130_fd_sc_hd__buf_8
XFILLER_44_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput644 _015_/Y vssd vssd vccd vccd la_data_in_mprj[32] sky130_fd_sc_hd__buf_8
Xoutput655 _025_/Y vssd vssd vccd vccd la_data_in_mprj[42] sky130_fd_sc_hd__buf_8
Xoutput666 _035_/Y vssd vssd vccd vccd la_data_in_mprj[52] sky130_fd_sc_hd__buf_8
Xoutput677 _045_/Y vssd vssd vccd vccd la_data_in_mprj[62] sky130_fd_sc_hd__buf_8
Xoutput688 _055_/Y vssd vssd vccd vccd la_data_in_mprj[72] sky130_fd_sc_hd__buf_8
XFILLER_25_2623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput699 _065_/Y vssd vssd vccd vccd la_data_in_mprj[82] sky130_fd_sc_hd__buf_8
XFILLER_3_3120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1408 wire1409/X vssd vssd vccd vccd wire1408/X sky130_fd_sc_hd__buf_6
XFILLER_42_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1419 wire1420/X vssd vssd vccd vccd wire1419/X sky130_fd_sc_hd__buf_6
XFILLER_25_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__369__B _369_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3030 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input253_A la_iena_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3700 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input420_A mprj_cyc_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__279__B _279_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_906 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_505_ _505_/A _505_/B vssd vssd vccd vccd _505_/X sky130_fd_sc_hd__and2_4
XTAP_2552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_436_ _564_/A _436_/B _436_/C vssd vssd vccd vccd _436_/X sky130_fd_sc_hd__and3b_4
XTAP_1862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_367_ _367_/A _367_/B vssd vssd vccd vccd _367_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_298_ _298_/A _298_/B vssd vssd vccd vccd _298_/X sky130_fd_sc_hd__and2_2
XANTENNA_output472_A _477_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xrebuffer3 split13/A vssd vssd vccd vccd rebuffer3/X sky130_fd_sc_hd__bufbuf_8
XFILLER_6_840 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_884 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output737_A wire1040/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1270_A wire1270/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1368_A wire1369/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output904_A _144_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1535_A wire1535/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2542 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2794 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1702_A wire1702/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__371__C _371_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput463 _369_/X vssd vssd vccd vccd la_data_in_core[0] sky130_fd_sc_hd__buf_8
XFILLER_9_3384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3154 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput474 _379_/X vssd vssd vccd vccd la_data_in_core[10] sky130_fd_sc_hd__buf_8
Xoutput485 _380_/X vssd vssd vccd vccd la_data_in_core[11] sky130_fd_sc_hd__buf_8
XFILLER_44_3799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput496 _383_/X vssd vssd vccd vccd la_data_in_core[14] sky130_fd_sc_hd__buf_8
XFILLER_5_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1205 _320_/X vssd vssd vccd vccd wire1205/X sky130_fd_sc_hd__buf_6
Xwire1216 _314_/X vssd vssd vccd vccd wire1216/X sky130_fd_sc_hd__buf_6
Xwire1227 wire1228/X vssd vssd vccd vccd wire1227/X sky130_fd_sc_hd__buf_6
Xwire1238 _299_/X vssd vssd vccd vccd wire1238/X sky130_fd_sc_hd__buf_6
Xwire1249 _294_/X vssd vssd vccd vccd wire1249/X sky130_fd_sc_hd__buf_6
XFILLER_38_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_221_ _221_/A _221_/B vssd vssd vccd vccd _221_/X sky130_fd_sc_hd__and2_4
XFILLER_11_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_152_ _152_/A vssd vssd vccd vccd _152_/Y sky130_fd_sc_hd__inv_2
XANTENNA__562__B _562_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_083_ _083_/A vssd vssd vccd vccd _083_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_input370_A la_oenb_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input64_A la_data_out_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__456__C _456_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1116_A wire1117/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output687_A wire991/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_419_ _547_/A _419_/B _419_/C vssd vssd vccd vccd _419_/X sky130_fd_sc_hd__and3b_4
XTAP_1692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__472__B _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output854_A wire1205/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1652_A wire1652/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[108\] la_data_out_core[108] _271_/X vssd vssd vccd vccd _091_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__370__A_N _498_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__382__B _382_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[8\]_A mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1002 wire1002/A vssd vssd vccd vccd _143_/A sky130_fd_sc_hd__buf_6
XFILLER_40_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[8\]_A la_data_out_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1013 wire1013/A vssd vssd vccd vccd wire1013/X sky130_fd_sc_hd__buf_6
XFILLER_25_2283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1024 wire1024/A vssd vssd vccd vccd _129_/A sky130_fd_sc_hd__buf_8
Xwire1035 _621_/X vssd vssd vccd vccd wire1035/X sky130_fd_sc_hd__buf_6
Xwire1046 _597_/X vssd vssd vccd vccd wire1046/X sky130_fd_sc_hd__buf_6
XFILLER_38_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1057 _472_/X vssd vssd vccd vccd wire1057/X sky130_fd_sc_hd__buf_6
Xwire1068 _440_/X vssd vssd vccd vccd wire1068/X sky130_fd_sc_hd__buf_6
XFILLER_25_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1079 _425_/X vssd vssd vccd vccd wire1079/X sky130_fd_sc_hd__buf_6
XFILLER_21_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__557__B _557_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input216_A la_iena_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__573__A _573_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_204_ _204_/A _204_/B vssd vssd vccd vccd _204_/X sky130_fd_sc_hd__and2_2
XFILLER_19_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__292__B _292_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_135_ _135_/A vssd vssd vccd vccd _135_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_7_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2530 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_066_ _066_/A vssd vssd vccd vccd _066_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_7_3811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__467__B _467_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1580 wire1581/X vssd vssd vccd vccd _610_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1591 wire1591/A vssd vssd vccd vccd _602_/B sky130_fd_sc_hd__buf_6
XANTENNA_wire1233_A wire1234/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__393__A_N _521_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__377__B _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input166_A la_iena_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_2209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input333_A la_oenb_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__568__A _568_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input27_A la_data_out_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_118_ _118_/A vssd vssd vccd vccd _118_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_29_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output552_A wire1071/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_049_ _049_/A vssd vssd vccd vccd _049_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output817_A _570_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1350_A wire1351/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1448_A wire1449/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[64\] la_data_out_core[64] _227_/X vssd vssd vccd vccd _047_/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA_wire1615_A wire1615/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2514 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire970_A _130_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input283_A la_oenb_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__570__B _570_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input450_A mprj_dat_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3847 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput330 la_oenb_mprj[48] vssd vssd vccd vccd _545_/A sky130_fd_sc_hd__buf_4
XANTENNA__298__A _298_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput341 la_oenb_mprj[58] vssd vssd vccd vccd _555_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput352 la_oenb_mprj[68] vssd vssd vccd vccd _565_/A sky130_fd_sc_hd__buf_4
Xinput363 la_oenb_mprj[78] vssd vssd vccd vccd _575_/A sky130_fd_sc_hd__clkbuf_4
Xinput374 la_oenb_mprj[88] vssd vssd vccd vccd _585_/A sky130_fd_sc_hd__buf_4
XFILLER_29_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput385 la_oenb_mprj[98] vssd vssd vccd vccd _595_/A sky130_fd_sc_hd__clkbuf_4
Xinput396 mprj_adr_o_core[17] vssd vssd vccd vccd wire1400/A sky130_fd_sc_hd__buf_6
XFILLER_35_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1029_A wire1029/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_598_ _598_/A _598_/B vssd vssd vccd vccd _598_/X sky130_fd_sc_hd__and2_1
XFILLER_34_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3270 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__431__A_N _559_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output767_A _525_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__480__B _480_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1 mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput804 _558_/X vssd vssd vccd vccd la_oenb_core[61] sky130_fd_sc_hd__buf_8
XANTENNA_output934_A wire1116/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput815 _568_/X vssd vssd vccd vccd la_oenb_core[71] sky130_fd_sc_hd__buf_8
Xoutput826 _578_/X vssd vssd vccd vccd la_oenb_core[81] sky130_fd_sc_hd__buf_8
Xoutput837 _588_/X vssd vssd vccd vccd la_oenb_core[91] sky130_fd_sc_hd__buf_8
XFILLER_6_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput848 wire1226/X vssd vssd vccd vccd mprj_adr_o_user[0] sky130_fd_sc_hd__buf_8
XFILLER_28_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput859 wire1225/X vssd vssd vccd vccd mprj_adr_o_user[1] sky130_fd_sc_hd__buf_8
XTAP_300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1732_A wire1732/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__374__C _374_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__390__B _390_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1062 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input129_A la_data_out_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_521_ _521_/A _521_/B vssd vssd vccd vccd _521_/X sky130_fd_sc_hd__and2_4
XTAP_2723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__565__B _565_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_452_ _580_/A _452_/B _452_/C vssd vssd vccd vccd _452_/X sky130_fd_sc_hd__and3b_4
XFILLER_19_3888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__454__A_N _582_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_383_ _511_/A _383_/B _383_/C vssd vssd vccd vccd _383_/X sky130_fd_sc_hd__and3b_4
XFILLER_25_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3590 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input94_A la_data_out_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__581__A _581_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__459__C _459_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output515_A wire1104/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_gates\[1\]_A user_irq_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput160 la_iena_mprj[125] vssd vssd vccd vccd _288_/B sky130_fd_sc_hd__clkbuf_4
Xinput171 la_iena_mprj[1] vssd vssd vccd vccd _164_/B sky130_fd_sc_hd__buf_4
XFILLER_4_2987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput182 la_iena_mprj[2] vssd vssd vccd vccd _165_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput193 la_iena_mprj[3] vssd vssd vccd vccd _166_/B sky130_fd_sc_hd__buf_4
XANTENNA_wire1146_A wire1147/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3310 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__475__B _475_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1313_A wire1313/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output884_A wire974/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1518 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[27\] la_data_out_core[27] _190_/X vssd vssd vccd vccd _010_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_18_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1682_A wire1683/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput601 _092_/Y vssd vssd vccd vccd la_data_in_mprj[109] sky130_fd_sc_hd__buf_8
Xoutput612 _102_/Y vssd vssd vccd vccd la_data_in_mprj[119] sky130_fd_sc_hd__buf_8
Xoutput623 _160_/Y vssd vssd vccd vccd la_data_in_mprj[13] sky130_fd_sc_hd__buf_8
Xoutput634 _006_/Y vssd vssd vccd vccd la_data_in_mprj[23] sky130_fd_sc_hd__buf_8
Xoutput645 _016_/Y vssd vssd vccd vccd la_data_in_mprj[33] sky130_fd_sc_hd__buf_8
Xoutput656 _026_/Y vssd vssd vccd vccd la_data_in_mprj[43] sky130_fd_sc_hd__buf_8
Xoutput667 _036_/Y vssd vssd vccd vccd la_data_in_mprj[53] sky130_fd_sc_hd__buf_8
XFILLER_25_2613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2782 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput678 _046_/Y vssd vssd vccd vccd la_data_in_mprj[63] sky130_fd_sc_hd__buf_8
XFILLER_28_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput689 _056_/Y vssd vssd vccd vccd la_data_in_mprj[73] sky130_fd_sc_hd__buf_8
XFILLER_42_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1409 wire1409/A vssd vssd vccd vccd wire1409/X sky130_fd_sc_hd__buf_6
XFILLER_41_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__369__C _369_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__477__A_N _605_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__385__B _385_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input246_A la_iena_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input413_A mprj_adr_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__576__A _576_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_504_ _504_/A _504_/B vssd vssd vccd vccd _504_/X sky130_fd_sc_hd__and2_4
XANTENNA__295__B _295_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_435_ _563_/A _435_/B _435_/C vssd vssd vccd vccd _435_/X sky130_fd_sc_hd__and3b_4
XTAP_1863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_366_ _366_/A _366_/B vssd vssd vccd vccd _366_/X sky130_fd_sc_hd__and2_4
XFILLER_31_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_297_ _297_/A _297_/B vssd vssd vccd vccd _297_/X sky130_fd_sc_hd__and2_1
XFILLER_13_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xrebuffer4 split13/A vssd vssd vccd vccd rebuffer4/X sky130_fd_sc_hd__bufbuf_8
XFILLER_6_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output465_A _470_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_896 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output632_A _004_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[40\]_A la_data_out_core[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1430_A wire1430/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1528_A wire1528/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput464 wire1059/X vssd vssd vccd vccd la_data_in_core[100] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[31\]_A la_data_out_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput475 _479_/X vssd vssd vccd vccd la_data_in_core[110] sky130_fd_sc_hd__buf_8
XFILLER_5_3227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3166 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput486 _489_/X vssd vssd vccd vccd la_data_in_core[120] sky130_fd_sc_hd__buf_8
Xoutput497 _384_/X vssd vssd vccd vccd la_data_in_core[15] sky130_fd_sc_hd__buf_8
XFILLER_9_2673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input1_A caravel_clk vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1206 _319_/X vssd vssd vccd vccd wire1206/X sky130_fd_sc_hd__buf_6
Xwire1217 _313_/X vssd vssd vccd vccd wire1217/X sky130_fd_sc_hd__buf_6
Xwire1228 _304_/X vssd vssd vccd vccd wire1228/X sky130_fd_sc_hd__buf_6
XFILLER_41_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1239 wire1240/X vssd vssd vccd vccd wire1239/X sky130_fd_sc_hd__buf_6
XFILLER_28_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[98\]_A la_data_out_core[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_940 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_220_ _220_/A _220_/B vssd vssd vccd vccd _220_/X sky130_fd_sc_hd__and2_4
XFILLER_10_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_151_ _151_/A vssd vssd vccd vccd _151_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_3424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input196_A la_iena_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3468 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_082_ _082_/A vssd vssd vccd vccd _082_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_13_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input363_A la_oenb_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input57_A la_data_out_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[22\]_A la_data_out_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3783 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3564 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_734 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[89\]_A la_data_out_core[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_418_ _546_/A _418_/B _418_/C vssd vssd vccd vccd _418_/X sky130_fd_sc_hd__and3b_2
XTAP_1693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output582_A wire1064/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_349_ _349_/A _349_/B vssd vssd vccd vccd _349_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output847_A wire961/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1380_A wire1381/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[94\] la_data_out_core[94] _257_/X vssd vssd vccd vccd _077_/A
+ sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[13\]_A la_data_out_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2824 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1645_A wire1645/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__382__C _382_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1003 wire1004/X vssd vssd vccd vccd _142_/A sky130_fd_sc_hd__buf_6
XANTENNA_user_to_mprj_in_gates\[8\]_B _171_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1014 wire1014/A vssd vssd vccd vccd _136_/A sky130_fd_sc_hd__buf_6
XFILLER_38_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1025 wire1025/A vssd vssd vccd vccd _128_/A sky130_fd_sc_hd__buf_8
XFILLER_22_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1036 _620_/X vssd vssd vccd vccd wire1036/X sky130_fd_sc_hd__buf_6
Xwire1047 _592_/X vssd vssd vccd vccd wire1047/X sky130_fd_sc_hd__buf_6
Xwire1058 _471_/X vssd vssd vccd vccd wire1058/X sky130_fd_sc_hd__buf_6
XFILLER_21_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1069 _439_/X vssd vssd vccd vccd wire1069/X sky130_fd_sc_hd__buf_6
XFILLER_38_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input111_A la_data_out_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input209_A la_iena_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__573__B _573_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_203_ _203_/A _203_/B vssd vssd vccd vccd _203_/X sky130_fd_sc_hd__and2_2
XFILLER_12_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_134_ _134_/A vssd vssd vccd vccd _134_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_11_497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2542 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_065_ _065_/A vssd vssd vccd vccd _065_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_27_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_818 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1570 wire1571/X vssd vssd vccd vccd _615_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1581 wire1581/A vssd vssd vccd vccd wire1581/X sky130_fd_sc_hd__buf_6
XFILLER_24_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1592 wire1592/A vssd vssd vccd vccd _601_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1226_A _305_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output797_A _552_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__483__B _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_wb_dat_gates\[22\] mprj_dat_i_user[22] rebuffer7/X vssd vssd vccd vccd wire1014/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA_wire1595_A wire1595/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[120\] la_data_out_core[120] _283_/X vssd vssd vccd vccd _103_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_2_2507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__377__C _377_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__393__B _393_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input159_A la_iena_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__568__B _568_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input326_A la_oenb_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__584__A _584_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3430 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_117_ _117_/A vssd vssd vccd vccd _117_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_10_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_048_ _048_/A vssd vssd vccd vccd _048_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output545_A wire1076/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1176_A wire1177/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_2700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output712_A _077_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__478__B _478_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1343_A wire1343/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[57\] la_data_out_core[57] _220_/X vssd vssd vccd vccd _040_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_19_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1510_A wire1510/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1608_A wire1608/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[119\]_A la_data_out_core[119] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_35_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__388__B _388_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_4131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input276_A la_oenb_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_rebuffer12_A wire1245/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3467 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__383__A_N _511_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input443_A mprj_dat_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__579__A _579_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3859 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput320 la_oenb_mprj[39] vssd vssd vccd vccd _536_/A sky130_fd_sc_hd__clkbuf_4
Xinput331 la_oenb_mprj[49] vssd vssd vccd vccd _546_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput342 la_oenb_mprj[59] vssd vssd vccd vccd _556_/A sky130_fd_sc_hd__buf_4
XANTENNA__298__B _298_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput353 la_oenb_mprj[69] vssd vssd vccd vccd _566_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput364 la_oenb_mprj[79] vssd vssd vccd vccd _576_/A sky130_fd_sc_hd__buf_4
Xinput375 la_oenb_mprj[89] vssd vssd vccd vccd _586_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput386 la_oenb_mprj[99] vssd vssd vccd vccd _596_/A sky130_fd_sc_hd__clkbuf_4
Xinput397 mprj_adr_o_core[18] vssd vssd vccd vccd wire1398/A sky130_fd_sc_hd__buf_6
XFILLER_2_3594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_597_ _597_/A _597_/B vssd vssd vccd vccd _597_/X sky130_fd_sc_hd__and2_1
XFILLER_38_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output495_A _382_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output662_A _032_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__480__C _480_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2 _437_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput805 _559_/X vssd vssd vccd vccd la_oenb_core[62] sky130_fd_sc_hd__buf_8
XFILLER_6_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput816 _569_/X vssd vssd vccd vccd la_oenb_core[72] sky130_fd_sc_hd__buf_8
Xoutput827 _579_/X vssd vssd vccd vccd la_oenb_core[82] sky130_fd_sc_hd__buf_8
Xoutput838 _589_/X vssd vssd vccd vccd la_oenb_core[92] sky130_fd_sc_hd__buf_8
XANTENNA_output927_A wire1130/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput849 wire1212/X vssd vssd vccd vccd mprj_adr_o_user[10] sky130_fd_sc_hd__buf_8
XFILLER_6_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1460_A wire1461/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1558_A wire1559/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1725_A wire1725/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__390__C _390_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2578 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1074 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_520_ _520_/A _520_/B vssd vssd vccd vccd _520_/X sky130_fd_sc_hd__and2_4
XTAP_2702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_451_ _579_/A _451_/B _451_/C vssd vssd vccd vccd _451_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_382_ _510_/A _382_/B _382_/C vssd vssd vccd vccd _382_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1711 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input393_A mprj_adr_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__581__B _581_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input87_A la_data_out_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__102__A _102_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput150 la_iena_mprj[116] vssd vssd vccd vccd _279_/B sky130_fd_sc_hd__clkbuf_4
Xinput161 la_iena_mprj[126] vssd vssd vccd vccd _289_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_irq_gates\[1\]_B _292_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput172 la_iena_mprj[20] vssd vssd vccd vccd _183_/B sky130_fd_sc_hd__clkbuf_4
Xinput183 la_iena_mprj[30] vssd vssd vccd vccd _193_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_output508_A _394_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput194 la_iena_mprj[40] vssd vssd vccd vccd _203_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1139_A _355_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__475__C _475_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1306_A wire1307/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output877_A wire1218/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__491__B _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1675_A wire1675/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput602 _157_/Y vssd vssd vccd vccd la_data_in_mprj[10] sky130_fd_sc_hd__buf_8
Xoutput613 _158_/Y vssd vssd vccd vccd la_data_in_mprj[11] sky130_fd_sc_hd__buf_8
Xoutput624 _161_/Y vssd vssd vccd vccd la_data_in_mprj[14] sky130_fd_sc_hd__buf_8
XFILLER_29_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput635 _007_/Y vssd vssd vccd vccd la_data_in_mprj[24] sky130_fd_sc_hd__buf_8
Xoutput646 _017_/Y vssd vssd vccd vccd la_data_in_mprj[34] sky130_fd_sc_hd__buf_8
Xoutput657 _027_/Y vssd vssd vccd vccd la_data_in_mprj[44] sky130_fd_sc_hd__buf_8
Xoutput668 _037_/Y vssd vssd vccd vccd la_data_in_mprj[54] sky130_fd_sc_hd__buf_8
Xoutput679 _047_/Y vssd vssd vccd vccd la_data_in_mprj[64] sky130_fd_sc_hd__buf_8
XFILLER_28_1025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2794 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__012__A _012_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__385__C _385_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input141_A la_iena_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input239_A la_iena_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__421__A_N _549_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__576__B _576_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input406_A mprj_adr_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_503_ _503_/A _503_/B vssd vssd vccd vccd _503_/X sky130_fd_sc_hd__and2_4
XTAP_2532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_434_ _562_/A _434_/B _434_/C vssd vssd vccd vccd _434_/X sky130_fd_sc_hd__and3b_2
XTAP_2587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__592__A _592_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_365_ _365_/A _365_/B vssd vssd vccd vccd _365_/X sky130_fd_sc_hd__and2_4
XFILLER_9_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_296_ _296_/A _296_/B vssd vssd vccd vccd _296_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xrebuffer5 split13/A vssd vssd vccd vccd rebuffer5/X sky130_fd_sc_hd__bufbuf_8
XFILLER_26_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1089_A _415_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output625_A _162_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__486__B _486_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1423_A input3/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__007__A _007_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[1\] la_data_out_core[1] _164_/X vssd vssd vccd vccd _148_/A
+ sky130_fd_sc_hd__nand2_2
Xoutput465 _470_/X vssd vssd vccd vccd la_data_in_core[101] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[31\]_B _194_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput476 _480_/X vssd vssd vccd vccd la_data_in_core[111] sky130_fd_sc_hd__buf_8
XANTENNA__444__A_N _572_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput487 _490_/X vssd vssd vccd vccd la_data_in_core[121] sky130_fd_sc_hd__buf_8
XFILLER_5_3239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput498 _385_/X vssd vssd vccd vccd la_data_in_core[16] sky130_fd_sc_hd__buf_8
XFILLER_25_3178 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1207 _318_/X vssd vssd vccd vccd wire1207/X sky130_fd_sc_hd__buf_6
Xwire1218 _312_/X vssd vssd vccd vccd wire1218/X sky130_fd_sc_hd__buf_6
XFILLER_25_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1229 wire1230/X vssd vssd vccd vccd wire1229/X sky130_fd_sc_hd__buf_6
XFILLER_45_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__396__B _396_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[98\]_B _261_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_150_ _150_/A vssd vssd vccd vccd _150_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_081_ _081_/A vssd vssd vccd vccd _081_/Y sky130_fd_sc_hd__inv_4
XFILLER_10_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input189_A la_iena_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input356_A la_oenb_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3795 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__587__A _587_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1730 wire1731/X vssd vssd vccd vccd wire1730/X sky130_fd_sc_hd__buf_6
XFILLER_19_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[89\]_B _252_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_417_ _545_/A _417_/B _417_/C vssd vssd vccd vccd _417_/X sky130_fd_sc_hd__and3b_4
XTAP_1672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_348_ _348_/A _348_/B vssd vssd vccd vccd _348_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1004_A wire1004/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output575_A _455_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_279_ _279_/A _279_/B vssd vssd vccd vccd _279_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__467__A_N _595_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output742_A _617_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1373_A wire1373/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[13\]_B _176_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[87\] la_data_out_core[87] _250_/X vssd vssd vccd vccd _070_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_29_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1540_A wire1540/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__497__A _497_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire993_A wire993/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1004 wire1004/A vssd vssd vccd vccd wire1004/X sky130_fd_sc_hd__buf_6
Xwire1015 wire1016/X vssd vssd vccd vccd _135_/A sky130_fd_sc_hd__buf_6
XFILLER_5_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1026 wire1026/A vssd vssd vccd vccd _127_/A sky130_fd_sc_hd__buf_8
Xwire1037 _619_/X vssd vssd vccd vccd wire1037/X sky130_fd_sc_hd__buf_6
Xwire1048 _557_/X vssd vssd vccd vccd wire1048/X sky130_fd_sc_hd__buf_6
XANTENNA__200__A _200_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1059 _469_/X vssd vssd vccd vccd wire1059/X sky130_fd_sc_hd__buf_6
XFILLER_38_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input104_A la_data_out_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_202_ _202_/A _202_/B vssd vssd vccd vccd _202_/X sky130_fd_sc_hd__and2_2
XFILLER_23_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_133_ _133_/A vssd vssd vccd vccd _133_/Y sky130_fd_sc_hd__inv_6
XFILLER_32_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_064_ _064_/A vssd vssd vccd vccd _064_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_3_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__110__A _110_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1560 wire1561/X vssd vssd vccd vccd _620_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1571 wire1571/A vssd vssd vccd vccd wire1571/X sky130_fd_sc_hd__buf_6
XFILLER_21_2672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1582 wire1582/A vssd vssd vccd vccd _609_/B sky130_fd_sc_hd__buf_6
Xwire1593 wire1593/A vssd vssd vccd vccd _600_/B sky130_fd_sc_hd__buf_6
XFILLER_46_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1121_A _364_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output692_A _059_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1219_A wire1220/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__483__C _483_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[15\] mprj_dat_i_user[15] rebuffer9/X vssd vssd vccd vccd wire1024/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA_wire1490_A wire1490/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__020__A _020_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[113\] la_data_out_core[113] _276_/X vssd vssd vccd vccd _096_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_2_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__393__C _393_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input221_A la_iena_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input319_A la_oenb_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__584__B _584_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_116_ _116_/A vssd vssd vccd vccd _116_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_7_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__105__A _105_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_047_ _047_/A vssd vssd vccd vccd _047_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_2403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output538_A wire1083/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1169_A _340_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__478__C _478_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output705_A _071_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1336_A wire1337/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1390 wire1390/A vssd vssd vccd vccd wire1390/X sky130_fd_sc_hd__buf_6
XFILLER_36_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__494__B _494_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[119\]_B _282_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1503_A wire1503/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__015__A _015_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[28\]_A mprj_dat_i_user[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__388__C _388_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input171_A la_iena_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input269_A la_oenb_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__579__B _579_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[19\]_A mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input436_A mprj_dat_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput310 la_oenb_mprj[2] vssd vssd vccd vccd _499_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_20_3619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput321 la_oenb_mprj[3] vssd vssd vccd vccd _500_/A sky130_fd_sc_hd__buf_4
XFILLER_27_1465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input32_A la_data_out_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput332 la_oenb_mprj[4] vssd vssd vccd vccd _501_/A sky130_fd_sc_hd__buf_4
Xinput343 la_oenb_mprj[5] vssd vssd vccd vccd wire1422/A sky130_fd_sc_hd__buf_6
XFILLER_40_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput354 la_oenb_mprj[6] vssd vssd vccd vccd _503_/A sky130_fd_sc_hd__buf_4
Xinput365 la_oenb_mprj[7] vssd vssd vccd vccd _504_/A sky130_fd_sc_hd__buf_4
Xinput376 la_oenb_mprj[8] vssd vssd vccd vccd _505_/A sky130_fd_sc_hd__buf_4
XFILLER_40_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput387 la_oenb_mprj[9] vssd vssd vccd vccd wire1421/A sky130_fd_sc_hd__buf_6
Xinput398 mprj_adr_o_core[19] vssd vssd vccd vccd wire1395/A sky130_fd_sc_hd__buf_6
XANTENNA__595__A _595_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_596_ _596_/A _596_/B vssd vssd vccd vccd _596_/X sky130_fd_sc_hd__and2_4
XFILLER_16_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1414 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output488_A _491_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_564 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output655_A _025_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_3 _439_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput806 _560_/X vssd vssd vccd vccd la_oenb_core[63] sky130_fd_sc_hd__buf_8
Xoutput817 _570_/X vssd vssd vccd vccd la_oenb_core[73] sky130_fd_sc_hd__buf_8
XFILLER_6_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput828 _580_/X vssd vssd vccd vccd la_oenb_core[83] sky130_fd_sc_hd__buf_8
XFILLER_29_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1286_A wire1287/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput839 _590_/X vssd vssd vccd vccd la_oenb_core[93] sky130_fd_sc_hd__buf_8
XFILLER_29_2954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output822_A _575_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__489__B _489_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1453_A wire1453/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1620_A wire1620/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1718_A wire1718/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_803 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__399__B _399_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_450_ _578_/A _450_/B _450_/C vssd vssd vccd vccd _450_/X sky130_fd_sc_hd__and3b_4
XTAP_2747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_381_ _509_/A _381_/B _381_/C vssd vssd vccd vccd _381_/X sky130_fd_sc_hd__and3b_4
XFILLER_17_3570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1723 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input386_A la_oenb_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput140 la_iena_mprj[107] vssd vssd vccd vccd _270_/B sky130_fd_sc_hd__clkbuf_4
Xinput151 la_iena_mprj[117] vssd vssd vccd vccd _280_/B sky130_fd_sc_hd__clkbuf_4
Xinput162 la_iena_mprj[127] vssd vssd vccd vccd _290_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput173 la_iena_mprj[21] vssd vssd vccd vccd _184_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput184 la_iena_mprj[31] vssd vssd vccd vccd _194_/B sky130_fd_sc_hd__clkbuf_4
Xinput195 la_iena_mprj[41] vssd vssd vccd vccd _204_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_37_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1034_A _622_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_579_ _579_/A _579_/B vssd vssd vccd vccd _579_/X sky130_fd_sc_hd__and2_4
XFILLER_38_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1201_A _323_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output772_A _529_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__491__C _491_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1570_A wire1571/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput603 _093_/Y vssd vssd vccd vccd la_data_in_mprj[110] sky130_fd_sc_hd__buf_8
Xoutput614 _103_/Y vssd vssd vccd vccd la_data_in_mprj[120] sky130_fd_sc_hd__buf_8
XANTENNA_wire1668_A wire1669/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput625 _162_/Y vssd vssd vccd vccd la_data_in_mprj[15] sky130_fd_sc_hd__buf_8
XFILLER_25_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput636 _008_/Y vssd vssd vccd vccd la_data_in_mprj[25] sky130_fd_sc_hd__buf_8
XFILLER_29_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput647 _018_/Y vssd vssd vccd vccd la_data_in_mprj[35] sky130_fd_sc_hd__buf_8
XFILLER_9_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput658 _028_/Y vssd vssd vccd vccd la_data_in_mprj[45] sky130_fd_sc_hd__buf_8
Xoutput669 _038_/Y vssd vssd vccd vccd la_data_in_mprj[55] sky130_fd_sc_hd__buf_8
XFILLER_28_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__373__A_N _501_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__203__A _203_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3736 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input134_A la_iena_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_502_ _502_/A _502_/B vssd vssd vccd vccd _502_/X sky130_fd_sc_hd__and2_4
XTAP_2533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input301_A la_oenb_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_433_ _561_/A _433_/B _433_/C vssd vssd vccd vccd _433_/X sky130_fd_sc_hd__and3b_1
XTAP_1843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__592__B _592_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_364_ _364_/A _364_/B vssd vssd vccd vccd _364_/X sky130_fd_sc_hd__and2_4
XTAP_1898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_295_ _295_/A_N _295_/B vssd vssd vccd vccd _295_/X sky130_fd_sc_hd__and2b_2
XFILLER_9_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xrebuffer6 wire1248/X vssd vssd vccd vccd rebuffer6/X sky130_fd_sc_hd__bufbuf_8
XFILLER_29_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__113__A _113_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output520_A wire1099/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output618_A _107_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1151_A _349_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__486__C _486_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__396__A_N _524_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[32\] la_data_out_core[32] _195_/X vssd vssd vccd vccd _015_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_33_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_2496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput466 wire1058/X vssd vssd vccd vccd la_data_in_core[102] sky130_fd_sc_hd__buf_8
Xoutput477 _481_/X vssd vssd vccd vccd la_data_in_core[112] sky130_fd_sc_hd__buf_8
Xoutput488 _491_/X vssd vssd vccd vccd la_data_in_core[122] sky130_fd_sc_hd__buf_8
Xoutput499 _386_/X vssd vssd vccd vccd la_data_in_core[17] sky130_fd_sc_hd__buf_8
XFILLER_29_1880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1208 wire1209/X vssd vssd vccd vccd wire1208/X sky130_fd_sc_hd__buf_6
XFILLER_41_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1219 wire1220/X vssd vssd vccd vccd wire1219/X sky130_fd_sc_hd__buf_6
XFILLER_25_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_080_ _080_/A vssd vssd vccd vccd _080_/Y sky130_fd_sc_hd__inv_4
XFILLER_6_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input251_A la_iena_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input349_A la_oenb_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1720 wire1720/A vssd vssd vccd vccd _449_/B sky130_fd_sc_hd__buf_6
Xwire1731 wire1732/X vssd vssd vccd vccd wire1731/X sky130_fd_sc_hd__buf_6
XANTENNA__587__B _587_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_416_ _544_/A _416_/B _416_/C vssd vssd vccd vccd _416_/X sky130_fd_sc_hd__and3b_2
XTAP_1673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__108__A _108_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_347_ _347_/A _347_/B vssd vssd vccd vccd _347_/X sky130_fd_sc_hd__and2_4
XFILLER_30_967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_278_ _278_/A _278_/B vssd vssd vccd vccd _278_/X sky130_fd_sc_hd__and2_4
XANTENNA_output470_A _475_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output568_A _376_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1199_A wire1200/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output735_A wire1041/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1366_A wire1366/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output902_A _143_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__497__B _497_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1533_A wire1533/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1700_A wire1700/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire986_A _114_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__018__A _018_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__411__A_N _539_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1005 wire1006/X vssd vssd vccd vccd _141_/A sky130_fd_sc_hd__buf_6
XFILLER_25_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1016 wire1016/A vssd vssd vccd vccd wire1016/X sky130_fd_sc_hd__buf_6
XFILLER_38_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1027 wire1027/A vssd vssd vccd vccd _126_/A sky130_fd_sc_hd__buf_8
XFILLER_25_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1038 _616_/X vssd vssd vccd vccd wire1038/X sky130_fd_sc_hd__buf_6
Xwire1049 _555_/X vssd vssd vccd vccd wire1049/X sky130_fd_sc_hd__buf_6
XFILLER_28_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_201_ _201_/A _201_/B vssd vssd vccd vccd _201_/X sky130_fd_sc_hd__and2_2
XFILLER_15_1209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input299_A la_oenb_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_132_ _132_/A vssd vssd vccd vccd _132_/Y sky130_fd_sc_hd__inv_6
XFILLER_8_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_063_ _063_/A vssd vssd vccd vccd _063_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input62_A la_data_out_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__598__A _598_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1550 wire1550/A vssd vssd vccd vccd _164_/A sky130_fd_sc_hd__buf_6
XFILLER_8_1292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1561 wire1561/A vssd vssd vccd vccd wire1561/X sky130_fd_sc_hd__buf_6
XFILLER_1_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1572 wire1573/X vssd vssd vccd vccd _614_/B sky130_fd_sc_hd__buf_6
XFILLER_46_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1583 wire1583/A vssd vssd vccd vccd _608_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1594 wire1594/A vssd vssd vccd vccd _599_/B sky130_fd_sc_hd__buf_6
XFILLER_21_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__434__A_N _562_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1114_A wire1115/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output852_A wire1207/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1483_A wire1483/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1650_A wire1650/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__301__A _301_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[106\] la_data_out_core[106] wire1251/X vssd vssd vccd vccd
+ _089_/A sky130_fd_sc_hd__nand2_8
XFILLER_25_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__211__A _211_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3683 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input214_A la_iena_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__457__A_N _585_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_115_ _115_/A vssd vssd vccd vccd _115_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_10_2341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_046_ _046_/A vssd vssd vccd vccd _046_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__121__A _121_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output600_A _091_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1380 wire1381/X vssd vssd vccd vccd _329_/B sky130_fd_sc_hd__buf_6
Xwire1391 wire1392/X vssd vssd vccd vccd _306_/B sky130_fd_sc_hd__buf_6
XANTENNA_wire1231_A wire1232/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1329_A wire1329/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__494__C _494_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1698_A wire1698/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[28\]_B split13/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__206__A _206_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input164_A la_iena_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput300 la_oenb_mprj[20] vssd vssd vccd vccd _517_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput311 la_oenb_mprj[30] vssd vssd vccd vccd _527_/A sky130_fd_sc_hd__buf_4
Xinput322 la_oenb_mprj[40] vssd vssd vccd vccd _537_/A sky130_fd_sc_hd__clkbuf_4
Xinput333 la_oenb_mprj[50] vssd vssd vccd vccd _547_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input331_A la_oenb_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput344 la_oenb_mprj[60] vssd vssd vccd vccd _557_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input429_A mprj_dat_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput355 la_oenb_mprj[70] vssd vssd vccd vccd _567_/A sky130_fd_sc_hd__buf_4
Xinput366 la_oenb_mprj[80] vssd vssd vccd vccd _577_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input25_A la_data_out_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput377 la_oenb_mprj[90] vssd vssd vccd vccd _587_/A sky130_fd_sc_hd__clkbuf_4
Xinput388 mprj_adr_o_core[0] vssd vssd vccd vccd wire1420/A sky130_fd_sc_hd__buf_6
XFILLER_40_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput399 mprj_adr_o_core[1] vssd vssd vccd vccd wire1393/A sky130_fd_sc_hd__buf_6
XFILLER_21_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__595__B _595_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_595_ _595_/A _595_/B vssd vssd vccd vccd _595_/X sky130_fd_sc_hd__and2_4
XFILLER_16_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__116__A _116_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_4 _439_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput807 _561_/X vssd vssd vccd vccd la_oenb_core[64] sky130_fd_sc_hd__buf_8
Xoutput818 _571_/X vssd vssd vccd vccd la_oenb_core[74] sky130_fd_sc_hd__buf_8
XANTENNA_output550_A _432_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[70\]_A la_data_out_core[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput829 _581_/X vssd vssd vccd vccd la_oenb_core[84] sky130_fd_sc_hd__buf_8
XFILLER_6_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_029_ _029_/A vssd vssd vccd vccd _029_/Y sky130_fd_sc_hd__inv_2
XANTENNA_wire1181_A _334_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1279_A wire1279/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3463 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__489__C _489_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output815_A _568_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1446_A wire1447/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[62\] la_data_out_core[62] _225_/X vssd vssd vccd vccd _045_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_39_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1613_A wire1613/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_826 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[61\]_A la_data_out_core[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__399__C _399_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_380_ _508_/A _380_/B _380_/C vssd vssd vccd vccd _380_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1779 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input281_A la_oenb_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input379_A la_oenb_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[52\]_A la_data_out_core[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput130 la_data_out_mprj[99] vssd vssd vccd vccd _468_/C sky130_fd_sc_hd__clkbuf_4
Xinput141 la_iena_mprj[108] vssd vssd vccd vccd _271_/B sky130_fd_sc_hd__clkbuf_4
Xinput152 la_iena_mprj[118] vssd vssd vccd vccd _281_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput163 la_iena_mprj[12] vssd vssd vccd vccd _175_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput174 la_iena_mprj[22] vssd vssd vccd vccd _185_/B sky130_fd_sc_hd__clkbuf_4
Xinput185 la_iena_mprj[32] vssd vssd vccd vccd _195_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput196 la_iena_mprj[42] vssd vssd vccd vccd _205_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_578_ _578_/A _578_/B vssd vssd vccd vccd _578_/X sky130_fd_sc_hd__and2_4
XFILLER_31_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1027_A wire1027/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output598_A _089_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output765_A wire1053/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1396_A wire1397/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output932_A wire1120/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput604 _094_/Y vssd vssd vccd vccd la_data_in_mprj[111] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[43\]_A la_data_out_core[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput615 _104_/Y vssd vssd vccd vccd la_data_in_mprj[121] sky130_fd_sc_hd__buf_8
XFILLER_44_3929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput626 _163_/Y vssd vssd vccd vccd la_data_in_mprj[16] sky130_fd_sc_hd__buf_8
XFILLER_25_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput637 _009_/Y vssd vssd vccd vccd la_data_in_mprj[26] sky130_fd_sc_hd__buf_8
XANTENNA_wire1563_A wire1563/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput648 _019_/Y vssd vssd vccd vccd la_data_in_mprj[36] sky130_fd_sc_hd__buf_8
XFILLER_28_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput659 _029_/Y vssd vssd vccd vccd la_data_in_mprj[46] sky130_fd_sc_hd__buf_8
XFILLER_29_2763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1730_A wire1731/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
.ends

