* NGSPICE file created from digital_pll.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_2 abstract view
.subckt sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_8 abstract view
.subckt sky130_fd_sc_hd__einvn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_4 abstract view
.subckt sky130_fd_sc_hd__einvn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_1 abstract view
.subckt sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

.subckt digital_pll VGND VPWR clockp[0] clockp[1] dco div[0] div[1] div[2] div[3]
+ div[4] enable ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12] ext_trim[13] ext_trim[14]
+ ext_trim[15] ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19] ext_trim[1] ext_trim[20]
+ ext_trim[21] ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25] ext_trim[2] ext_trim[3]
+ ext_trim[4] ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8] ext_trim[9] osc resetb
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__338__A1 ext_trim[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_363_ _312_/X ext_trim[25] dco VGND VGND VPWR VPWR _363_/X sky130_fd_sc_hd__mux2_1
X_294_ _305_/A _376_/Q _378_/Q _375_/Q _292_/X VGND VGND VPWR VPWR _294_/X sky130_fd_sc_hd__o41a_2
Xringosc.dstage\[1\].id.delayint0 ringosc.dstage\[1\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XANTENNA__214__A div[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_346_ _298_/X ext_trim[7] dco VGND VGND VPWR VPWR _346_/X sky130_fd_sc_hd__mux2_1
X_277_ _368_/Q _367_/Q _369_/Q _370_/Q VGND VGND VPWR VPWR _277_/X sky130_fd_sc_hd__a31o_2
X_200_ _369_/Q _384_/Q VGND VGND VPWR VPWR _200_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__209__A div[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_329_ _335_/A VGND VGND VPWR VPWR _329_/X sky130_fd_sc_hd__buf_1
Xringosc.dstage\[11\].id.delayen1 ringosc.dstage\[11\].id.delayen1/A _339_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[11\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[10\].id.delayenb0 ringosc.dstage\[10\].id.delayenb1/A _340_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XFILLER_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[9\].id.delayenb0 ringosc.dstage\[9\].id.delayenb1/A _342_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[9\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_362_ _290_/X ext_trim[12] dco VGND VGND VPWR VPWR _362_/X sky130_fd_sc_hd__mux2_1
X_293_ _305_/A _376_/Q _378_/Q _305_/C _292_/X VGND VGND VPWR VPWR _293_/X sky130_fd_sc_hd__o41a_2
XANTENNA__320__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_276_ _371_/Q _275_/Y _187_/Y VGND VGND VPWR VPWR _371_/D sky130_fd_sc_hd__o21a_2
X_345_ _301_/X ext_trim[21] dco VGND VGND VPWR VPWR _345_/X sky130_fd_sc_hd__mux2_1
XANTENNA__315__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_328_ _335_/A VGND VGND VPWR VPWR _328_/X sky130_fd_sc_hd__buf_1
X_259_ _264_/A _264_/B VGND VGND VPWR VPWR _259_/X sky130_fd_sc_hd__or2_2
XFILLER_20_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[10\].id.delayenb1 ringosc.dstage\[10\].id.delayenb1/A _341_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[9\].id.delayenb1 ringosc.dstage\[9\].id.delayenb1/A _343_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[9\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XANTENNA__323__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__318__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_361_ _299_/X ext_trim[13] dco VGND VGND VPWR VPWR _361_/X sky130_fd_sc_hd__mux2_1
X_292_ _378_/Q _310_/C _296_/B VGND VGND VPWR VPWR _292_/X sky130_fd_sc_hd__o21a_2
X_275_ _275_/A VGND VGND VPWR VPWR _275_/Y sky130_fd_sc_hd__inv_2
X_344_ _289_/X ext_trim[8] dco VGND VGND VPWR VPWR _344_/X sky130_fd_sc_hd__mux2_1
XANTENNA__331__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[4\].id.delayen0 ringosc.dstage\[4\].id.delayen0/A _352_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_327_ _335_/A VGND VGND VPWR VPWR _327_/X sky130_fd_sc_hd__buf_1
XANTENNA__326__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_189_ enable resetb VGND VGND VPWR VPWR _190_/B sky130_fd_sc_hd__nand2_2
X_258_ _309_/A _273_/B _257_/X VGND VGND VPWR VPWR _378_/D sky130_fd_sc_hd__o21ai_2
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__359__A1 ext_trim[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[5\].id.delayenb0 ringosc.dstage\[5\].id.delayenb1/A _350_/X VGND
+ VGND VPWR VPWR ringosc.ibufp10/A sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[10\].id.delaybuf0 ringosc.dstage\[9\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[9\].id.delaybuf0 ringosc.dstage\[8\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_360_ _240_/C ext_trim[0] dco VGND VGND VPWR VPWR _360_/X sky130_fd_sc_hd__mux2_1
X_291_ _378_/Q _310_/C _296_/A _296_/B VGND VGND VPWR VPWR _291_/X sky130_fd_sc_hd__o31a_2
XANTENNA__329__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_274_ _274_/A _282_/B _274_/C _274_/D VGND VGND VPWR VPWR _275_/A sky130_fd_sc_hd__or4_2
X_343_ _304_/X ext_trim[22] dco VGND VGND VPWR VPWR _343_/X sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[4\].id.delayen1 ringosc.dstage\[4\].id.delayen1/A _353_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_326_ _335_/A VGND VGND VPWR VPWR _326_/X sky130_fd_sc_hd__buf_1
X_188_ _386_/Q _187_/Y _371_/Q _233_/B VGND VGND VPWR VPWR _386_/D sky130_fd_sc_hd__a22o_2
X_257_ _254_/Y _256_/A _254_/A _256_/Y _243_/Y VGND VGND VPWR VPWR _257_/X sky130_fd_sc_hd__a221o_2
XFILLER_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_309_ _309_/A _309_/B VGND VGND VPWR VPWR _309_/Y sky130_fd_sc_hd__nor2_2
XFILLER_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[5\].id.delayenb1 ringosc.dstage\[5\].id.delayenb1/A _351_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[5\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[10\].id.delaybuf1 ringosc.dstage\[10\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[9\].id.delaybuf1 ringosc.dstage\[9\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_290_ _378_/Q _310_/C _375_/Q _296_/B VGND VGND VPWR VPWR _290_/X sky130_fd_sc_hd__o31a_2
X_273_ _372_/Q _273_/B VGND VGND VPWR VPWR _372_/D sky130_fd_sc_hd__xor2_1
X_342_ _293_/X ext_trim[9] dco VGND VGND VPWR VPWR _342_/X sky130_fd_sc_hd__mux2_1
X_187_ _233_/B VGND VGND VPWR VPWR _187_/Y sky130_fd_sc_hd__inv_2
X_256_ _256_/A VGND VGND VPWR VPWR _256_/Y sky130_fd_sc_hd__inv_2
X_325_ _335_/A VGND VGND VPWR VPWR _325_/X sky130_fd_sc_hd__buf_1
X_308_ _268_/A _374_/Q _309_/A _310_/C _304_/X VGND VGND VPWR VPWR _308_/X sky130_fd_sc_hd__o41a_2
X_239_ _378_/Q _239_/B VGND VGND VPWR VPWR _240_/C sky130_fd_sc_hd__or2_2
XFILLER_20_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[5\].id.delaybuf0 ringosc.dstage\[4\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[1\].id.delayenb0 ringosc.dstage\[1\].id.delayenb1/A _358_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[1\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
X_341_ _334_/X ext_trim[23] dco VGND VGND VPWR VPWR _341_/X sky130_fd_sc_hd__mux2_1
X_272_ _231_/A _273_/B _243_/Y _271_/X VGND VGND VPWR VPWR _373_/D sky130_fd_sc_hd__o22ai_2
XFILLER_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__340__A1 ext_trim[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[8\].id.delayint0 ringosc.dstage\[8\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_186_ _366_/D _366_/Q VGND VGND VPWR VPWR _233_/B sky130_fd_sc_hd__xor2_1
X_255_ _378_/Q _255_/B VGND VGND VPWR VPWR _256_/A sky130_fd_sc_hd__xor2_1
X_324_ _335_/A VGND VGND VPWR VPWR _324_/X sky130_fd_sc_hd__buf_1
X_169_ _386_/Q VGND VGND VPWR VPWR _219_/B sky130_fd_sc_hd__inv_2
X_238_ _305_/C _310_/B VGND VGND VPWR VPWR _239_/B sky130_fd_sc_hd__or2_2
X_307_ _337_/X _307_/B VGND VGND VPWR VPWR _307_/X sky130_fd_sc_hd__and2_2
XFILLER_19_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[5\].id.delaybuf1 ringosc.dstage\[5\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[1\].id.delayenb1 ringosc.dstage\[1\].id.delayenb1/A _359_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[1\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_340_ _296_/X ext_trim[10] dco VGND VGND VPWR VPWR _340_/X sky130_fd_sc_hd__mux2_1
X_271_ _372_/Q _271_/B VGND VGND VPWR VPWR _271_/X sky130_fd_sc_hd__xor2_1
Xringosc.dstage\[1\].id.delayen0 ringosc.dstage\[1\].id.delayen0/A _358_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
X_185_ div[0] VGND VGND VPWR VPWR _185_/Y sky130_fd_sc_hd__inv_2
X_323_ _335_/A VGND VGND VPWR VPWR _323_/X sky130_fd_sc_hd__buf_1
X_254_ _254_/A VGND VGND VPWR VPWR _254_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_168_ _371_/Q VGND VGND VPWR VPWR _168_/Y sky130_fd_sc_hd__inv_2
X_306_ _309_/A _310_/C _268_/A _305_/X _304_/X VGND VGND VPWR VPWR _306_/X sky130_fd_sc_hd__o311a_2
X_237_ _310_/B VGND VGND VPWR VPWR _309_/B sky130_fd_sc_hd__inv_2
XFILLER_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_270_ _243_/Y _269_/X _374_/Q _243_/Y VGND VGND VPWR VPWR _374_/D sky130_fd_sc_hd__a2bb2o_2
XFILLER_4_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[1\].id.delayen1 ringosc.dstage\[1\].id.delayen1/A _359_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_3_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[1\].id.delaybuf0 ringosc.dstage\[0\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_322_ _335_/A VGND VGND VPWR VPWR _322_/X sky130_fd_sc_hd__buf_1
Xringosc.dstage\[4\].id.delayint0 ringosc.dstage\[4\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_184_ _372_/Q VGND VGND VPWR VPWR _231_/B sky130_fd_sc_hd__inv_2
X_253_ _264_/B _252_/A _264_/A _250_/B _309_/B VGND VGND VPWR VPWR _254_/A sky130_fd_sc_hd__o32a_2
X_236_ _377_/Q _376_/Q VGND VGND VPWR VPWR _310_/B sky130_fd_sc_hd__or2_2
X_305_ _305_/A _376_/Q _305_/C _309_/A VGND VGND VPWR VPWR _305_/X sky130_fd_sc_hd__or4_2
XFILLER_19_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_219_ _371_/Q _219_/B VGND VGND VPWR VPWR _221_/A sky130_fd_sc_hd__xor2_1
Xringosc.dstage\[9\].id.delayen0 ringosc.dstage\[9\].id.delayen0/A _342_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__361__A1 ext_trim[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__352__A1 ext_trim[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__343__A1 ext_trim[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[1\].id.delaybuf1 ringosc.dstage\[1\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_321_ _335_/A VGND VGND VPWR VPWR _321_/X sky130_fd_sc_hd__buf_1
X_183_ _373_/Q VGND VGND VPWR VPWR _231_/A sky130_fd_sc_hd__inv_2
X_252_ _252_/A VGND VGND VPWR VPWR _252_/Y sky130_fd_sc_hd__inv_2
XANTENNA__225__B1 div[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_235_ _305_/C VGND VGND VPWR VPWR _246_/B sky130_fd_sc_hd__inv_2
X_304_ _375_/Q _247_/A _310_/C _309_/A _303_/X VGND VGND VPWR VPWR _304_/X sky130_fd_sc_hd__o41a_2
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_218_ div[1] _214_/B _217_/X VGND VGND VPWR VPWR _218_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__364__D osc VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[9\].id.delayen1 ringosc.dstage\[9\].id.delayen1/A _343_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__341__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_182_ _374_/Q VGND VGND VPWR VPWR _247_/A sky130_fd_sc_hd__inv_2
X_251_ _305_/A _255_/B VGND VGND VPWR VPWR _252_/A sky130_fd_sc_hd__xor2_1
X_320_ _335_/A VGND VGND VPWR VPWR _320_/X sky130_fd_sc_hd__buf_1
X_234_ _375_/Q _374_/Q VGND VGND VPWR VPWR _305_/C sky130_fd_sc_hd__or2_2
X_303_ _309_/A _310_/B _268_/A _302_/X _301_/X VGND VGND VPWR VPWR _303_/X sky130_fd_sc_hd__o311a_2
Xringosc.dstage\[0\].id.delayint0 ringosc.dstage\[0\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.iss.reseten0 ringosc.iss.const1/HI _190_/B VGND VGND VPWR VPWR ringosc.ibufp00/A
+ sky130_fd_sc_hd__einvp_1
X_217_ div[1] _214_/B div[0] _216_/Y _214_/Y VGND VGND VPWR VPWR _217_/X sky130_fd_sc_hd__o221a_2
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__344__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__339__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[8\].id.delayenb0 ringosc.dstage\[8\].id.delayenb1/A _344_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[8\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__352__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_250_ _376_/Q _250_/B VGND VGND VPWR VPWR _264_/B sky130_fd_sc_hd__xor2_1
X_181_ _375_/Q VGND VGND VPWR VPWR _268_/A sky130_fd_sc_hd__inv_2
X_379_ _336_/A _379_/D _318_/X VGND VGND VPWR VPWR _379_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__347__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_302_ _305_/C _310_/C _309_/A VGND VGND VPWR VPWR _302_/X sky130_fd_sc_hd__or3_2
X_233_ _380_/Q _233_/B _381_/Q _379_/Q VGND VGND VPWR VPWR _233_/X sky130_fd_sc_hd__and4_2
XFILLER_19_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_216_ _216_/A VGND VGND VPWR VPWR _216_/Y sky130_fd_sc_hd__inv_2
Xringosc.iss.delayint0 ringosc.iss.delayen1/Z VGND VGND VPWR VPWR ringosc.iss.delayen0/A
+ sky130_fd_sc_hd__clkinv_1
XANTENNA__360__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__355__A1 ext_trim[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__346__A1 ext_trim[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__355__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[8\].id.delayenb1 ringosc.dstage\[8\].id.delayenb1/A _345_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[8\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_180_ _376_/Q VGND VGND VPWR VPWR _288_/B sky130_fd_sc_hd__inv_2
X_378_ _336_/A _378_/D _319_/X VGND VGND VPWR VPWR _378_/Q sky130_fd_sc_hd__dfrtp_2
X_232_ _185_/Y _216_/A _217_/X _212_/A _223_/Y VGND VGND VPWR VPWR _232_/Y sky130_fd_sc_hd__o2111ai_2
XANTENNA__363__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_301_ _375_/Q _247_/A _310_/B _378_/Q _239_/B VGND VGND VPWR VPWR _301_/X sky130_fd_sc_hd__o311a_2
XFILLER_19_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__358__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[6\].id.delayen0 ringosc.dstage\[6\].id.delayen0/A _348_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
X_215_ _282_/B _215_/B VGND VGND VPWR VPWR _216_/A sky130_fd_sc_hd__xor2_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_377_ _336_/A _377_/D _320_/X VGND VGND VPWR VPWR _377_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[4\].id.delayenb0 ringosc.dstage\[4\].id.delayenb1/A _352_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[4\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[8\].id.delaybuf0 ringosc.dstage\[7\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_231_ _231_/A _231_/B _300_/B VGND VGND VPWR VPWR _231_/X sky130_fd_sc_hd__or3_2
X_300_ _309_/A _300_/B VGND VGND VPWR VPWR _307_/B sky130_fd_sc_hd__nand2_2
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[10\].id.delayen0 ringosc.dstage\[10\].id.delayen0/A _340_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
Xringosc.dstage\[6\].id.delayen1 ringosc.dstage\[6\].id.delayen1/A _349_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_214_ div[1] _214_/B VGND VGND VPWR VPWR _214_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__313__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__223__A div[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__321__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[4\].id.delayenb1 ringosc.dstage\[4\].id.delayenb1/A _353_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[4\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_376_ _336_/A _376_/D _321_/X VGND VGND VPWR VPWR _376_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[8\].id.delaybuf1 ringosc.dstage\[8\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_230_ _305_/A _288_/B _230_/C VGND VGND VPWR VPWR _300_/B sky130_fd_sc_hd__or3_2
XANTENNA__316__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_359_ _306_/X ext_trim[14] dco VGND VGND VPWR VPWR _359_/X sky130_fd_sc_hd__mux2_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[10\].id.delayen1 ringosc.dstage\[10\].id.delayen1/A _341_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_10_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_213_ _201_/X _202_/X _201_/X _202_/X VGND VGND VPWR VPWR _214_/B sky130_fd_sc_hd__a2bb2o_2
XANTENNA__358__A1 ext_trim[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__349__A1 ext_trim[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__324__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__319__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_375_ _336_/A _375_/D _322_/X VGND VGND VPWR VPWR _375_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__332__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_358_ _297_/X ext_trim[1] dco VGND VGND VPWR VPWR _358_/X sky130_fd_sc_hd__mux2_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__327__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[4\].id.delaybuf0 ringosc.dstage\[3\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_289_ _305_/C _310_/C _378_/Q _296_/B VGND VGND VPWR VPWR _289_/X sky130_fd_sc_hd__o31a_2
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_212_ _212_/A VGND VGND VPWR VPWR _212_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[7\].id.delayint0 ringosc.dstage\[7\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[0\].id.delayenb0 ringosc.dstage\[0\].id.delayenb1/A _360_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[0\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__335__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_374_ _336_/A _374_/D _323_/X VGND VGND VPWR VPWR _374_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[3\].id.delayen0 ringosc.dstage\[3\].id.delayen0/A _354_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_357_ _303_/X ext_trim[15] dco VGND VGND VPWR VPWR _357_/X sky130_fd_sc_hd__mux2_1
X_288_ _377_/Q _288_/B VGND VGND VPWR VPWR _310_/C sky130_fd_sc_hd__or2_2
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[4\].id.delaybuf1 ringosc.dstage\[4\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_211_ div[2] _207_/X _210_/A _208_/Y VGND VGND VPWR VPWR _212_/A sky130_fd_sc_hd__o211a_2
Xringosc.dstage\[0\].id.delayenb1 ringosc.dstage\[0\].id.delayenb1/A _361_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[0\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.iss.delayenb0 ringosc.iss.delayenb1/A ringosc.iss.ctrlen0/X VGND VGND VPWR
+ VPWR ringosc.ibufp00/A sky130_fd_sc_hd__einvn_8
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_373_ _336_/A _373_/D _324_/X VGND VGND VPWR VPWR _373_/Q sky130_fd_sc_hd__dfrtp_2
X_287_ _375_/Q _296_/B VGND VGND VPWR VPWR _287_/X sky130_fd_sc_hd__or2_2
X_356_ _292_/X ext_trim[2] dco VGND VGND VPWR VPWR _356_/X sky130_fd_sc_hd__mux2_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[3\].id.delayen1 ringosc.dstage\[3\].id.delayen1/A _355_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_210_ _210_/A VGND VGND VPWR VPWR _210_/Y sky130_fd_sc_hd__inv_2
X_339_ _310_/X ext_trim[24] dco VGND VGND VPWR VPWR _339_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.iss.delayenb1 ringosc.iss.delayenb1/A _363_/X VGND VGND VPWR VPWR ringosc.iss.delayen1/Z
+ sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[0\].id.delaybuf0 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.dstage\[0\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[3\].id.delayint0 ringosc.dstage\[3\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_372_ _336_/A _372_/D _325_/X VGND VGND VPWR VPWR _372_/Q sky130_fd_sc_hd__dfrtp_2
X_286_ _378_/Q _310_/B VGND VGND VPWR VPWR _296_/B sky130_fd_sc_hd__or2_2
X_355_ _307_/X ext_trim[16] dco VGND VGND VPWR VPWR _355_/X sky130_fd_sc_hd__mux2_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_338_ _295_/X ext_trim[11] dco VGND VGND VPWR VPWR _338_/X sky130_fd_sc_hd__mux2_1
X_269_ _269_/A _269_/B VGND VGND VPWR VPWR _269_/X sky130_fd_sc_hd__xor2_1
Xringosc.dstage\[0\].id.delaybuf1 ringosc.dstage\[0\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__190__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.iss.delaybuf0 ringosc.iss.delayenb1/A VGND VGND VPWR VPWR ringosc.iss.delayen1/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__185__A div[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_371_ _336_/A _371_/D _326_/X VGND VGND VPWR VPWR _371_/Q sky130_fd_sc_hd__dfrtp_2
X_354_ _296_/B ext_trim[3] dco VGND VGND VPWR VPWR _354_/X sky130_fd_sc_hd__mux2_1
X_285_ _371_/Q _275_/Y _282_/B _233_/B VGND VGND VPWR VPWR _367_/D sky130_fd_sc_hd__a211o_2
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_199_ _370_/Q _199_/B VGND VGND VPWR VPWR _199_/X sky130_fd_sc_hd__xor2_1
XFILLER_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_268_ _268_/A _268_/B VGND VGND VPWR VPWR _375_/D sky130_fd_sc_hd__xor2_1
X_337_ _300_/B _239_/B _378_/Q VGND VGND VPWR VPWR _337_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__360__A1 ext_trim[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__351__A1 ext_trim[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__342__A1 ext_trim[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__385__RESET_B _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_370_ _336_/A _370_/D _327_/X VGND VGND VPWR VPWR _370_/Q sky130_fd_sc_hd__dfrtp_2
X_284_ _284_/A VGND VGND VPWR VPWR _368_/D sky130_fd_sc_hd__inv_2
Xringosc.dstage\[0\].id.delayen0 ringosc.dstage\[0\].id.delayen0/A _360_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
X_353_ _308_/X ext_trim[17] dco VGND VGND VPWR VPWR _353_/X sky130_fd_sc_hd__mux2_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_198_ _370_/Q _385_/Q VGND VGND VPWR VPWR _198_/Y sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[7\].id.delayenb0 ringosc.dstage\[7\].id.delayenb1/A _346_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[7\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
X_336_ _336_/A VGND VGND VPWR VPWR clockp[0] sky130_fd_sc_hd__buf_2
X_267_ _247_/A _250_/B _273_/B _266_/X VGND VGND VPWR VPWR _268_/B sky130_fd_sc_hd__o211ai_2
X_319_ _335_/A VGND VGND VPWR VPWR _319_/X sky130_fd_sc_hd__buf_1
Xringosc.dstage\[0\].id.delayen1 ringosc.dstage\[0\].id.delayen1/A _361_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_352_ _294_/X ext_trim[4] dco VGND VGND VPWR VPWR _352_/X sky130_fd_sc_hd__mux2_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ _168_/Y _275_/A _233_/B _233_/B _282_/X VGND VGND VPWR VPWR _284_/A sky130_fd_sc_hd__o32a_2
XFILLER_14_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[7\].id.delayenb1 ringosc.dstage\[7\].id.delayenb1/A _347_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[7\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_266_ _374_/Q _255_/B _269_/A VGND VGND VPWR VPWR _266_/X sky130_fd_sc_hd__mux2_1
X_197_ _379_/Q _233_/B VGND VGND VPWR VPWR _379_/D sky130_fd_sc_hd__or2_2
X_335_ _335_/A VGND VGND VPWR VPWR _335_/X sky130_fd_sc_hd__buf_1
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_249_ _246_/Y _248_/Y _269_/A _250_/B _246_/B VGND VGND VPWR VPWR _264_/A sky130_fd_sc_hd__o32a_2
X_318_ _335_/A VGND VGND VPWR VPWR _318_/X sky130_fd_sc_hd__buf_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[8\].id.delayen0 ringosc.dstage\[8\].id.delayen0/A _344_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[8\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XANTENNA__342__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_282_ _368_/Q _282_/B VGND VGND VPWR VPWR _282_/X sky130_fd_sc_hd__xor2_1
XFILLER_14_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_351_ _309_/Y ext_trim[18] dco VGND VGND VPWR VPWR _351_/X sky130_fd_sc_hd__mux2_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_334_ _378_/Q VGND VGND VPWR VPWR _334_/X sky130_fd_sc_hd__buf_1
XANTENNA__363__A1 ext_trim[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_265_ _273_/B _259_/X _264_/Y _376_/Q _243_/Y VGND VGND VPWR VPWR _376_/D sky130_fd_sc_hd__a32o_2
X_196_ _380_/Q _187_/Y _379_/Q _233_/B VGND VGND VPWR VPWR _380_/D sky130_fd_sc_hd__a22o_2
XANTENNA__354__A1 ext_trim[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__350__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_248_ _269_/B VGND VGND VPWR VPWR _248_/Y sky130_fd_sc_hd__inv_2
XANTENNA__345__A1 ext_trim[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_179_ _377_/Q VGND VGND VPWR VPWR _305_/A sky130_fd_sc_hd__inv_2
X_317_ _335_/A VGND VGND VPWR VPWR _317_/X sky130_fd_sc_hd__buf_1
Xringosc.dstage\[3\].id.delayenb0 ringosc.dstage\[3\].id.delayenb1/A _354_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[3\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[7\].id.delaybuf0 ringosc.dstage\[6\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[11\].id.delayint0 ringosc.dstage\[11\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XANTENNA__345__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[8\].id.delayen1 ringosc.dstage\[8\].id.delayen1/A _345_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[8\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_350_ _291_/X ext_trim[5] dco VGND VGND VPWR VPWR _350_/X sky130_fd_sc_hd__mux2_1
X_281_ _371_/Q _275_/Y _187_/Y _280_/X VGND VGND VPWR VPWR _369_/D sky130_fd_sc_hd__a31o_2
XANTENNA__353__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__348__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_333_ _335_/A VGND VGND VPWR VPWR _333_/X sky130_fd_sc_hd__buf_1
X_264_ _264_/A _264_/B VGND VGND VPWR VPWR _264_/Y sky130_fd_sc_hd__nand2_2
X_195_ _380_/Q _233_/B _381_/Q _187_/Y VGND VGND VPWR VPWR _381_/D sky130_fd_sc_hd__a22o_2
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_247_ _247_/A _250_/B VGND VGND VPWR VPWR _269_/B sky130_fd_sc_hd__xor2_1
X_316_ _335_/A VGND VGND VPWR VPWR _316_/X sky130_fd_sc_hd__buf_1
Xringosc.dstage\[3\].id.delayenb1 ringosc.dstage\[3\].id.delayenb1/A _355_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[3\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[7\].id.delaybuf1 ringosc.dstage\[7\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_178_ _378_/Q VGND VGND VPWR VPWR _309_/A sky130_fd_sc_hd__inv_2
XANTENNA__361__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__356__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__218__A1 div[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_280_ _274_/A _282_/B _274_/C _187_/Y _279_/Y VGND VGND VPWR VPWR _280_/X sky130_fd_sc_hd__o311a_2
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_194_ _382_/Q _187_/Y _367_/Q _233_/B VGND VGND VPWR VPWR _382_/D sky130_fd_sc_hd__a22o_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_332_ _335_/A VGND VGND VPWR VPWR _332_/X sky130_fd_sc_hd__buf_1
X_263_ _305_/A _273_/B _262_/X VGND VGND VPWR VPWR _377_/D sky130_fd_sc_hd__o21ai_2
XANTENNA__359__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_177_ _382_/Q VGND VGND VPWR VPWR _215_/B sky130_fd_sc_hd__inv_2
X_315_ _335_/A VGND VGND VPWR VPWR _315_/X sky130_fd_sc_hd__buf_1
X_246_ _296_/A _246_/B VGND VGND VPWR VPWR _246_/Y sky130_fd_sc_hd__nor2_2
XFILLER_22_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_229_ _230_/C VGND VGND VPWR VPWR _296_/A sky130_fd_sc_hd__inv_2
Xringosc.dstage\[3\].id.delaybuf0 ringosc.dstage\[2\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[6\].id.delayint0 ringosc.dstage\[6\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_17_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.ibufp10 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.ibufp11/A sky130_fd_sc_hd__clkinv_2
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_193_ _383_/Q _187_/Y _368_/Q _233_/B VGND VGND VPWR VPWR _383_/D sky130_fd_sc_hd__a22o_2
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ _335_/A VGND VGND VPWR VPWR _331_/X sky130_fd_sc_hd__buf_1
X_262_ _252_/Y _261_/A _252_/A _261_/Y _243_/Y VGND VGND VPWR VPWR _262_/X sky130_fd_sc_hd__a221o_2
XANTENNA__357__A1 ext_trim[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__348__A1 ext_trim[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__339__A1 ext_trim[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_176_ _367_/Q VGND VGND VPWR VPWR _282_/B sky130_fd_sc_hd__inv_2
X_314_ _335_/A VGND VGND VPWR VPWR _314_/X sky130_fd_sc_hd__buf_1
X_245_ _231_/A _250_/B _231_/B _271_/B VGND VGND VPWR VPWR _269_/A sky130_fd_sc_hd__o22a_2
Xringosc.dstage\[5\].id.delayen0 ringosc.dstage\[5\].id.delayen0/A _350_/X VGND VGND
+ VPWR VPWR ringosc.ibufp10/A sky130_fd_sc_hd__einvp_2
XANTENNA__314__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[3\].id.delaybuf1 ringosc.dstage\[3\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_228_ _268_/A _247_/A VGND VGND VPWR VPWR _230_/C sky130_fd_sc_hd__or2_2
XANTENNA__322__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.ibufp11 ringosc.ibufp11/A VGND VGND VPWR VPWR clockp[1] sky130_fd_sc_hd__clkinv_8
Xringosc.ibufp00 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.ibufp01/A sky130_fd_sc_hd__clkinv_2
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__317__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_192_ _384_/Q _187_/Y _369_/Q _233_/B VGND VGND VPWR VPWR _384_/D sky130_fd_sc_hd__a22o_2
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ _335_/A VGND VGND VPWR VPWR _330_/X sky130_fd_sc_hd__buf_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ _261_/A VGND VGND VPWR VPWR _261_/Y sky130_fd_sc_hd__inv_2
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_313_ _335_/A VGND VGND VPWR VPWR _313_/X sky130_fd_sc_hd__buf_1
X_175_ _383_/Q VGND VGND VPWR VPWR _202_/B sky130_fd_sc_hd__inv_2
X_244_ _373_/Q _250_/B VGND VGND VPWR VPWR _271_/B sky130_fd_sc_hd__xor2_1
Xringosc.dstage\[5\].id.delayen1 ringosc.dstage\[5\].id.delayen1/A _351_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[5\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XANTENNA__330__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_227_ _250_/B VGND VGND VPWR VPWR _255_/B sky130_fd_sc_hd__inv_2
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__325__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[2\].id.delayint0 ringosc.dstage\[2\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_14_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.ibufp01 ringosc.ibufp01/A VGND VGND VPWR VPWR _336_/A sky130_fd_sc_hd__clkinv_8
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__333__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ _288_/B _250_/B _259_/X VGND VGND VPWR VPWR _261_/A sky130_fd_sc_hd__o21ai_2
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_191_ _385_/Q _187_/Y _370_/Q _233_/B VGND VGND VPWR VPWR _385_/D sky130_fd_sc_hd__a22o_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__328__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_174_ _368_/Q VGND VGND VPWR VPWR _274_/A sky130_fd_sc_hd__inv_2
X_243_ _273_/B VGND VGND VPWR VPWR _243_/Y sky130_fd_sc_hd__inv_2
X_312_ _296_/A _246_/B _310_/B _378_/Q _239_/B VGND VGND VPWR VPWR _312_/X sky130_fd_sc_hd__o311a_2
XFILLER_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[11\].id.delayenb0 ringosc.dstage\[11\].id.delayenb1/A _338_/X VGND
+ VGND VPWR VPWR ringosc.iss.delayenb1/A sky130_fd_sc_hd__einvn_8
XFILLER_8_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_226_ _226_/A _226_/B VGND VGND VPWR VPWR _250_/B sky130_fd_sc_hd__or2_2
X_209_ div[3] _209_/B VGND VGND VPWR VPWR _210_/A sky130_fd_sc_hd__or2_2
XFILLER_5_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_190_ dco _190_/B VGND VGND VPWR VPWR _335_/A sky130_fd_sc_hd__nor2_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_173_ _384_/Q VGND VGND VPWR VPWR _206_/B sky130_fd_sc_hd__inv_2
X_311_ _305_/A _376_/Q _375_/Q _310_/X VGND VGND VPWR VPWR _311_/X sky130_fd_sc_hd__o31a_2
X_242_ _309_/A _255_/B _231_/X _241_/X VGND VGND VPWR VPWR _273_/B sky130_fd_sc_hd__o31a_2
X_225_ _168_/Y _219_/B div[4] _223_/B _221_/X VGND VGND VPWR VPWR _226_/B sky130_fd_sc_hd__o221ai_2
Xringosc.dstage\[11\].id.delayenb1 ringosc.dstage\[11\].id.delayenb1/A _339_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[11\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_208_ div[3] _209_/B div[2] _207_/X VGND VGND VPWR VPWR _208_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__211__A1 div[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_310_ _378_/Q _310_/B _310_/C VGND VGND VPWR VPWR _310_/X sky130_fd_sc_hd__and3_2
X_172_ _369_/Q VGND VGND VPWR VPWR _274_/C sky130_fd_sc_hd__inv_2
Xringosc.dstage\[2\].id.delayen0 ringosc.dstage\[2\].id.delayen0/A _356_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
Xringosc.iss.const1 VGND VGND VPWR VPWR ringosc.iss.const1/HI ringosc.iss.const1/LO
+ sky130_fd_sc_hd__conb_1
X_241_ _226_/B _232_/Y _250_/B _240_/X _233_/X VGND VGND VPWR VPWR _241_/X sky130_fd_sc_hd__o221a_2
X_224_ _208_/Y _210_/Y _212_/Y _218_/Y _223_/Y VGND VGND VPWR VPWR _226_/A sky130_fd_sc_hd__o221a_2
XFILLER_8_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_207_ _207_/A _207_/B VGND VGND VPWR VPWR _207_/X sky130_fd_sc_hd__xor2_1
Xringosc.dstage\[6\].id.delayenb0 ringosc.dstage\[6\].id.delayenb1/A _348_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[6\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[11\].id.delaybuf0 ringosc.dstage\[10\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_386_ _336_/A _386_/D _335_/X VGND VGND VPWR VPWR _386_/Q sky130_fd_sc_hd__dfrtp_2
X_171_ _385_/Q VGND VGND VPWR VPWR _199_/B sky130_fd_sc_hd__inv_2
Xringosc.dstage\[2\].id.delayen1 ringosc.dstage\[2\].id.delayen1/A _357_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_240_ _373_/Q _372_/Q _240_/C VGND VGND VPWR VPWR _240_/X sky130_fd_sc_hd__or3_2
X_369_ _336_/A _369_/D _328_/X VGND VGND VPWR VPWR _369_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__350__A1 ext_trim[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_223_ div[4] _223_/B VGND VGND VPWR VPWR _223_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__341__A1 ext_trim[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_206_ _274_/C _206_/B VGND VGND VPWR VPWR _207_/B sky130_fd_sc_hd__xor2_1
Xringosc.dstage\[6\].id.delayenb1 ringosc.dstage\[6\].id.delayenb1/A _349_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[6\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[11\].id.delaybuf1 ringosc.dstage\[11\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_385_ _336_/A _385_/D _335_/A VGND VGND VPWR VPWR _385_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.iss.delayen0 ringosc.iss.delayen0/A _362_/X VGND VGND VPWR VPWR ringosc.ibufp00/A
+ sky130_fd_sc_hd__einvp_2
X_170_ _370_/Q VGND VGND VPWR VPWR _274_/D sky130_fd_sc_hd__inv_2
X_368_ _336_/A _368_/D _329_/X VGND VGND VPWR VPWR _368_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__189__A enable VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_299_ _377_/Q _376_/Q _375_/Q _378_/Q VGND VGND VPWR VPWR _299_/X sky130_fd_sc_hd__a31o_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_222_ _221_/A _221_/B _221_/X VGND VGND VPWR VPWR _223_/B sky130_fd_sc_hd__a21bo_2
XFILLER_6_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_205_ _199_/X _204_/X _199_/X _204_/X VGND VGND VPWR VPWR _209_/B sky130_fd_sc_hd__a2bb2o_2
Xringosc.dstage\[6\].id.delaybuf0 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.dstage\[6\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[2\].id.delayenb0 ringosc.dstage\[2\].id.delayenb1/A _356_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[2\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[10\].id.delayint0 ringosc.dstage\[10\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[9\].id.delayint0 ringosc.dstage\[9\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_384_ _336_/A _384_/D _313_/X VGND VGND VPWR VPWR _384_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.iss.delayen1 ringosc.iss.delayen1/A _363_/X VGND VGND VPWR VPWR ringosc.iss.delayen1/Z
+ sky130_fd_sc_hd__einvp_2
XFILLER_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_298_ _377_/Q _376_/Q _305_/C _378_/Q VGND VGND VPWR VPWR _298_/X sky130_fd_sc_hd__a31o_2
X_367_ _336_/A _367_/D _330_/X VGND VGND VPWR VPWR _367_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__189__B resetb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_221_ _221_/A _221_/B VGND VGND VPWR VPWR _221_/X sky130_fd_sc_hd__or2_2
X_204_ _274_/C _206_/B _200_/Y _207_/A VGND VGND VPWR VPWR _204_/X sky130_fd_sc_hd__o22a_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[6\].id.delaybuf1 ringosc.dstage\[6\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[2\].id.delayenb1 ringosc.dstage\[2\].id.delayenb1/A _357_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[2\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_383_ _336_/A _383_/D _314_/X VGND VGND VPWR VPWR _383_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__362__A1 ext_trim[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__353__A1 ext_trim[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__340__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_366_ _336_/A _366_/D _331_/X VGND VGND VPWR VPWR _366_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__344__A1 ext_trim[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_297_ _305_/A _376_/Q _378_/Q _292_/X VGND VGND VPWR VPWR _297_/X sky130_fd_sc_hd__o31a_2
X_220_ _274_/D _199_/B _198_/Y _204_/X VGND VGND VPWR VPWR _221_/B sky130_fd_sc_hd__o22a_2
X_349_ _307_/B ext_trim[19] dco VGND VGND VPWR VPWR _349_/X sky130_fd_sc_hd__mux2_1
X_203_ _274_/A _202_/B _201_/X _202_/X VGND VGND VPWR VPWR _207_/A sky130_fd_sc_hd__o22a_2
Xringosc.iss.ctrlen0 _190_/B _362_/X VGND VGND VPWR VPWR ringosc.iss.ctrlen0/X sky130_fd_sc_hd__or2_2
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__217__B1 div[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__208__B1 div[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__343__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[2\].id.delaybuf0 ringosc.dstage\[1\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[5\].id.delayint0 ringosc.dstage\[5\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_382_ _336_/A _382_/D _315_/X VGND VGND VPWR VPWR _382_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__338__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_365_ _336_/A _365_/D _332_/X VGND VGND VPWR VPWR _366_/D sky130_fd_sc_hd__dfrtp_2
X_296_ _296_/A _296_/B VGND VGND VPWR VPWR _296_/X sky130_fd_sc_hd__or2_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__351__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_348_ _287_/X ext_trim[6] dco VGND VGND VPWR VPWR _348_/X sky130_fd_sc_hd__mux2_1
X_279_ _274_/A _282_/B _274_/C VGND VGND VPWR VPWR _279_/Y sky130_fd_sc_hd__o21ai_2
X_202_ _368_/Q _202_/B VGND VGND VPWR VPWR _202_/X sky130_fd_sc_hd__xor2_1
XANTENNA__346__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__217__A1 div[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[7\].id.delayen0 ringosc.dstage\[7\].id.delayen0/A _346_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[7\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XANTENNA__208__A1 div[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[2\].id.delaybuf1 ringosc.dstage\[2\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__354__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_381_ _336_/A _381_/D _316_/X VGND VGND VPWR VPWR _381_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__349__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_364_ _336_/A osc _333_/X VGND VGND VPWR VPWR _365_/D sky130_fd_sc_hd__dfrtp_2
X_295_ _305_/A _376_/Q _378_/Q _296_/A _292_/X VGND VGND VPWR VPWR _295_/X sky130_fd_sc_hd__o41a_2
X_278_ _371_/Q _275_/A _187_/Y _277_/X VGND VGND VPWR VPWR _370_/D sky130_fd_sc_hd__o211a_2
X_347_ _311_/X ext_trim[20] dco VGND VGND VPWR VPWR _347_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_201_ _282_/B _215_/B VGND VGND VPWR VPWR _201_/X sky130_fd_sc_hd__or2_2
XANTENNA__362__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[11\].id.delayen0 ringosc.dstage\[11\].id.delayen0/A _338_/X VGND
+ VGND VPWR VPWR ringosc.iss.delayenb1/A sky130_fd_sc_hd__einvp_2
Xringosc.dstage\[7\].id.delayen1 ringosc.dstage\[7\].id.delayen1/A _347_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[7\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XANTENNA__357__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__356__A1 ext_trim[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_380_ _336_/A _380_/D _317_/X VGND VGND VPWR VPWR _380_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__347__A1 ext_trim[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

