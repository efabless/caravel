magic
tech sky130A
magscale 1 2
timestamp 1638477072
<< locali >>
rect 8125 9911 8159 10149
rect 13093 5627 13127 5797
rect 15669 3519 15703 3621
rect 3985 2839 4019 3009
<< viali >>
rect 7297 10761 7331 10795
rect 10425 10761 10459 10795
rect 12909 10761 12943 10795
rect 14013 10761 14047 10795
rect 18337 10761 18371 10795
rect 10333 10693 10367 10727
rect 11529 10693 11563 10727
rect 13553 10693 13587 10727
rect 13645 10693 13679 10727
rect 15209 10693 15243 10727
rect 1593 10625 1627 10659
rect 2329 10625 2363 10659
rect 2605 10625 2639 10659
rect 2697 10625 2731 10659
rect 2789 10625 2823 10659
rect 7481 10625 7515 10659
rect 10149 10625 10183 10659
rect 10609 10625 10643 10659
rect 11345 10625 11379 10659
rect 12081 10625 12115 10659
rect 13093 10625 13127 10659
rect 15117 10625 15151 10659
rect 15393 10625 15427 10659
rect 18061 10625 18095 10659
rect 18245 10625 18279 10659
rect 18521 10625 18555 10659
rect 1685 10557 1719 10591
rect 2053 10557 2087 10591
rect 2973 10557 3007 10591
rect 11621 10557 11655 10591
rect 13369 10557 13403 10591
rect 17877 10557 17911 10591
rect 14473 10489 14507 10523
rect 18061 10489 18095 10523
rect 1409 10421 1443 10455
rect 2237 10421 2271 10455
rect 11069 10421 11103 10455
rect 12725 10421 12759 10455
rect 14197 10421 14231 10455
rect 15025 10421 15059 10455
rect 15945 10421 15979 10455
rect 1409 10217 1443 10251
rect 5825 10217 5859 10251
rect 13093 10217 13127 10251
rect 17831 10217 17865 10251
rect 8125 10149 8159 10183
rect 8309 10149 8343 10183
rect 2697 10081 2731 10115
rect 6101 10081 6135 10115
rect 1501 10013 1535 10047
rect 2973 10013 3007 10047
rect 3157 10013 3191 10047
rect 3525 10013 3559 10047
rect 3709 10013 3743 10047
rect 3985 9945 4019 9979
rect 6377 9945 6411 9979
rect 8493 10081 8527 10115
rect 11345 10081 11379 10115
rect 16405 10081 16439 10115
rect 8861 10013 8895 10047
rect 11069 10013 11103 10047
rect 13277 10013 13311 10047
rect 13369 10013 13403 10047
rect 13553 10013 13587 10047
rect 13921 10013 13955 10047
rect 15761 10013 15795 10047
rect 15853 10013 15887 10047
rect 16037 10013 16071 10047
rect 18245 10013 18279 10047
rect 18521 10013 18555 10047
rect 10609 9945 10643 9979
rect 11161 9945 11195 9979
rect 11621 9945 11655 9979
rect 3249 9877 3283 9911
rect 3433 9877 3467 9911
rect 5457 9877 5491 9911
rect 7849 9877 7883 9911
rect 8125 9877 8159 9911
rect 10287 9877 10321 9911
rect 10885 9877 10919 9911
rect 15347 9877 15381 9911
rect 18337 9877 18371 9911
rect 2053 9673 2087 9707
rect 2697 9673 2731 9707
rect 3985 9673 4019 9707
rect 8585 9673 8619 9707
rect 11805 9673 11839 9707
rect 581 9605 615 9639
rect 2237 9605 2271 9639
rect 4997 9605 5031 9639
rect 16635 9605 16669 9639
rect 2145 9537 2179 9571
rect 2329 9537 2363 9571
rect 2513 9537 2547 9571
rect 2789 9537 2823 9571
rect 2973 9537 3007 9571
rect 3709 9537 3743 9571
rect 3893 9537 3927 9571
rect 4353 9537 4387 9571
rect 5089 9537 5123 9571
rect 7665 9537 7699 9571
rect 8677 9537 8711 9571
rect 9321 9537 9355 9571
rect 9505 9537 9539 9571
rect 10057 9537 10091 9571
rect 10425 9537 10459 9571
rect 10692 9537 10726 9571
rect 12541 9537 12575 9571
rect 14289 9537 14323 9571
rect 305 9469 339 9503
rect 4445 9469 4479 9503
rect 4537 9469 4571 9503
rect 5365 9469 5399 9503
rect 5641 9469 5675 9503
rect 7757 9469 7791 9503
rect 7941 9469 7975 9503
rect 8861 9469 8895 9503
rect 9413 9469 9447 9503
rect 9965 9469 9999 9503
rect 14841 9469 14875 9503
rect 15209 9469 15243 9503
rect 7113 9401 7147 9435
rect 8217 9401 8251 9435
rect 9689 9401 9723 9435
rect 3157 9333 3191 9367
rect 3525 9333 3559 9367
rect 3801 9333 3835 9367
rect 5273 9333 5307 9367
rect 7297 9333 7331 9367
rect 12449 9333 12483 9367
rect 14657 9333 14691 9367
rect 2789 9129 2823 9163
rect 6285 9129 6319 9163
rect 9045 9129 9079 9163
rect 12357 9129 12391 9163
rect 2145 9061 2179 9095
rect 2237 9061 2271 9095
rect 2513 9061 2547 9095
rect 2329 8993 2363 9027
rect 3157 8993 3191 9027
rect 4813 8993 4847 9027
rect 6469 8993 6503 9027
rect 6561 8993 6595 9027
rect 10241 8993 10275 9027
rect 11713 8993 11747 9027
rect 13001 8993 13035 9027
rect 15025 8993 15059 9027
rect 581 8925 615 8959
rect 1777 8925 1811 8959
rect 2605 8925 2639 8959
rect 2697 8925 2731 8959
rect 3065 8925 3099 8959
rect 3341 8925 3375 8959
rect 3525 8925 3559 8959
rect 4537 8925 4571 8959
rect 4721 8925 4755 8959
rect 4905 8925 4939 8959
rect 5089 8925 5123 8959
rect 7021 8925 7055 8959
rect 8769 8925 8803 8959
rect 9229 8925 9263 8959
rect 9321 8925 9355 8959
rect 9781 8925 9815 8959
rect 10057 8925 10091 8959
rect 10333 8925 10367 8959
rect 11621 8925 11655 8959
rect 12725 8925 12759 8959
rect 15853 8925 15887 8959
rect 5733 8857 5767 8891
rect 5917 8857 5951 8891
rect 7113 8857 7147 8891
rect 7297 8857 7331 8891
rect 9873 8857 9907 8891
rect 11529 8857 11563 8891
rect 14749 8857 14783 8891
rect 16129 8857 16163 8891
rect 17877 8857 17911 8891
rect 489 8789 523 8823
rect 2329 8789 2363 8823
rect 3433 8789 3467 8823
rect 4629 8789 4663 8823
rect 6929 8789 6963 8823
rect 7021 8789 7055 8823
rect 8861 8789 8895 8823
rect 9689 8789 9723 8823
rect 9781 8789 9815 8823
rect 10701 8789 10735 8823
rect 11161 8789 11195 8823
rect 12265 8789 12299 8823
rect 12817 8789 12851 8823
rect 13277 8789 13311 8823
rect 15209 8789 15243 8823
rect 15669 8789 15703 8823
rect 2099 8585 2133 8619
rect 4905 8585 4939 8619
rect 6469 8585 6503 8619
rect 7113 8585 7147 8619
rect 7297 8585 7331 8619
rect 10701 8585 10735 8619
rect 11069 8585 11103 8619
rect 12449 8585 12483 8619
rect 14289 8585 14323 8619
rect 5549 8517 5583 8551
rect 7389 8517 7423 8551
rect 7573 8517 7607 8551
rect 9781 8517 9815 8551
rect 10149 8517 10183 8551
rect 10425 8517 10459 8551
rect 11161 8517 11195 8551
rect 12817 8517 12851 8551
rect 305 8449 339 8483
rect 673 8449 707 8483
rect 2881 8449 2915 8483
rect 3065 8449 3099 8483
rect 3893 8449 3927 8483
rect 4169 8449 4203 8483
rect 4261 8449 4295 8483
rect 5181 8449 5215 8483
rect 5365 8449 5399 8483
rect 6653 8449 6687 8483
rect 7297 8449 7331 8483
rect 8217 8449 8251 8483
rect 8677 8449 8711 8483
rect 8769 8449 8803 8483
rect 9689 8449 9723 8483
rect 9965 8449 9999 8483
rect 10241 8449 10275 8483
rect 10333 8449 10367 8483
rect 12541 8449 12575 8483
rect 14473 8449 14507 8483
rect 14657 8449 14691 8483
rect 18245 8449 18279 8483
rect 18521 8449 18555 8483
rect 3985 8381 4019 8415
rect 4905 8381 4939 8415
rect 5089 8381 5123 8415
rect 6745 8381 6779 8415
rect 8309 8381 8343 8415
rect 8493 8381 8527 8415
rect 11253 8381 11287 8415
rect 14841 8381 14875 8415
rect 15209 8381 15243 8415
rect 4077 8313 4111 8347
rect 9873 8313 9907 8347
rect 14657 8313 14691 8347
rect 18337 8313 18371 8347
rect 2329 8245 2363 8279
rect 2973 8245 3007 8279
rect 7849 8245 7883 8279
rect 16635 8245 16669 8279
rect 15117 8041 15151 8075
rect 1961 7973 1995 8007
rect 2743 7973 2777 8007
rect 7297 7973 7331 8007
rect 10057 7973 10091 8007
rect 13645 7973 13679 8007
rect 1777 7905 1811 7939
rect 2329 7905 2363 7939
rect 2513 7905 2547 7939
rect 4353 7905 4387 7939
rect 7941 7905 7975 7939
rect 13277 7905 13311 7939
rect 14013 7905 14047 7939
rect 14473 7905 14507 7939
rect 15761 7905 15795 7939
rect 16129 7905 16163 7939
rect 17509 7905 17543 7939
rect 2053 7837 2087 7871
rect 2237 7837 2271 7871
rect 2421 7837 2455 7871
rect 4537 7837 4571 7871
rect 4721 7837 4755 7871
rect 4997 7837 5031 7871
rect 5089 7837 5123 7871
rect 5457 7837 5491 7871
rect 5549 7837 5583 7871
rect 5733 7837 5767 7871
rect 6285 7837 6319 7871
rect 7665 7837 7699 7871
rect 9413 7837 9447 7871
rect 9505 7837 9539 7871
rect 9597 7837 9631 7871
rect 9873 7837 9907 7871
rect 10057 7837 10091 7871
rect 10333 7837 10367 7871
rect 10425 7837 10459 7871
rect 10517 7837 10551 7871
rect 10701 7837 10735 7871
rect 13461 7837 13495 7871
rect 14105 7837 14139 7871
rect 14749 7837 14783 7871
rect 4077 7769 4111 7803
rect 5181 7769 5215 7803
rect 5365 7769 5399 7803
rect 6837 7769 6871 7803
rect 7021 7769 7055 7803
rect 9781 7769 9815 7803
rect 11345 7769 11379 7803
rect 1777 7701 1811 7735
rect 3709 7701 3743 7735
rect 4169 7701 4203 7735
rect 4813 7701 4847 7735
rect 5273 7701 5307 7735
rect 5641 7701 5675 7735
rect 6193 7701 6227 7735
rect 7757 7701 7791 7735
rect 10425 7701 10459 7735
rect 11437 7701 11471 7735
rect 14657 7701 14691 7735
rect 15485 7701 15519 7735
rect 2237 7497 2271 7531
rect 2697 7497 2731 7531
rect 3065 7497 3099 7531
rect 3157 7497 3191 7531
rect 9781 7497 9815 7531
rect 9965 7497 9999 7531
rect 12633 7497 12667 7531
rect 13461 7497 13495 7531
rect 581 7429 615 7463
rect 13553 7429 13587 7463
rect 14197 7429 14231 7463
rect 2329 7361 2363 7395
rect 5181 7361 5215 7395
rect 5549 7361 5583 7395
rect 6975 7361 7009 7395
rect 7481 7361 7515 7395
rect 8769 7361 8803 7395
rect 10425 7361 10459 7395
rect 11851 7361 11885 7395
rect 12265 7361 12299 7395
rect 12909 7361 12943 7395
rect 13185 7361 13219 7395
rect 13369 7361 13403 7395
rect 13461 7361 13495 7395
rect 13734 7361 13768 7395
rect 14013 7361 14047 7395
rect 14289 7361 14323 7395
rect 17049 7361 17083 7395
rect 305 7293 339 7327
rect 2053 7293 2087 7327
rect 3341 7293 3375 7327
rect 7389 7293 7423 7327
rect 8493 7293 8527 7327
rect 10057 7293 10091 7327
rect 12173 7293 12207 7327
rect 14473 7293 14507 7327
rect 14841 7293 14875 7327
rect 8953 7225 8987 7259
rect 13277 7225 13311 7259
rect 13829 7225 13863 7259
rect 2605 7157 2639 7191
rect 5089 7157 5123 7191
rect 8585 7157 8619 7191
rect 13001 7157 13035 7191
rect 16267 7157 16301 7191
rect 16865 7157 16899 7191
rect 2145 6953 2179 6987
rect 11621 6953 11655 6987
rect 14381 6953 14415 6987
rect 16116 6953 16150 6987
rect 2605 6885 2639 6919
rect 7941 6885 7975 6919
rect 15301 6885 15335 6919
rect 1961 6817 1995 6851
rect 3065 6817 3099 6851
rect 4353 6817 4387 6851
rect 9137 6817 9171 6851
rect 11345 6817 11379 6851
rect 14105 6817 14139 6851
rect 14841 6817 14875 6851
rect 14933 6817 14967 6851
rect 2237 6749 2271 6783
rect 2605 6749 2639 6783
rect 2789 6749 2823 6783
rect 2881 6749 2915 6783
rect 2973 6749 3007 6783
rect 3157 6749 3191 6783
rect 6561 6749 6595 6783
rect 8125 6749 8159 6783
rect 8309 6749 8343 6783
rect 11069 6749 11103 6783
rect 11253 6749 11287 6783
rect 11721 6749 11755 6783
rect 14013 6749 14047 6783
rect 14197 6749 14231 6783
rect 15393 6749 15427 6783
rect 15853 6749 15887 6783
rect 18245 6749 18279 6783
rect 18521 6749 18555 6783
rect 2329 6681 2363 6715
rect 2513 6681 2547 6715
rect 6806 6681 6840 6715
rect 10701 6681 10735 6715
rect 11805 6681 11839 6715
rect 15761 6681 15795 6715
rect 17877 6681 17911 6715
rect 1961 6613 1995 6647
rect 3709 6613 3743 6647
rect 4077 6613 4111 6647
rect 4169 6613 4203 6647
rect 8217 6613 8251 6647
rect 10885 6613 10919 6647
rect 13645 6613 13679 6647
rect 13829 6613 13863 6647
rect 14749 6613 14783 6647
rect 18337 6613 18371 6647
rect 3893 6409 3927 6443
rect 4905 6409 4939 6443
rect 5365 6409 5399 6443
rect 8401 6409 8435 6443
rect 16681 6409 16715 6443
rect 16865 6409 16899 6443
rect 17233 6409 17267 6443
rect 17693 6409 17727 6443
rect 18061 6409 18095 6443
rect 9965 6341 9999 6375
rect 15209 6341 15243 6375
rect 305 6273 339 6307
rect 2145 6273 2179 6307
rect 2329 6273 2363 6307
rect 2789 6273 2823 6307
rect 4261 6273 4295 6307
rect 4353 6273 4387 6307
rect 5273 6273 5307 6307
rect 8125 6273 8159 6307
rect 8493 6273 8527 6307
rect 9045 6273 9079 6307
rect 9229 6273 9263 6307
rect 9321 6273 9355 6307
rect 9689 6273 9723 6307
rect 12081 6273 12115 6307
rect 14657 6273 14691 6307
rect 14933 6273 14967 6307
rect 17325 6273 17359 6307
rect 581 6205 615 6239
rect 2237 6205 2271 6239
rect 2513 6205 2547 6239
rect 2697 6205 2731 6239
rect 4445 6205 4479 6239
rect 5457 6205 5491 6239
rect 8401 6205 8435 6239
rect 11713 6205 11747 6239
rect 12357 6205 12391 6239
rect 17417 6205 17451 6239
rect 18153 6205 18187 6239
rect 18245 6205 18279 6239
rect 2605 6137 2639 6171
rect 8217 6137 8251 6171
rect 2053 6069 2087 6103
rect 2881 6069 2915 6103
rect 8769 6069 8803 6103
rect 8953 6069 8987 6103
rect 11897 6069 11931 6103
rect 13829 6069 13863 6103
rect 14565 6069 14599 6103
rect 14749 6069 14783 6103
rect 2421 5865 2455 5899
rect 3249 5865 3283 5899
rect 5641 5865 5675 5899
rect 7481 5865 7515 5899
rect 7849 5865 7883 5899
rect 10609 5865 10643 5899
rect 17831 5865 17865 5899
rect 11161 5797 11195 5831
rect 11989 5797 12023 5831
rect 12265 5797 12299 5831
rect 13093 5797 13127 5831
rect 14657 5797 14691 5831
rect 2973 5729 3007 5763
rect 3433 5729 3467 5763
rect 4997 5729 5031 5763
rect 12817 5729 12851 5763
rect 765 5661 799 5695
rect 2329 5661 2363 5695
rect 2881 5661 2915 5695
rect 3341 5661 3375 5695
rect 3525 5661 3559 5695
rect 3709 5661 3743 5695
rect 3985 5661 4019 5695
rect 4537 5661 4571 5695
rect 6101 5661 6135 5695
rect 7573 5661 7607 5695
rect 10425 5661 10459 5695
rect 11805 5661 11839 5695
rect 12725 5661 12759 5695
rect 13737 5729 13771 5763
rect 14289 5729 14323 5763
rect 15301 5729 15335 5763
rect 16405 5729 16439 5763
rect 13553 5661 13587 5695
rect 13823 5661 13857 5695
rect 14170 5661 14204 5695
rect 16037 5661 16071 5695
rect 18245 5661 18279 5695
rect 18521 5661 18555 5695
rect 5181 5593 5215 5627
rect 6368 5593 6402 5627
rect 8677 5593 8711 5627
rect 10977 5593 11011 5627
rect 12633 5593 12667 5627
rect 13093 5593 13127 5627
rect 15117 5593 15151 5627
rect 673 5525 707 5559
rect 3985 5525 4019 5559
rect 5273 5525 5307 5559
rect 8033 5525 8067 5559
rect 13829 5525 13863 5559
rect 14565 5525 14599 5559
rect 15025 5525 15059 5559
rect 15853 5525 15887 5559
rect 18337 5525 18371 5559
rect 2283 5321 2317 5355
rect 4445 5321 4479 5355
rect 8861 5321 8895 5355
rect 9137 5253 9171 5287
rect 9321 5253 9355 5287
rect 17233 5253 17267 5287
rect 489 5185 523 5219
rect 857 5185 891 5219
rect 4077 5185 4111 5219
rect 7481 5185 7515 5219
rect 7748 5185 7782 5219
rect 9045 5185 9079 5219
rect 13461 5185 13495 5219
rect 14933 5185 14967 5219
rect 16957 5185 16991 5219
rect 3985 5117 4019 5151
rect 9873 5117 9907 5151
rect 10149 5117 10183 5151
rect 13553 5117 13587 5151
rect 15209 5117 15243 5151
rect 9045 5049 9079 5083
rect 2605 4981 2639 5015
rect 9689 4981 9723 5015
rect 11621 4981 11655 5015
rect 13829 4981 13863 5015
rect 14749 4981 14783 5015
rect 16681 4981 16715 5015
rect 11161 4777 11195 4811
rect 13737 4777 13771 4811
rect 11805 4709 11839 4743
rect 3709 4641 3743 4675
rect 6101 4641 6135 4675
rect 8493 4641 8527 4675
rect 11621 4641 11655 4675
rect 15209 4641 15243 4675
rect 15485 4641 15519 4675
rect 17601 4641 17635 4675
rect 765 4573 799 4607
rect 6469 4573 6503 4607
rect 7941 4573 7975 4607
rect 8033 4573 8067 4607
rect 11529 4573 11563 4607
rect 11805 4573 11839 4607
rect 11897 4573 11931 4607
rect 12173 4573 12207 4607
rect 12357 4573 12391 4607
rect 17877 4573 17911 4607
rect 3985 4505 4019 4539
rect 8769 4505 8803 4539
rect 12081 4505 12115 4539
rect 15853 4505 15887 4539
rect 673 4437 707 4471
rect 2513 4437 2547 4471
rect 3433 4437 3467 4471
rect 5457 4437 5491 4471
rect 5917 4437 5951 4471
rect 8217 4437 8251 4471
rect 10241 4437 10275 4471
rect 12265 4437 12299 4471
rect 13553 4437 13587 4471
rect 15669 4437 15703 4471
rect 2513 4233 2547 4267
rect 3525 4233 3559 4267
rect 3985 4233 4019 4267
rect 6285 4233 6319 4267
rect 7665 4233 7699 4267
rect 8125 4233 8159 4267
rect 8493 4233 8527 4267
rect 8953 4233 8987 4267
rect 10057 4233 10091 4267
rect 10517 4233 10551 4267
rect 3341 4165 3375 4199
rect 7021 4165 7055 4199
rect 14565 4165 14599 4199
rect 489 4097 523 4131
rect 2789 4097 2823 4131
rect 3065 4097 3099 4131
rect 3249 4097 3283 4131
rect 3801 4097 3835 4131
rect 3893 4097 3927 4131
rect 4169 4087 4203 4121
rect 4353 4097 4387 4131
rect 4997 4097 5031 4131
rect 5181 4097 5215 4131
rect 6469 4097 6503 4131
rect 7757 4097 7791 4131
rect 8585 4097 8619 4131
rect 9137 4097 9171 4131
rect 10885 4097 10919 4131
rect 11493 4097 11527 4131
rect 11621 4097 11655 4131
rect 11713 4097 11747 4131
rect 12081 4097 12115 4131
rect 12265 4097 12299 4131
rect 18245 4097 18279 4131
rect 18521 4097 18555 4131
rect 857 4029 891 4063
rect 2513 4029 2547 4063
rect 2973 4029 3007 4063
rect 7849 4029 7883 4063
rect 8769 4029 8803 4063
rect 10149 4029 10183 4063
rect 10241 4029 10275 4063
rect 10977 4029 11011 4063
rect 11069 4029 11103 4063
rect 12449 4029 12483 4063
rect 12817 4029 12851 4063
rect 14749 4029 14783 4063
rect 16497 4029 16531 4063
rect 2283 3961 2317 3995
rect 6837 3961 6871 3995
rect 7297 3961 7331 3995
rect 9689 3961 9723 3995
rect 12173 3961 12207 3995
rect 2697 3893 2731 3927
rect 3709 3893 3743 3927
rect 4261 3893 4295 3927
rect 4997 3893 5031 3927
rect 11897 3893 11931 3927
rect 14243 3893 14277 3927
rect 16239 3893 16273 3927
rect 18337 3893 18371 3927
rect 2789 3689 2823 3723
rect 10057 3689 10091 3723
rect 12909 3689 12943 3723
rect 18153 3689 18187 3723
rect 2697 3621 2731 3655
rect 4353 3621 4387 3655
rect 14289 3621 14323 3655
rect 14565 3621 14599 3655
rect 15669 3621 15703 3655
rect 2237 3553 2271 3587
rect 3709 3553 3743 3587
rect 6193 3553 6227 3587
rect 6285 3553 6319 3587
rect 6469 3553 6503 3587
rect 9689 3553 9723 3587
rect 12541 3553 12575 3587
rect 13921 3553 13955 3587
rect 15117 3553 15151 3587
rect 1777 3485 1811 3519
rect 1869 3485 1903 3519
rect 2881 3485 2915 3519
rect 3157 3485 3191 3519
rect 3341 3485 3375 3519
rect 3893 3485 3927 3519
rect 3985 3485 4019 3519
rect 4077 3485 4111 3519
rect 4537 3485 4571 3519
rect 5733 3485 5767 3519
rect 5917 3485 5951 3519
rect 6561 3485 6595 3519
rect 7849 3485 7883 3519
rect 8125 3485 8159 3519
rect 8309 3485 8343 3519
rect 9781 3485 9815 3519
rect 12633 3485 12667 3519
rect 15025 3485 15059 3519
rect 15669 3485 15703 3519
rect 15761 3485 15795 3519
rect 16129 3485 16163 3519
rect 2329 3417 2363 3451
rect 7757 3417 7791 3451
rect 14933 3417 14967 3451
rect 17877 3417 17911 3451
rect 18245 3417 18279 3451
rect 1593 3349 1627 3383
rect 3065 3349 3099 3383
rect 5825 3349 5859 3383
rect 6193 3349 6227 3383
rect 8585 3349 8619 3383
rect 12265 3349 12299 3383
rect 14381 3349 14415 3383
rect 15485 3349 15519 3383
rect 2053 3145 2087 3179
rect 2605 3145 2639 3179
rect 3157 3145 3191 3179
rect 5457 3145 5491 3179
rect 5917 3145 5951 3179
rect 14657 3145 14691 3179
rect 14887 3145 14921 3179
rect 581 3077 615 3111
rect 4537 3077 4571 3111
rect 7389 3077 7423 3111
rect 7573 3077 7607 3111
rect 7941 3077 7975 3111
rect 2697 3009 2731 3043
rect 3065 3009 3099 3043
rect 3249 3009 3283 3043
rect 3709 3009 3743 3043
rect 3893 3009 3927 3043
rect 3985 3009 4019 3043
rect 4169 3009 4203 3043
rect 4261 3009 4295 3043
rect 4445 3009 4479 3043
rect 4629 3009 4663 3043
rect 5825 3009 5859 3043
rect 7665 3009 7699 3043
rect 7757 3009 7791 3043
rect 8217 3009 8251 3043
rect 9965 3009 9999 3043
rect 10057 3009 10091 3043
rect 11851 3009 11885 3043
rect 12449 3009 12483 3043
rect 13553 3009 13587 3043
rect 13737 3009 13771 3043
rect 14289 3009 14323 3043
rect 14565 3009 14599 3043
rect 14749 3009 14783 3043
rect 16313 3009 16347 3043
rect 305 2941 339 2975
rect 6009 2941 6043 2975
rect 6285 2941 6319 2975
rect 9873 2941 9907 2975
rect 10425 2941 10459 2975
rect 12357 2941 12391 2975
rect 14105 2941 14139 2975
rect 16681 2941 16715 2975
rect 8401 2873 8435 2907
rect 12817 2873 12851 2907
rect 2237 2805 2271 2839
rect 3801 2805 3835 2839
rect 3985 2805 4019 2839
rect 6745 2805 6779 2839
rect 7849 2805 7883 2839
rect 9413 2805 9447 2839
rect 3249 2601 3283 2635
rect 6745 2601 6779 2635
rect 7573 2601 7607 2635
rect 10287 2601 10321 2635
rect 6469 2533 6503 2567
rect 13001 2533 13035 2567
rect 3065 2465 3099 2499
rect 3709 2465 3743 2499
rect 3985 2465 4019 2499
rect 4813 2465 4847 2499
rect 8861 2465 8895 2499
rect 11529 2465 11563 2499
rect 13277 2465 13311 2499
rect 13829 2465 13863 2499
rect 15853 2465 15887 2499
rect 17877 2465 17911 2499
rect 3341 2397 3375 2431
rect 6285 2397 6319 2431
rect 6469 2397 6503 2431
rect 6929 2397 6963 2431
rect 7113 2397 7147 2431
rect 7573 2397 7607 2431
rect 8125 2397 8159 2431
rect 8217 2397 8251 2431
rect 8493 2397 8527 2431
rect 12357 2397 12391 2431
rect 12449 2397 12483 2431
rect 12541 2397 12575 2431
rect 12725 2397 12759 2431
rect 12817 2397 12851 2431
rect 13553 2397 13587 2431
rect 13691 2397 13725 2431
rect 18245 2397 18279 2431
rect 18521 2397 18555 2431
rect 4905 2329 4939 2363
rect 6837 2329 6871 2363
rect 7297 2329 7331 2363
rect 7481 2329 7515 2363
rect 11345 2329 11379 2363
rect 12909 2329 12943 2363
rect 13093 2329 13127 2363
rect 14096 2329 14130 2363
rect 17601 2329 17635 2363
rect 3065 2261 3099 2295
rect 4997 2261 5031 2295
rect 5365 2261 5399 2295
rect 7941 2261 7975 2295
rect 10885 2261 10919 2295
rect 11253 2261 11287 2295
rect 13461 2261 13495 2295
rect 15209 2261 15243 2295
rect 15393 2261 15427 2295
rect 15669 2261 15703 2295
rect 18337 2261 18371 2295
rect 3801 2057 3835 2091
rect 4905 2057 4939 2091
rect 5273 2057 5307 2091
rect 5365 2057 5399 2091
rect 6377 2057 6411 2091
rect 9045 2057 9079 2091
rect 10609 2057 10643 2091
rect 11069 2057 11103 2091
rect 12633 2057 12667 2091
rect 857 1989 891 2023
rect 9229 1989 9263 2023
rect 14749 1989 14783 2023
rect 3065 1921 3099 1955
rect 3341 1921 3375 1955
rect 3433 1921 3467 1955
rect 3617 1921 3651 1955
rect 3893 1921 3927 1955
rect 6469 1921 6503 1955
rect 7297 1921 7331 1955
rect 9137 1921 9171 1955
rect 9413 1921 9447 1955
rect 9873 1921 9907 1955
rect 10701 1921 10735 1955
rect 11161 1921 11195 1955
rect 12541 1921 12575 1955
rect 13001 1921 13035 1955
rect 14289 1921 14323 1955
rect 14473 1921 14507 1955
rect 14657 1921 14691 1955
rect 14933 1921 14967 1955
rect 15301 1921 15335 1955
rect 15568 1921 15602 1955
rect 581 1853 615 1887
rect 2329 1853 2363 1887
rect 2789 1853 2823 1887
rect 3525 1853 3559 1887
rect 5549 1853 5583 1887
rect 6285 1853 6319 1887
rect 7573 1853 7607 1887
rect 9965 1853 9999 1887
rect 10241 1853 10275 1887
rect 10517 1853 10551 1887
rect 14013 1853 14047 1887
rect 14565 1853 14599 1887
rect 15209 1853 15243 1887
rect 3249 1785 3283 1819
rect 14105 1785 14139 1819
rect 15117 1785 15151 1819
rect 2513 1717 2547 1751
rect 2881 1717 2915 1751
rect 2973 1717 3007 1751
rect 6837 1717 6871 1751
rect 7113 1717 7147 1751
rect 9137 1717 9171 1751
rect 11253 1717 11287 1751
rect 12909 1717 12943 1751
rect 14197 1717 14231 1751
rect 16681 1717 16715 1751
rect 3801 1513 3835 1547
rect 5917 1513 5951 1547
rect 6101 1513 6135 1547
rect 10241 1513 10275 1547
rect 11161 1513 11195 1547
rect 14841 1513 14875 1547
rect 17601 1513 17635 1547
rect 1317 1377 1351 1411
rect 1593 1377 1627 1411
rect 3065 1377 3099 1411
rect 5641 1377 5675 1411
rect 6745 1377 6779 1411
rect 9137 1377 9171 1411
rect 9965 1377 9999 1411
rect 12909 1377 12943 1411
rect 13829 1377 13863 1411
rect 15209 1377 15243 1411
rect 16129 1377 16163 1411
rect 3433 1309 3467 1343
rect 3525 1309 3559 1343
rect 3893 1309 3927 1343
rect 5549 1309 5583 1343
rect 6469 1309 6503 1343
rect 8493 1309 8527 1343
rect 8677 1309 8711 1343
rect 8769 1309 8803 1343
rect 9873 1309 9907 1343
rect 10241 1309 10275 1343
rect 10425 1309 10459 1343
rect 11161 1309 11195 1343
rect 11253 1309 11287 1343
rect 12817 1309 12851 1343
rect 13737 1309 13771 1343
rect 15025 1309 15059 1343
rect 15853 1309 15887 1343
rect 17785 1309 17819 1343
rect 17877 1309 17911 1343
rect 18061 1309 18095 1343
rect 18153 1309 18187 1343
rect 3249 1241 3283 1275
rect 6561 1241 6595 1275
rect 10885 1241 10919 1275
rect 11069 1241 11103 1275
rect 11345 1241 11379 1275
rect 12725 1241 12759 1275
rect 14289 1241 14323 1275
rect 15669 1241 15703 1275
rect 18337 1241 18371 1275
rect 3525 1173 3559 1207
rect 4077 1173 4111 1207
rect 9413 1173 9447 1207
rect 9781 1173 9815 1207
rect 12357 1173 12391 1207
rect 13277 1173 13311 1207
rect 13645 1173 13679 1207
rect 18061 1173 18095 1207
rect 18521 1173 18555 1207
rect 2329 969 2363 1003
rect 5917 969 5951 1003
rect 7113 969 7147 1003
rect 10333 969 10367 1003
rect 11437 969 11471 1003
rect 14197 969 14231 1003
rect 18245 969 18279 1003
rect 5457 901 5491 935
rect 9183 901 9217 935
rect 9781 901 9815 935
rect 11805 901 11839 935
rect 14473 901 14507 935
rect 17110 901 17144 935
rect 2513 833 2547 867
rect 4307 833 4341 867
rect 4629 833 4663 867
rect 4997 833 5031 867
rect 5181 833 5215 867
rect 5733 833 5767 867
rect 5825 833 5859 867
rect 6009 833 6043 867
rect 6469 833 6503 867
rect 7389 833 7423 867
rect 9689 833 9723 867
rect 9965 833 9999 867
rect 10701 833 10735 867
rect 10793 833 10827 867
rect 11621 833 11655 867
rect 11897 833 11931 867
rect 12081 833 12115 867
rect 14013 833 14047 867
rect 16497 833 16531 867
rect 16865 833 16899 867
rect 18521 833 18555 867
rect 2881 765 2915 799
rect 6285 765 6319 799
rect 6377 765 6411 799
rect 7757 765 7791 799
rect 10885 765 10919 799
rect 12357 765 12391 799
rect 13829 765 13863 799
rect 16221 765 16255 799
rect 18337 697 18371 731
rect 4537 629 4571 663
rect 6837 629 6871 663
rect 9689 629 9723 663
rect 11897 629 11931 663
rect 3157 425 3191 459
rect 3249 425 3283 459
rect 5733 425 5767 459
rect 8493 425 8527 459
rect 10517 425 10551 459
rect 12817 425 12851 459
rect 14749 425 14783 459
rect 15117 425 15151 459
rect 17325 425 17359 459
rect 17693 425 17727 459
rect 18153 425 18187 459
rect 18521 425 18555 459
rect 6101 357 6135 391
rect 3065 289 3099 323
rect 3801 289 3835 323
rect 5365 289 5399 323
rect 6653 289 6687 323
rect 8769 289 8803 323
rect 9137 289 9171 323
rect 10149 289 10183 323
rect 12173 289 12207 323
rect 12541 289 12575 323
rect 12633 289 12667 323
rect 3341 221 3375 255
rect 3709 221 3743 255
rect 3893 221 3927 255
rect 5457 221 5491 255
rect 6469 221 6503 255
rect 8677 221 8711 255
rect 10241 221 10275 255
rect 14657 221 14691 255
rect 14933 221 14967 255
rect 17233 221 17267 255
rect 18061 221 18095 255
rect 6561 153 6595 187
<< metal1 >>
rect 0 10906 18860 10928
rect 0 10854 4660 10906
rect 4712 10854 4724 10906
rect 4776 10854 4788 10906
rect 4840 10854 4852 10906
rect 4904 10854 4916 10906
rect 4968 10854 7760 10906
rect 7812 10854 7824 10906
rect 7876 10854 7888 10906
rect 7940 10854 7952 10906
rect 8004 10854 8016 10906
rect 8068 10854 10860 10906
rect 10912 10854 10924 10906
rect 10976 10854 10988 10906
rect 11040 10854 11052 10906
rect 11104 10854 11116 10906
rect 11168 10854 13960 10906
rect 14012 10854 14024 10906
rect 14076 10854 14088 10906
rect 14140 10854 14152 10906
rect 14204 10854 14216 10906
rect 14268 10854 17060 10906
rect 17112 10854 17124 10906
rect 17176 10854 17188 10906
rect 17240 10854 17252 10906
rect 17304 10854 17316 10906
rect 17368 10854 18860 10906
rect 0 10832 18860 10854
rect 2406 10752 2412 10804
rect 2464 10792 2470 10804
rect 2464 10764 2728 10792
rect 2464 10752 2470 10764
rect 2038 10724 2044 10736
rect 1596 10696 2044 10724
rect 1596 10665 1624 10696
rect 2038 10684 2044 10696
rect 2096 10724 2102 10736
rect 2096 10696 2636 10724
rect 2096 10684 2102 10696
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10625 1639 10659
rect 1581 10619 1639 10625
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2406 10656 2412 10668
rect 2363 10628 2412 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 2406 10616 2412 10628
rect 2464 10616 2470 10668
rect 2608 10665 2636 10696
rect 2700 10665 2728 10764
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 7285 10795 7343 10801
rect 7285 10792 7297 10795
rect 7156 10764 7297 10792
rect 7156 10752 7162 10764
rect 7285 10761 7297 10764
rect 7331 10761 7343 10795
rect 7285 10755 7343 10761
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10413 10795 10471 10801
rect 10413 10792 10425 10795
rect 10008 10764 10425 10792
rect 10008 10752 10014 10764
rect 10413 10761 10425 10764
rect 10459 10761 10471 10795
rect 10413 10755 10471 10761
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 12897 10795 12955 10801
rect 12897 10792 12909 10795
rect 12860 10764 12909 10792
rect 12860 10752 12866 10764
rect 12897 10761 12909 10764
rect 12943 10761 12955 10795
rect 12897 10755 12955 10761
rect 14001 10795 14059 10801
rect 14001 10761 14013 10795
rect 14047 10792 14059 10795
rect 14734 10792 14740 10804
rect 14047 10764 14740 10792
rect 14047 10761 14059 10764
rect 14001 10755 14059 10761
rect 14734 10752 14740 10764
rect 14792 10752 14798 10804
rect 18325 10795 18383 10801
rect 18325 10761 18337 10795
rect 18371 10761 18383 10795
rect 18325 10755 18383 10761
rect 10321 10727 10379 10733
rect 10321 10693 10333 10727
rect 10367 10724 10379 10727
rect 11517 10727 11575 10733
rect 11517 10724 11529 10727
rect 10367 10696 11529 10724
rect 10367 10693 10379 10696
rect 10321 10687 10379 10693
rect 11517 10693 11529 10696
rect 11563 10693 11575 10727
rect 13538 10724 13544 10736
rect 13499 10696 13544 10724
rect 11517 10687 11575 10693
rect 13538 10684 13544 10696
rect 13596 10684 13602 10736
rect 13633 10727 13691 10733
rect 13633 10693 13645 10727
rect 13679 10724 13691 10727
rect 15197 10727 15255 10733
rect 15197 10724 15209 10727
rect 13679 10696 15209 10724
rect 13679 10693 13691 10696
rect 13633 10687 13691 10693
rect 15197 10693 15209 10696
rect 15243 10693 15255 10727
rect 15197 10687 15255 10693
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10625 2651 10659
rect 2593 10619 2651 10625
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10625 2743 10659
rect 2685 10619 2743 10625
rect 2777 10659 2835 10665
rect 2777 10625 2789 10659
rect 2823 10656 2835 10659
rect 2866 10656 2872 10668
rect 2823 10628 2872 10656
rect 2823 10625 2835 10628
rect 2777 10619 2835 10625
rect 2866 10616 2872 10628
rect 2924 10616 2930 10668
rect 7466 10656 7472 10668
rect 7427 10628 7472 10656
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10625 10195 10659
rect 10137 10619 10195 10625
rect 10597 10659 10655 10665
rect 10597 10625 10609 10659
rect 10643 10656 10655 10659
rect 11238 10656 11244 10668
rect 10643 10628 11244 10656
rect 10643 10625 10655 10628
rect 10597 10619 10655 10625
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10557 1731 10591
rect 1673 10551 1731 10557
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10588 2099 10591
rect 2958 10588 2964 10600
rect 2087 10560 2964 10588
rect 2087 10557 2099 10560
rect 2041 10551 2099 10557
rect 566 10412 572 10464
rect 624 10452 630 10464
rect 1397 10455 1455 10461
rect 1397 10452 1409 10455
rect 624 10424 1409 10452
rect 624 10412 630 10424
rect 1397 10421 1409 10424
rect 1443 10421 1455 10455
rect 1688 10452 1716 10551
rect 2958 10548 2964 10560
rect 3016 10548 3022 10600
rect 10152 10520 10180 10619
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 11333 10659 11391 10665
rect 11333 10625 11345 10659
rect 11379 10656 11391 10659
rect 11790 10656 11796 10668
rect 11379 10628 11796 10656
rect 11379 10625 11391 10628
rect 11333 10619 11391 10625
rect 11790 10616 11796 10628
rect 11848 10656 11854 10668
rect 12069 10659 12127 10665
rect 12069 10656 12081 10659
rect 11848 10628 12081 10656
rect 11848 10616 11854 10628
rect 12069 10625 12081 10628
rect 12115 10625 12127 10659
rect 12069 10619 12127 10625
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10656 13139 10659
rect 13127 10628 15056 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 11609 10591 11667 10597
rect 11609 10588 11621 10591
rect 11204 10560 11621 10588
rect 11204 10548 11210 10560
rect 11609 10557 11621 10560
rect 11655 10557 11667 10591
rect 11609 10551 11667 10557
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10588 13415 10591
rect 14642 10588 14648 10600
rect 13403 10560 14648 10588
rect 13403 10557 13415 10560
rect 13357 10551 13415 10557
rect 14642 10548 14648 10560
rect 14700 10548 14706 10600
rect 13722 10520 13728 10532
rect 10152 10492 13728 10520
rect 13722 10480 13728 10492
rect 13780 10480 13786 10532
rect 13906 10480 13912 10532
rect 13964 10520 13970 10532
rect 14461 10523 14519 10529
rect 14461 10520 14473 10523
rect 13964 10492 14473 10520
rect 13964 10480 13970 10492
rect 14461 10489 14473 10492
rect 14507 10489 14519 10523
rect 15028 10520 15056 10628
rect 15102 10616 15108 10668
rect 15160 10656 15166 10668
rect 15160 10628 15205 10656
rect 15160 10616 15166 10628
rect 15286 10616 15292 10668
rect 15344 10656 15350 10668
rect 15381 10659 15439 10665
rect 15381 10656 15393 10659
rect 15344 10628 15393 10656
rect 15344 10616 15350 10628
rect 15381 10625 15393 10628
rect 15427 10625 15439 10659
rect 18046 10656 18052 10668
rect 18007 10628 18052 10656
rect 15381 10619 15439 10625
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 18233 10659 18291 10665
rect 18233 10625 18245 10659
rect 18279 10656 18291 10659
rect 18340 10656 18368 10755
rect 18279 10628 18368 10656
rect 18509 10659 18567 10665
rect 18279 10625 18291 10628
rect 18233 10619 18291 10625
rect 18509 10625 18521 10659
rect 18555 10656 18567 10659
rect 18782 10656 18788 10668
rect 18555 10628 18788 10656
rect 18555 10625 18567 10628
rect 18509 10619 18567 10625
rect 17865 10591 17923 10597
rect 17865 10557 17877 10591
rect 17911 10588 17923 10591
rect 18524 10588 18552 10619
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 17911 10560 18552 10588
rect 17911 10557 17923 10560
rect 17865 10551 17923 10557
rect 18049 10523 18107 10529
rect 18049 10520 18061 10523
rect 15028 10492 18061 10520
rect 14461 10483 14519 10489
rect 18049 10489 18061 10492
rect 18095 10489 18107 10523
rect 18049 10483 18107 10489
rect 2225 10455 2283 10461
rect 2225 10452 2237 10455
rect 1688 10424 2237 10452
rect 1397 10415 1455 10421
rect 2225 10421 2237 10424
rect 2271 10452 2283 10455
rect 2498 10452 2504 10464
rect 2271 10424 2504 10452
rect 2271 10421 2283 10424
rect 2225 10415 2283 10421
rect 2498 10412 2504 10424
rect 2556 10412 2562 10464
rect 11054 10452 11060 10464
rect 11015 10424 11060 10452
rect 11054 10412 11060 10424
rect 11112 10412 11118 10464
rect 11606 10412 11612 10464
rect 11664 10452 11670 10464
rect 12713 10455 12771 10461
rect 12713 10452 12725 10455
rect 11664 10424 12725 10452
rect 11664 10412 11670 10424
rect 12713 10421 12725 10424
rect 12759 10421 12771 10455
rect 12713 10415 12771 10421
rect 14185 10455 14243 10461
rect 14185 10421 14197 10455
rect 14231 10452 14243 10455
rect 14366 10452 14372 10464
rect 14231 10424 14372 10452
rect 14231 10421 14243 10424
rect 14185 10415 14243 10421
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 14826 10412 14832 10464
rect 14884 10452 14890 10464
rect 15013 10455 15071 10461
rect 15013 10452 15025 10455
rect 14884 10424 15025 10452
rect 14884 10412 14890 10424
rect 15013 10421 15025 10424
rect 15059 10421 15071 10455
rect 15013 10415 15071 10421
rect 15933 10455 15991 10461
rect 15933 10421 15945 10455
rect 15979 10452 15991 10455
rect 16206 10452 16212 10464
rect 15979 10424 16212 10452
rect 15979 10421 15991 10424
rect 15933 10415 15991 10421
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 0 10362 18860 10384
rect 0 10310 3110 10362
rect 3162 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 3302 10362
rect 3354 10310 3366 10362
rect 3418 10310 6210 10362
rect 6262 10310 6274 10362
rect 6326 10310 6338 10362
rect 6390 10310 6402 10362
rect 6454 10310 6466 10362
rect 6518 10310 9310 10362
rect 9362 10310 9374 10362
rect 9426 10310 9438 10362
rect 9490 10310 9502 10362
rect 9554 10310 9566 10362
rect 9618 10310 12410 10362
rect 12462 10310 12474 10362
rect 12526 10310 12538 10362
rect 12590 10310 12602 10362
rect 12654 10310 12666 10362
rect 12718 10310 15510 10362
rect 15562 10310 15574 10362
rect 15626 10310 15638 10362
rect 15690 10310 15702 10362
rect 15754 10310 15766 10362
rect 15818 10310 18860 10362
rect 0 10288 18860 10310
rect 1394 10248 1400 10260
rect 1355 10220 1400 10248
rect 1394 10208 1400 10220
rect 1452 10208 1458 10260
rect 4430 10248 4436 10260
rect 2976 10220 4436 10248
rect 2685 10115 2743 10121
rect 2685 10081 2697 10115
rect 2731 10112 2743 10115
rect 2976 10112 3004 10220
rect 4430 10208 4436 10220
rect 4488 10248 4494 10260
rect 5813 10251 5871 10257
rect 5813 10248 5825 10251
rect 4488 10220 5825 10248
rect 4488 10208 4494 10220
rect 5813 10217 5825 10220
rect 5859 10248 5871 10251
rect 5902 10248 5908 10260
rect 5859 10220 5908 10248
rect 5859 10217 5871 10220
rect 5813 10211 5871 10217
rect 5902 10208 5908 10220
rect 5960 10248 5966 10260
rect 6822 10248 6828 10260
rect 5960 10220 6828 10248
rect 5960 10208 5966 10220
rect 6822 10208 6828 10220
rect 6880 10248 6886 10260
rect 6880 10220 7420 10248
rect 6880 10208 6886 10220
rect 3694 10180 3700 10192
rect 2731 10084 3004 10112
rect 3528 10152 3700 10180
rect 2731 10081 2743 10084
rect 2685 10075 2743 10081
rect 1394 10004 1400 10056
rect 1452 10044 1458 10056
rect 1489 10047 1547 10053
rect 1489 10044 1501 10047
rect 1452 10016 1501 10044
rect 1452 10004 1458 10016
rect 1489 10013 1501 10016
rect 1535 10013 1547 10047
rect 2958 10044 2964 10056
rect 2919 10016 2964 10044
rect 1489 10007 1547 10013
rect 2958 10004 2964 10016
rect 3016 10004 3022 10056
rect 3145 10047 3203 10053
rect 3145 10013 3157 10047
rect 3191 10044 3203 10047
rect 3326 10044 3332 10056
rect 3191 10016 3332 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 3326 10004 3332 10016
rect 3384 10004 3390 10056
rect 3528 10053 3556 10152
rect 3694 10140 3700 10152
rect 3752 10140 3758 10192
rect 7392 10180 7420 10220
rect 7466 10208 7472 10260
rect 7524 10248 7530 10260
rect 12986 10248 12992 10260
rect 7524 10220 12992 10248
rect 7524 10208 7530 10220
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 13081 10251 13139 10257
rect 13081 10217 13093 10251
rect 13127 10248 13139 10251
rect 13538 10248 13544 10260
rect 13127 10220 13544 10248
rect 13127 10217 13139 10220
rect 13081 10211 13139 10217
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 17819 10251 17877 10257
rect 17819 10217 17831 10251
rect 17865 10248 17877 10251
rect 18046 10248 18052 10260
rect 17865 10220 18052 10248
rect 17865 10217 17877 10220
rect 17819 10211 17877 10217
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 8113 10183 8171 10189
rect 8113 10180 8125 10183
rect 7392 10152 8125 10180
rect 8113 10149 8125 10152
rect 8159 10180 8171 10183
rect 8297 10183 8355 10189
rect 8297 10180 8309 10183
rect 8159 10152 8309 10180
rect 8159 10149 8171 10152
rect 8113 10143 8171 10149
rect 8297 10149 8309 10152
rect 8343 10149 8355 10183
rect 8297 10143 8355 10149
rect 14918 10140 14924 10192
rect 14976 10180 14982 10192
rect 14976 10152 15792 10180
rect 14976 10140 14982 10152
rect 3970 10112 3976 10124
rect 3804 10084 3976 10112
rect 3513 10047 3571 10053
rect 3513 10013 3525 10047
rect 3559 10013 3571 10047
rect 3513 10007 3571 10013
rect 3697 10047 3755 10053
rect 3697 10013 3709 10047
rect 3743 10044 3755 10047
rect 3804 10044 3832 10084
rect 3970 10072 3976 10084
rect 4028 10112 4034 10124
rect 6086 10112 6092 10124
rect 4028 10084 6092 10112
rect 4028 10072 4034 10084
rect 6086 10072 6092 10084
rect 6144 10112 6150 10124
rect 8481 10115 8539 10121
rect 8481 10112 8493 10115
rect 6144 10084 8493 10112
rect 6144 10072 6150 10084
rect 8481 10081 8493 10084
rect 8527 10081 8539 10115
rect 11330 10112 11336 10124
rect 11243 10084 11336 10112
rect 8481 10075 8539 10081
rect 11330 10072 11336 10084
rect 11388 10112 11394 10124
rect 15010 10112 15016 10124
rect 11388 10084 15016 10112
rect 11388 10072 11394 10084
rect 15010 10072 15016 10084
rect 15068 10072 15074 10124
rect 8846 10044 8852 10056
rect 3743 10016 3832 10044
rect 8807 10016 8852 10044
rect 3743 10013 3755 10016
rect 3697 10007 3755 10013
rect 8846 10004 8852 10016
rect 8904 10004 8910 10056
rect 11054 10044 11060 10056
rect 11015 10016 11060 10044
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 12986 10004 12992 10056
rect 13044 10044 13050 10056
rect 13265 10047 13323 10053
rect 13265 10044 13277 10047
rect 13044 10016 13277 10044
rect 13044 10004 13050 10016
rect 13265 10013 13277 10016
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 13357 10047 13415 10053
rect 13357 10013 13369 10047
rect 13403 10044 13415 10047
rect 13541 10047 13599 10053
rect 13541 10044 13553 10047
rect 13403 10016 13553 10044
rect 13403 10013 13415 10016
rect 13357 10007 13415 10013
rect 13541 10013 13553 10016
rect 13587 10013 13599 10047
rect 13906 10044 13912 10056
rect 13867 10016 13912 10044
rect 13541 10007 13599 10013
rect 13906 10004 13912 10016
rect 13964 10004 13970 10056
rect 15764 10053 15792 10152
rect 16393 10115 16451 10121
rect 16393 10081 16405 10115
rect 16439 10112 16451 10115
rect 16574 10112 16580 10124
rect 16439 10084 16580 10112
rect 16439 10081 16451 10084
rect 16393 10075 16451 10081
rect 16574 10072 16580 10084
rect 16632 10072 16638 10124
rect 15749 10047 15807 10053
rect 15749 10013 15761 10047
rect 15795 10013 15807 10047
rect 15749 10007 15807 10013
rect 15841 10047 15899 10053
rect 15841 10013 15853 10047
rect 15887 10044 15899 10047
rect 16025 10047 16083 10053
rect 16025 10044 16037 10047
rect 15887 10016 16037 10044
rect 15887 10013 15899 10016
rect 15841 10007 15899 10013
rect 16025 10013 16037 10016
rect 16071 10013 16083 10047
rect 16025 10007 16083 10013
rect 18233 10047 18291 10053
rect 18233 10013 18245 10047
rect 18279 10044 18291 10047
rect 18509 10047 18567 10053
rect 18509 10044 18521 10047
rect 18279 10016 18521 10044
rect 18279 10013 18291 10016
rect 18233 10007 18291 10013
rect 18509 10013 18521 10016
rect 18555 10044 18567 10047
rect 18598 10044 18604 10056
rect 18555 10016 18604 10044
rect 18555 10013 18567 10016
rect 18509 10007 18567 10013
rect 18598 10004 18604 10016
rect 18656 10004 18662 10056
rect 3970 9976 3976 9988
rect 3931 9948 3976 9976
rect 3970 9936 3976 9948
rect 4028 9936 4034 9988
rect 4430 9936 4436 9988
rect 4488 9936 4494 9988
rect 6365 9979 6423 9985
rect 6365 9945 6377 9979
rect 6411 9945 6423 9979
rect 6365 9939 6423 9945
rect 3234 9908 3240 9920
rect 3195 9880 3240 9908
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 3418 9908 3424 9920
rect 3379 9880 3424 9908
rect 3418 9868 3424 9880
rect 3476 9868 3482 9920
rect 3694 9868 3700 9920
rect 3752 9908 3758 9920
rect 4154 9908 4160 9920
rect 3752 9880 4160 9908
rect 3752 9868 3758 9880
rect 4154 9868 4160 9880
rect 4212 9908 4218 9920
rect 5258 9908 5264 9920
rect 4212 9880 5264 9908
rect 4212 9868 4218 9880
rect 5258 9868 5264 9880
rect 5316 9908 5322 9920
rect 5445 9911 5503 9917
rect 5445 9908 5457 9911
rect 5316 9880 5457 9908
rect 5316 9868 5322 9880
rect 5445 9877 5457 9880
rect 5491 9877 5503 9911
rect 6380 9908 6408 9939
rect 6822 9936 6828 9988
rect 6880 9936 6886 9988
rect 10597 9979 10655 9985
rect 10597 9976 10609 9979
rect 9890 9962 10609 9976
rect 9876 9948 10609 9962
rect 6546 9908 6552 9920
rect 6380 9880 6552 9908
rect 5445 9871 5503 9877
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 7650 9868 7656 9920
rect 7708 9908 7714 9920
rect 7837 9911 7895 9917
rect 7837 9908 7849 9911
rect 7708 9880 7849 9908
rect 7708 9868 7714 9880
rect 7837 9877 7849 9880
rect 7883 9877 7895 9911
rect 7837 9871 7895 9877
rect 8113 9911 8171 9917
rect 8113 9877 8125 9911
rect 8159 9908 8171 9911
rect 9876 9908 9904 9948
rect 10597 9945 10609 9948
rect 10643 9976 10655 9979
rect 11146 9976 11152 9988
rect 10643 9948 11152 9976
rect 10643 9945 10655 9948
rect 10597 9939 10655 9945
rect 11146 9936 11152 9948
rect 11204 9936 11210 9988
rect 11606 9976 11612 9988
rect 11567 9948 11612 9976
rect 11606 9936 11612 9948
rect 11664 9936 11670 9988
rect 10318 9917 10324 9920
rect 8159 9880 9904 9908
rect 10275 9911 10324 9917
rect 8159 9877 8171 9880
rect 8113 9871 8171 9877
rect 10275 9877 10287 9911
rect 10321 9877 10324 9911
rect 10275 9871 10324 9877
rect 10318 9868 10324 9871
rect 10376 9868 10382 9920
rect 10686 9868 10692 9920
rect 10744 9908 10750 9920
rect 10873 9911 10931 9917
rect 10873 9908 10885 9911
rect 10744 9880 10885 9908
rect 10744 9868 10750 9880
rect 10873 9877 10885 9880
rect 10919 9877 10931 9911
rect 11164 9908 11192 9936
rect 12084 9908 12112 9962
rect 14458 9936 14464 9988
rect 14516 9936 14522 9988
rect 16758 9936 16764 9988
rect 16816 9936 16822 9988
rect 13170 9908 13176 9920
rect 11164 9880 13176 9908
rect 10873 9871 10931 9877
rect 13170 9868 13176 9880
rect 13228 9868 13234 9920
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 15335 9911 15393 9917
rect 15335 9908 15347 9911
rect 15252 9880 15347 9908
rect 15252 9868 15258 9880
rect 15335 9877 15347 9880
rect 15381 9877 15393 9911
rect 18322 9908 18328 9920
rect 18283 9880 18328 9908
rect 15335 9871 15393 9877
rect 18322 9868 18328 9880
rect 18380 9868 18386 9920
rect 0 9818 18860 9840
rect 0 9766 4660 9818
rect 4712 9766 4724 9818
rect 4776 9766 4788 9818
rect 4840 9766 4852 9818
rect 4904 9766 4916 9818
rect 4968 9766 7760 9818
rect 7812 9766 7824 9818
rect 7876 9766 7888 9818
rect 7940 9766 7952 9818
rect 8004 9766 8016 9818
rect 8068 9766 10860 9818
rect 10912 9766 10924 9818
rect 10976 9766 10988 9818
rect 11040 9766 11052 9818
rect 11104 9766 11116 9818
rect 11168 9766 13960 9818
rect 14012 9766 14024 9818
rect 14076 9766 14088 9818
rect 14140 9766 14152 9818
rect 14204 9766 14216 9818
rect 14268 9766 17060 9818
rect 17112 9766 17124 9818
rect 17176 9766 17188 9818
rect 17240 9766 17252 9818
rect 17304 9766 17316 9818
rect 17368 9766 18860 9818
rect 0 9744 18860 9766
rect 2038 9704 2044 9716
rect 1999 9676 2044 9704
rect 2038 9664 2044 9676
rect 2096 9664 2102 9716
rect 2590 9704 2596 9716
rect 2148 9676 2596 9704
rect 566 9636 572 9648
rect 527 9608 572 9636
rect 566 9596 572 9608
rect 624 9596 630 9648
rect 2148 9636 2176 9676
rect 2590 9664 2596 9676
rect 2648 9664 2654 9716
rect 2685 9707 2743 9713
rect 2685 9673 2697 9707
rect 2731 9704 2743 9707
rect 2774 9704 2780 9716
rect 2731 9676 2780 9704
rect 2731 9673 2743 9676
rect 2685 9667 2743 9673
rect 2774 9664 2780 9676
rect 2832 9704 2838 9716
rect 3418 9704 3424 9716
rect 2832 9676 3424 9704
rect 2832 9664 2838 9676
rect 3418 9664 3424 9676
rect 3476 9664 3482 9716
rect 3694 9664 3700 9716
rect 3752 9664 3758 9716
rect 3973 9707 4031 9713
rect 3973 9704 3985 9707
rect 3804 9676 3985 9704
rect 1794 9608 2176 9636
rect 2225 9639 2283 9645
rect 2225 9605 2237 9639
rect 2271 9636 2283 9639
rect 2271 9608 2820 9636
rect 2271 9605 2283 9608
rect 2225 9599 2283 9605
rect 2130 9568 2136 9580
rect 2091 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9537 2375 9571
rect 2498 9568 2504 9580
rect 2459 9540 2504 9568
rect 2317 9531 2375 9537
rect 290 9500 296 9512
rect 251 9472 296 9500
rect 290 9460 296 9472
rect 348 9460 354 9512
rect 2038 9460 2044 9512
rect 2096 9500 2102 9512
rect 2332 9500 2360 9531
rect 2498 9528 2504 9540
rect 2556 9528 2562 9580
rect 2792 9577 2820 9608
rect 3510 9596 3516 9648
rect 3568 9636 3574 9648
rect 3712 9636 3740 9664
rect 3568 9608 3740 9636
rect 3568 9596 3574 9608
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9537 2835 9571
rect 2958 9568 2964 9580
rect 2919 9540 2964 9568
rect 2777 9531 2835 9537
rect 2958 9528 2964 9540
rect 3016 9528 3022 9580
rect 3694 9568 3700 9580
rect 3655 9540 3700 9568
rect 3694 9528 3700 9540
rect 3752 9528 3758 9580
rect 2096 9472 2360 9500
rect 2096 9460 2102 9472
rect 3326 9460 3332 9512
rect 3384 9500 3390 9512
rect 3804 9500 3832 9676
rect 3973 9673 3985 9676
rect 4019 9673 4031 9707
rect 3973 9667 4031 9673
rect 4062 9664 4068 9716
rect 4120 9704 4126 9716
rect 4120 9676 5212 9704
rect 4120 9664 4126 9676
rect 5184 9648 5212 9676
rect 7650 9664 7656 9716
rect 7708 9664 7714 9716
rect 8570 9704 8576 9716
rect 8531 9676 8576 9704
rect 8570 9664 8576 9676
rect 8628 9664 8634 9716
rect 11790 9704 11796 9716
rect 11751 9676 11796 9704
rect 11790 9664 11796 9676
rect 11848 9664 11854 9716
rect 12986 9664 12992 9716
rect 13044 9704 13050 9716
rect 14918 9704 14924 9716
rect 13044 9676 14924 9704
rect 13044 9664 13050 9676
rect 14918 9664 14924 9676
rect 14976 9664 14982 9716
rect 4985 9639 5043 9645
rect 4985 9636 4997 9639
rect 3896 9608 4997 9636
rect 3896 9577 3924 9608
rect 4985 9605 4997 9608
rect 5031 9605 5043 9639
rect 4985 9599 5043 9605
rect 5166 9596 5172 9648
rect 5224 9596 5230 9648
rect 5902 9596 5908 9648
rect 5960 9636 5966 9648
rect 7668 9636 7696 9664
rect 10318 9636 10324 9648
rect 5960 9608 6118 9636
rect 7668 9608 9352 9636
rect 5960 9596 5966 9608
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9537 3939 9571
rect 3881 9531 3939 9537
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9568 4399 9571
rect 4798 9568 4804 9580
rect 4387 9540 4804 9568
rect 4387 9537 4399 9540
rect 4341 9531 4399 9537
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9568 5135 9571
rect 5258 9568 5264 9580
rect 5123 9540 5264 9568
rect 5123 9537 5135 9540
rect 5077 9531 5135 9537
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 9324 9577 9352 9608
rect 9508 9608 10324 9636
rect 9508 9577 9536 9608
rect 10318 9596 10324 9608
rect 10376 9596 10382 9648
rect 11330 9636 11336 9648
rect 10428 9608 11336 9636
rect 7653 9571 7711 9577
rect 7653 9568 7665 9571
rect 7576 9540 7665 9568
rect 3384 9472 3832 9500
rect 3384 9460 3390 9472
rect 3970 9460 3976 9512
rect 4028 9500 4034 9512
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 4028 9472 4445 9500
rect 4028 9460 4034 9472
rect 4433 9469 4445 9472
rect 4479 9469 4491 9503
rect 4433 9463 4491 9469
rect 4522 9460 4528 9512
rect 4580 9500 4586 9512
rect 5353 9503 5411 9509
rect 4580 9472 4625 9500
rect 4580 9460 4586 9472
rect 5353 9469 5365 9503
rect 5399 9469 5411 9503
rect 5626 9500 5632 9512
rect 5587 9472 5632 9500
rect 5353 9463 5411 9469
rect 3050 9432 3056 9444
rect 1964 9404 3056 9432
rect 750 9324 756 9376
rect 808 9364 814 9376
rect 1964 9364 1992 9404
rect 3050 9392 3056 9404
rect 3108 9392 3114 9444
rect 808 9336 1992 9364
rect 808 9324 814 9336
rect 2590 9324 2596 9376
rect 2648 9364 2654 9376
rect 3145 9367 3203 9373
rect 3145 9364 3157 9367
rect 2648 9336 3157 9364
rect 2648 9324 2654 9336
rect 3145 9333 3157 9336
rect 3191 9364 3203 9367
rect 3510 9364 3516 9376
rect 3191 9336 3516 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 3789 9367 3847 9373
rect 3789 9364 3801 9367
rect 3660 9336 3801 9364
rect 3660 9324 3666 9336
rect 3789 9333 3801 9336
rect 3835 9333 3847 9367
rect 5258 9364 5264 9376
rect 5219 9336 5264 9364
rect 3789 9327 3847 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5368 9364 5396 9463
rect 5626 9460 5632 9472
rect 5684 9460 5690 9512
rect 7101 9435 7159 9441
rect 7101 9401 7113 9435
rect 7147 9432 7159 9435
rect 7190 9432 7196 9444
rect 7147 9404 7196 9432
rect 7147 9401 7159 9404
rect 7101 9395 7159 9401
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 7576 9432 7604 9540
rect 7653 9537 7665 9540
rect 7699 9537 7711 9571
rect 8665 9571 8723 9577
rect 8665 9568 8677 9571
rect 7653 9531 7711 9537
rect 7760 9540 8677 9568
rect 7760 9512 7788 9540
rect 8665 9537 8677 9540
rect 8711 9537 8723 9571
rect 8665 9531 8723 9537
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 9674 9528 9680 9580
rect 9732 9568 9738 9580
rect 10428 9577 10456 9608
rect 11330 9596 11336 9608
rect 11388 9596 11394 9648
rect 11606 9596 11612 9648
rect 11664 9636 11670 9648
rect 14366 9636 14372 9648
rect 11664 9608 14372 9636
rect 11664 9596 11670 9608
rect 14366 9596 14372 9608
rect 14424 9596 14430 9648
rect 16206 9596 16212 9648
rect 16264 9596 16270 9648
rect 16574 9596 16580 9648
rect 16632 9645 16638 9648
rect 16632 9639 16681 9645
rect 16632 9605 16635 9639
rect 16669 9605 16681 9639
rect 16632 9599 16681 9605
rect 16632 9596 16638 9599
rect 10686 9577 10692 9580
rect 10045 9571 10103 9577
rect 10045 9568 10057 9571
rect 9732 9540 10057 9568
rect 9732 9528 9738 9540
rect 10045 9537 10057 9540
rect 10091 9537 10103 9571
rect 10045 9531 10103 9537
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9537 10471 9571
rect 10680 9568 10692 9577
rect 10647 9540 10692 9568
rect 10413 9531 10471 9537
rect 10680 9531 10692 9540
rect 10686 9528 10692 9531
rect 10744 9528 10750 9580
rect 12529 9571 12587 9577
rect 12529 9537 12541 9571
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 7742 9460 7748 9512
rect 7800 9500 7806 9512
rect 7929 9503 7987 9509
rect 7800 9472 7845 9500
rect 7800 9460 7806 9472
rect 7929 9469 7941 9503
rect 7975 9500 7987 9503
rect 8110 9500 8116 9512
rect 7975 9472 8116 9500
rect 7975 9469 7987 9472
rect 7929 9463 7987 9469
rect 8110 9460 8116 9472
rect 8168 9500 8174 9512
rect 8849 9503 8907 9509
rect 8168 9472 8340 9500
rect 8168 9460 8174 9472
rect 8205 9435 8263 9441
rect 8205 9432 8217 9435
rect 7576 9404 8217 9432
rect 8205 9401 8217 9404
rect 8251 9401 8263 9435
rect 8205 9395 8263 9401
rect 6086 9364 6092 9376
rect 5368 9336 6092 9364
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 7282 9364 7288 9376
rect 7243 9336 7288 9364
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 8312 9364 8340 9472
rect 8849 9469 8861 9503
rect 8895 9500 8907 9503
rect 8938 9500 8944 9512
rect 8895 9472 8944 9500
rect 8895 9469 8907 9472
rect 8849 9463 8907 9469
rect 8938 9460 8944 9472
rect 8996 9460 9002 9512
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9500 9459 9503
rect 9953 9503 10011 9509
rect 9953 9500 9965 9503
rect 9447 9472 9965 9500
rect 9447 9469 9459 9472
rect 9401 9463 9459 9469
rect 9953 9469 9965 9472
rect 9999 9469 10011 9503
rect 9953 9463 10011 9469
rect 8570 9392 8576 9444
rect 8628 9432 8634 9444
rect 9677 9435 9735 9441
rect 9677 9432 9689 9435
rect 8628 9404 9689 9432
rect 8628 9392 8634 9404
rect 9677 9401 9689 9404
rect 9723 9401 9735 9435
rect 9677 9395 9735 9401
rect 10686 9364 10692 9376
rect 8312 9336 10692 9364
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 12544 9364 12572 9531
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 13780 9540 14289 9568
rect 13780 9528 13786 9540
rect 14277 9537 14289 9540
rect 14323 9568 14335 9571
rect 15286 9568 15292 9580
rect 14323 9540 15292 9568
rect 14323 9537 14335 9540
rect 14277 9531 14335 9537
rect 15286 9528 15292 9540
rect 15344 9528 15350 9580
rect 16224 9568 16252 9596
rect 16758 9568 16764 9580
rect 16224 9540 16764 9568
rect 16758 9528 16764 9540
rect 16816 9528 16822 9580
rect 14826 9500 14832 9512
rect 14787 9472 14832 9500
rect 14826 9460 14832 9472
rect 14884 9460 14890 9512
rect 15194 9500 15200 9512
rect 15155 9472 15200 9500
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 14366 9392 14372 9444
rect 14424 9432 14430 9444
rect 14424 9404 14872 9432
rect 14424 9392 14430 9404
rect 12802 9364 12808 9376
rect 12483 9336 12808 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 13170 9324 13176 9376
rect 13228 9364 13234 9376
rect 13722 9364 13728 9376
rect 13228 9336 13728 9364
rect 13228 9324 13234 9336
rect 13722 9324 13728 9336
rect 13780 9364 13786 9376
rect 14458 9364 14464 9376
rect 13780 9336 14464 9364
rect 13780 9324 13786 9336
rect 14458 9324 14464 9336
rect 14516 9364 14522 9376
rect 14645 9367 14703 9373
rect 14645 9364 14657 9367
rect 14516 9336 14657 9364
rect 14516 9324 14522 9336
rect 14645 9333 14657 9336
rect 14691 9333 14703 9367
rect 14844 9364 14872 9404
rect 17494 9364 17500 9376
rect 14844 9336 17500 9364
rect 14645 9327 14703 9333
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 0 9274 18860 9296
rect 0 9222 3110 9274
rect 3162 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 3302 9274
rect 3354 9222 3366 9274
rect 3418 9222 6210 9274
rect 6262 9222 6274 9274
rect 6326 9222 6338 9274
rect 6390 9222 6402 9274
rect 6454 9222 6466 9274
rect 6518 9222 9310 9274
rect 9362 9222 9374 9274
rect 9426 9222 9438 9274
rect 9490 9222 9502 9274
rect 9554 9222 9566 9274
rect 9618 9222 12410 9274
rect 12462 9222 12474 9274
rect 12526 9222 12538 9274
rect 12590 9222 12602 9274
rect 12654 9222 12666 9274
rect 12718 9222 15510 9274
rect 15562 9222 15574 9274
rect 15626 9222 15638 9274
rect 15690 9222 15702 9274
rect 15754 9222 15766 9274
rect 15818 9222 18860 9274
rect 0 9200 18860 9222
rect 2406 9160 2412 9172
rect 2148 9132 2412 9160
rect 2148 9101 2176 9132
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 2777 9163 2835 9169
rect 2777 9129 2789 9163
rect 2823 9160 2835 9163
rect 3694 9160 3700 9172
rect 2823 9132 3700 9160
rect 2823 9129 2835 9132
rect 2777 9123 2835 9129
rect 2133 9095 2191 9101
rect 2133 9061 2145 9095
rect 2179 9061 2191 9095
rect 2133 9055 2191 9061
rect 2225 9095 2283 9101
rect 2225 9061 2237 9095
rect 2271 9092 2283 9095
rect 2501 9095 2559 9101
rect 2501 9092 2513 9095
rect 2271 9064 2513 9092
rect 2271 9061 2283 9064
rect 2225 9055 2283 9061
rect 2501 9061 2513 9064
rect 2547 9061 2559 9095
rect 2501 9055 2559 9061
rect 2317 9027 2375 9033
rect 2317 8993 2329 9027
rect 2363 9024 2375 9027
rect 2774 9024 2780 9036
rect 2363 8996 2780 9024
rect 2363 8993 2375 8996
rect 2317 8987 2375 8993
rect 2774 8984 2780 8996
rect 2832 8984 2838 9036
rect 290 8916 296 8968
rect 348 8956 354 8968
rect 569 8959 627 8965
rect 569 8956 581 8959
rect 348 8928 581 8956
rect 348 8916 354 8928
rect 569 8925 581 8928
rect 615 8956 627 8959
rect 750 8956 756 8968
rect 615 8928 756 8956
rect 615 8925 627 8928
rect 569 8919 627 8925
rect 750 8916 756 8928
rect 808 8916 814 8968
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8956 1823 8959
rect 2038 8956 2044 8968
rect 1811 8928 2044 8956
rect 1811 8925 1823 8928
rect 1765 8919 1823 8925
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8925 2651 8959
rect 2593 8919 2651 8925
rect 2608 8888 2636 8919
rect 2682 8916 2688 8968
rect 2740 8956 2746 8968
rect 2740 8928 2785 8956
rect 2740 8916 2746 8928
rect 2884 8888 2912 9132
rect 3694 9120 3700 9132
rect 3752 9120 3758 9172
rect 4798 9120 4804 9172
rect 4856 9160 4862 9172
rect 4856 9132 5580 9160
rect 4856 9120 4862 9132
rect 3160 9064 5120 9092
rect 2958 8984 2964 9036
rect 3016 9024 3022 9036
rect 3160 9033 3188 9064
rect 3145 9027 3203 9033
rect 3145 9024 3157 9027
rect 3016 8996 3157 9024
rect 3016 8984 3022 8996
rect 3145 8993 3157 8996
rect 3191 8993 3203 9027
rect 4154 9024 4160 9036
rect 3145 8987 3203 8993
rect 3252 8996 3464 9024
rect 3050 8916 3056 8968
rect 3108 8956 3114 8968
rect 3252 8956 3280 8996
rect 3108 8928 3280 8956
rect 3329 8959 3387 8965
rect 3108 8916 3114 8928
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 2608 8860 2912 8888
rect 290 8780 296 8832
rect 348 8820 354 8832
rect 477 8823 535 8829
rect 477 8820 489 8823
rect 348 8792 489 8820
rect 348 8780 354 8792
rect 477 8789 489 8792
rect 523 8789 535 8823
rect 477 8783 535 8789
rect 658 8780 664 8832
rect 716 8820 722 8832
rect 2317 8823 2375 8829
rect 2317 8820 2329 8823
rect 716 8792 2329 8820
rect 716 8780 722 8792
rect 2317 8789 2329 8792
rect 2363 8789 2375 8823
rect 2317 8783 2375 8789
rect 2682 8780 2688 8832
rect 2740 8820 2746 8832
rect 3344 8820 3372 8919
rect 3436 8888 3464 8996
rect 3528 8996 4160 9024
rect 3528 8965 3556 8996
rect 4154 8984 4160 8996
rect 4212 8984 4218 9036
rect 4798 9024 4804 9036
rect 4759 8996 4804 9024
rect 4798 8984 4804 8996
rect 4856 8984 4862 9036
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8925 3571 8959
rect 3513 8919 3571 8925
rect 3602 8916 3608 8968
rect 3660 8956 3666 8968
rect 5092 8965 5120 9064
rect 5552 9024 5580 9132
rect 5626 9120 5632 9172
rect 5684 9160 5690 9172
rect 6273 9163 6331 9169
rect 6273 9160 6285 9163
rect 5684 9132 6285 9160
rect 5684 9120 5690 9132
rect 6273 9129 6285 9132
rect 6319 9129 6331 9163
rect 7742 9160 7748 9172
rect 6273 9123 6331 9129
rect 6380 9132 7748 9160
rect 5810 9052 5816 9104
rect 5868 9092 5874 9104
rect 6380 9092 6408 9132
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 8846 9120 8852 9172
rect 8904 9160 8910 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 8904 9132 9045 9160
rect 8904 9120 8910 9132
rect 9033 9129 9045 9132
rect 9079 9129 9091 9163
rect 9033 9123 9091 9129
rect 11238 9120 11244 9172
rect 11296 9160 11302 9172
rect 12345 9163 12403 9169
rect 12345 9160 12357 9163
rect 11296 9132 12357 9160
rect 11296 9120 11302 9132
rect 12345 9129 12357 9132
rect 12391 9129 12403 9163
rect 12345 9123 12403 9129
rect 12894 9120 12900 9172
rect 12952 9160 12958 9172
rect 18322 9160 18328 9172
rect 12952 9132 18328 9160
rect 12952 9120 12958 9132
rect 18322 9120 18328 9132
rect 18380 9120 18386 9172
rect 8754 9092 8760 9104
rect 5868 9064 6408 9092
rect 6472 9064 8760 9092
rect 5868 9052 5874 9064
rect 6472 9036 6500 9064
rect 8754 9052 8760 9064
rect 8812 9052 8818 9104
rect 8938 9052 8944 9104
rect 8996 9092 9002 9104
rect 8996 9064 10456 9092
rect 8996 9052 9002 9064
rect 10428 9036 10456 9064
rect 12912 9064 13400 9092
rect 6454 9024 6460 9036
rect 5552 8996 6460 9024
rect 6454 8984 6460 8996
rect 6512 8984 6518 9036
rect 6549 9027 6607 9033
rect 6549 8993 6561 9027
rect 6595 9024 6607 9027
rect 7282 9024 7288 9036
rect 6595 8996 7288 9024
rect 6595 8993 6607 8996
rect 6549 8987 6607 8993
rect 7282 8984 7288 8996
rect 7340 8984 7346 9036
rect 9674 9024 9680 9036
rect 8772 8996 9680 9024
rect 4525 8959 4583 8965
rect 4525 8956 4537 8959
rect 3660 8928 4537 8956
rect 3660 8916 3666 8928
rect 4525 8925 4537 8928
rect 4571 8925 4583 8959
rect 4525 8919 4583 8925
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8956 4767 8959
rect 4893 8959 4951 8965
rect 4893 8956 4905 8959
rect 4755 8928 4905 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 4893 8925 4905 8928
rect 4939 8925 4951 8959
rect 4893 8919 4951 8925
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5350 8956 5356 8968
rect 5123 8928 5356 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 3786 8888 3792 8900
rect 3436 8860 3792 8888
rect 3786 8848 3792 8860
rect 3844 8848 3850 8900
rect 4908 8888 4936 8919
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 7006 8956 7012 8968
rect 6967 8928 7012 8956
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 7190 8916 7196 8968
rect 7248 8956 7254 8968
rect 8772 8965 8800 8996
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 9950 8984 9956 9036
rect 10008 9024 10014 9036
rect 10229 9027 10287 9033
rect 10229 9024 10241 9027
rect 10008 8996 10241 9024
rect 10008 8984 10014 8996
rect 10229 8993 10241 8996
rect 10275 8993 10287 9027
rect 10229 8987 10287 8993
rect 10410 8984 10416 9036
rect 10468 9024 10474 9036
rect 11701 9027 11759 9033
rect 11701 9024 11713 9027
rect 10468 8996 11713 9024
rect 10468 8984 10474 8996
rect 11701 8993 11713 8996
rect 11747 8993 11759 9027
rect 11701 8987 11759 8993
rect 8757 8959 8815 8965
rect 8757 8956 8769 8959
rect 7248 8928 8769 8956
rect 7248 8916 7254 8928
rect 4982 8888 4988 8900
rect 4895 8860 4988 8888
rect 4982 8848 4988 8860
rect 5040 8888 5046 8900
rect 5721 8891 5779 8897
rect 5721 8888 5733 8891
rect 5040 8860 5733 8888
rect 5040 8848 5046 8860
rect 5721 8857 5733 8860
rect 5767 8857 5779 8891
rect 5721 8851 5779 8857
rect 5905 8891 5963 8897
rect 5905 8857 5917 8891
rect 5951 8888 5963 8891
rect 7024 8888 7052 8916
rect 7300 8897 7328 8928
rect 8757 8925 8769 8928
rect 8803 8925 8815 8959
rect 8757 8919 8815 8925
rect 8846 8916 8852 8968
rect 8904 8956 8910 8968
rect 9217 8959 9275 8965
rect 9217 8956 9229 8959
rect 8904 8928 9229 8956
rect 8904 8916 8910 8928
rect 9217 8925 9229 8928
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 9306 8916 9312 8968
rect 9364 8956 9370 8968
rect 9766 8956 9772 8968
rect 9364 8928 9409 8956
rect 9727 8928 9772 8956
rect 9364 8916 9370 8928
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 10045 8959 10103 8965
rect 10045 8925 10057 8959
rect 10091 8956 10103 8959
rect 10318 8956 10324 8968
rect 10091 8928 10324 8956
rect 10091 8925 10103 8928
rect 10045 8919 10103 8925
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 11606 8956 11612 8968
rect 11567 8928 11612 8956
rect 11606 8916 11612 8928
rect 11664 8916 11670 8968
rect 12713 8959 12771 8965
rect 12713 8925 12725 8959
rect 12759 8956 12771 8959
rect 12912 8956 12940 9064
rect 12989 9027 13047 9033
rect 12989 8993 13001 9027
rect 13035 9024 13047 9027
rect 13372 9024 13400 9064
rect 14734 9024 14740 9036
rect 13035 8996 13308 9024
rect 13372 8996 14740 9024
rect 13035 8993 13047 8996
rect 12989 8987 13047 8993
rect 12759 8928 12940 8956
rect 12759 8925 12771 8928
rect 12713 8919 12771 8925
rect 5951 8860 7052 8888
rect 7101 8891 7159 8897
rect 5951 8857 5963 8860
rect 5905 8851 5963 8857
rect 7101 8857 7113 8891
rect 7147 8857 7159 8891
rect 7101 8851 7159 8857
rect 7285 8891 7343 8897
rect 7285 8857 7297 8891
rect 7331 8857 7343 8891
rect 9861 8891 9919 8897
rect 9861 8888 9873 8891
rect 7285 8851 7343 8857
rect 7484 8860 9873 8888
rect 2740 8792 3372 8820
rect 3421 8823 3479 8829
rect 2740 8780 2746 8792
rect 3421 8789 3433 8823
rect 3467 8820 3479 8823
rect 3878 8820 3884 8832
rect 3467 8792 3884 8820
rect 3467 8789 3479 8792
rect 3421 8783 3479 8789
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 4522 8780 4528 8832
rect 4580 8820 4586 8832
rect 4617 8823 4675 8829
rect 4617 8820 4629 8823
rect 4580 8792 4629 8820
rect 4580 8780 4586 8792
rect 4617 8789 4629 8792
rect 4663 8820 4675 8823
rect 5074 8820 5080 8832
rect 4663 8792 5080 8820
rect 4663 8789 4675 8792
rect 4617 8783 4675 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 6917 8823 6975 8829
rect 6917 8789 6929 8823
rect 6963 8820 6975 8823
rect 7009 8823 7067 8829
rect 7009 8820 7021 8823
rect 6963 8792 7021 8820
rect 6963 8789 6975 8792
rect 6917 8783 6975 8789
rect 7009 8789 7021 8792
rect 7055 8789 7067 8823
rect 7116 8820 7144 8851
rect 7374 8820 7380 8832
rect 7116 8792 7380 8820
rect 7009 8783 7067 8789
rect 7374 8780 7380 8792
rect 7432 8820 7438 8832
rect 7484 8820 7512 8860
rect 9861 8857 9873 8860
rect 9907 8888 9919 8891
rect 10502 8888 10508 8900
rect 9907 8860 10508 8888
rect 9907 8857 9919 8860
rect 9861 8851 9919 8857
rect 10502 8848 10508 8860
rect 10560 8848 10566 8900
rect 11517 8891 11575 8897
rect 11517 8888 11529 8891
rect 10704 8860 11529 8888
rect 8846 8820 8852 8832
rect 7432 8792 7512 8820
rect 8807 8792 8852 8820
rect 7432 8780 7438 8792
rect 8846 8780 8852 8792
rect 8904 8780 8910 8832
rect 10704 8829 10732 8860
rect 11517 8857 11529 8860
rect 11563 8857 11575 8891
rect 11517 8851 11575 8857
rect 9677 8823 9735 8829
rect 9677 8789 9689 8823
rect 9723 8820 9735 8823
rect 9769 8823 9827 8829
rect 9769 8820 9781 8823
rect 9723 8792 9781 8820
rect 9723 8789 9735 8792
rect 9677 8783 9735 8789
rect 9769 8789 9781 8792
rect 9815 8789 9827 8823
rect 9769 8783 9827 8789
rect 10689 8823 10747 8829
rect 10689 8789 10701 8823
rect 10735 8789 10747 8823
rect 10689 8783 10747 8789
rect 11149 8823 11207 8829
rect 11149 8789 11161 8823
rect 11195 8820 11207 8823
rect 11238 8820 11244 8832
rect 11195 8792 11244 8820
rect 11195 8789 11207 8792
rect 11149 8783 11207 8789
rect 11238 8780 11244 8792
rect 11296 8780 11302 8832
rect 12250 8820 12256 8832
rect 12211 8792 12256 8820
rect 12250 8780 12256 8792
rect 12308 8780 12314 8832
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 13280 8829 13308 8996
rect 14734 8984 14740 8996
rect 14792 8984 14798 9036
rect 15010 9024 15016 9036
rect 14971 8996 15016 9024
rect 15010 8984 15016 8996
rect 15068 8984 15074 9036
rect 15102 8916 15108 8968
rect 15160 8956 15166 8968
rect 15841 8959 15899 8965
rect 15841 8956 15853 8959
rect 15160 8928 15853 8956
rect 15160 8916 15166 8928
rect 15841 8925 15853 8928
rect 15887 8925 15899 8959
rect 15841 8919 15899 8925
rect 13722 8848 13728 8900
rect 13780 8848 13786 8900
rect 14642 8848 14648 8900
rect 14700 8888 14706 8900
rect 14737 8891 14795 8897
rect 14737 8888 14749 8891
rect 14700 8860 14749 8888
rect 14700 8848 14706 8860
rect 14737 8857 14749 8860
rect 14783 8888 14795 8891
rect 14826 8888 14832 8900
rect 14783 8860 14832 8888
rect 14783 8857 14795 8860
rect 14737 8851 14795 8857
rect 14826 8848 14832 8860
rect 14884 8848 14890 8900
rect 15010 8888 15016 8900
rect 14936 8860 15016 8888
rect 12805 8823 12863 8829
rect 12805 8820 12817 8823
rect 12584 8792 12817 8820
rect 12584 8780 12590 8792
rect 12805 8789 12817 8792
rect 12851 8789 12863 8823
rect 12805 8783 12863 8789
rect 13265 8823 13323 8829
rect 13265 8789 13277 8823
rect 13311 8820 13323 8823
rect 14458 8820 14464 8832
rect 13311 8792 14464 8820
rect 13311 8789 13323 8792
rect 13265 8783 13323 8789
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 14550 8780 14556 8832
rect 14608 8820 14614 8832
rect 14936 8820 14964 8860
rect 15010 8848 15016 8860
rect 15068 8888 15074 8900
rect 16114 8888 16120 8900
rect 15068 8860 15792 8888
rect 16075 8860 16120 8888
rect 15068 8848 15074 8860
rect 14608 8792 14964 8820
rect 15197 8823 15255 8829
rect 14608 8780 14614 8792
rect 15197 8789 15209 8823
rect 15243 8820 15255 8823
rect 15286 8820 15292 8832
rect 15243 8792 15292 8820
rect 15243 8789 15255 8792
rect 15197 8783 15255 8789
rect 15286 8780 15292 8792
rect 15344 8820 15350 8832
rect 15657 8823 15715 8829
rect 15657 8820 15669 8823
rect 15344 8792 15669 8820
rect 15344 8780 15350 8792
rect 15657 8789 15669 8792
rect 15703 8789 15715 8823
rect 15764 8820 15792 8860
rect 16114 8848 16120 8860
rect 16172 8848 16178 8900
rect 16758 8848 16764 8900
rect 16816 8848 16822 8900
rect 17865 8891 17923 8897
rect 17865 8857 17877 8891
rect 17911 8857 17923 8891
rect 17865 8851 17923 8857
rect 17880 8820 17908 8851
rect 15764 8792 17908 8820
rect 15657 8783 15715 8789
rect 0 8730 18860 8752
rect 0 8678 4660 8730
rect 4712 8678 4724 8730
rect 4776 8678 4788 8730
rect 4840 8678 4852 8730
rect 4904 8678 4916 8730
rect 4968 8678 7760 8730
rect 7812 8678 7824 8730
rect 7876 8678 7888 8730
rect 7940 8678 7952 8730
rect 8004 8678 8016 8730
rect 8068 8678 10860 8730
rect 10912 8678 10924 8730
rect 10976 8678 10988 8730
rect 11040 8678 11052 8730
rect 11104 8678 11116 8730
rect 11168 8678 13960 8730
rect 14012 8678 14024 8730
rect 14076 8678 14088 8730
rect 14140 8678 14152 8730
rect 14204 8678 14216 8730
rect 14268 8678 17060 8730
rect 17112 8678 17124 8730
rect 17176 8678 17188 8730
rect 17240 8678 17252 8730
rect 17304 8678 17316 8730
rect 17368 8678 18860 8730
rect 0 8656 18860 8678
rect 2130 8625 2136 8628
rect 2087 8619 2136 8625
rect 2087 8616 2099 8619
rect 2043 8588 2099 8616
rect 2087 8585 2099 8588
rect 2133 8585 2136 8619
rect 2087 8579 2136 8585
rect 2130 8576 2136 8579
rect 2188 8616 2194 8628
rect 2682 8616 2688 8628
rect 2188 8588 2688 8616
rect 2188 8576 2194 8588
rect 2682 8576 2688 8588
rect 2740 8576 2746 8628
rect 4893 8619 4951 8625
rect 4893 8585 4905 8619
rect 4939 8616 4951 8619
rect 4982 8616 4988 8628
rect 4939 8588 4988 8616
rect 4939 8585 4951 8588
rect 4893 8579 4951 8585
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 6457 8619 6515 8625
rect 6457 8585 6469 8619
rect 6503 8616 6515 8619
rect 6546 8616 6552 8628
rect 6503 8588 6552 8616
rect 6503 8585 6515 8588
rect 6457 8579 6515 8585
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8616 7159 8619
rect 7285 8619 7343 8625
rect 7285 8616 7297 8619
rect 7147 8588 7297 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 7285 8585 7297 8588
rect 7331 8585 7343 8619
rect 7285 8579 7343 8585
rect 7484 8588 8892 8616
rect 5537 8551 5595 8557
rect 290 8480 296 8492
rect 251 8452 296 8480
rect 290 8440 296 8452
rect 348 8440 354 8492
rect 658 8480 664 8492
rect 619 8452 664 8480
rect 658 8440 664 8452
rect 716 8440 722 8492
rect 1688 8276 1716 8534
rect 4172 8520 5304 8548
rect 2866 8480 2872 8492
rect 2827 8452 2872 8480
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3878 8480 3884 8492
rect 3099 8452 3740 8480
rect 3839 8452 3884 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 3712 8344 3740 8452
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 4172 8489 4200 8520
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8449 4215 8483
rect 4157 8443 4215 8449
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8480 4307 8483
rect 5166 8480 5172 8492
rect 4295 8478 5028 8480
rect 5092 8478 5172 8480
rect 4295 8452 5172 8478
rect 4295 8449 4307 8452
rect 5000 8450 5120 8452
rect 4249 8443 4307 8449
rect 5166 8440 5172 8452
rect 5224 8440 5230 8492
rect 3970 8412 3976 8424
rect 3883 8384 3976 8412
rect 3970 8372 3976 8384
rect 4028 8412 4034 8424
rect 4893 8415 4951 8421
rect 4893 8412 4905 8415
rect 4028 8384 4905 8412
rect 4028 8372 4034 8384
rect 4893 8381 4905 8384
rect 4939 8381 4951 8415
rect 4893 8375 4951 8381
rect 5077 8415 5135 8421
rect 5077 8381 5089 8415
rect 5123 8412 5135 8415
rect 5276 8412 5304 8520
rect 5537 8517 5549 8551
rect 5583 8548 5595 8551
rect 5718 8548 5724 8560
rect 5583 8520 5724 8548
rect 5583 8517 5595 8520
rect 5537 8511 5595 8517
rect 5718 8508 5724 8520
rect 5776 8548 5782 8560
rect 7374 8548 7380 8560
rect 5776 8520 7380 8548
rect 5776 8508 5782 8520
rect 7374 8508 7380 8520
rect 7432 8508 7438 8560
rect 5350 8440 5356 8492
rect 5408 8480 5414 8492
rect 5408 8452 5453 8480
rect 5408 8440 5414 8452
rect 6454 8440 6460 8492
rect 6512 8480 6518 8492
rect 6641 8483 6699 8489
rect 6641 8480 6653 8483
rect 6512 8452 6653 8480
rect 6512 8440 6518 8452
rect 6641 8449 6653 8452
rect 6687 8449 6699 8483
rect 6641 8443 6699 8449
rect 7006 8440 7012 8492
rect 7064 8480 7070 8492
rect 7285 8483 7343 8489
rect 7285 8480 7297 8483
rect 7064 8452 7297 8480
rect 7064 8440 7070 8452
rect 7285 8449 7297 8452
rect 7331 8480 7343 8483
rect 7484 8480 7512 8588
rect 7561 8551 7619 8557
rect 7561 8517 7573 8551
rect 7607 8548 7619 8551
rect 7650 8548 7656 8560
rect 7607 8520 7656 8548
rect 7607 8517 7619 8520
rect 7561 8511 7619 8517
rect 7650 8508 7656 8520
rect 7708 8548 7714 8560
rect 8864 8548 8892 8588
rect 9306 8576 9312 8628
rect 9364 8616 9370 8628
rect 10689 8619 10747 8625
rect 10689 8616 10701 8619
rect 9364 8588 10701 8616
rect 9364 8576 9370 8588
rect 10689 8585 10701 8588
rect 10735 8585 10747 8619
rect 10689 8579 10747 8585
rect 11057 8619 11115 8625
rect 11057 8585 11069 8619
rect 11103 8616 11115 8619
rect 11238 8616 11244 8628
rect 11103 8588 11244 8616
rect 11103 8585 11115 8588
rect 11057 8579 11115 8585
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 12250 8576 12256 8628
rect 12308 8616 12314 8628
rect 12437 8619 12495 8625
rect 12437 8616 12449 8619
rect 12308 8588 12449 8616
rect 12308 8576 12314 8588
rect 12437 8585 12449 8588
rect 12483 8616 12495 8619
rect 13722 8616 13728 8628
rect 12483 8588 13728 8616
rect 12483 8585 12495 8588
rect 12437 8579 12495 8585
rect 13722 8576 13728 8588
rect 13780 8616 13786 8628
rect 14277 8619 14335 8625
rect 13780 8588 14044 8616
rect 13780 8576 13786 8588
rect 9582 8548 9588 8560
rect 7708 8520 8800 8548
rect 8864 8520 9588 8548
rect 7708 8508 7714 8520
rect 8772 8489 8800 8520
rect 9582 8508 9588 8520
rect 9640 8508 9646 8560
rect 9769 8551 9827 8557
rect 9769 8517 9781 8551
rect 9815 8548 9827 8551
rect 10137 8551 10195 8557
rect 10137 8548 10149 8551
rect 9815 8520 10149 8548
rect 9815 8517 9827 8520
rect 9769 8511 9827 8517
rect 10137 8517 10149 8520
rect 10183 8517 10195 8551
rect 10410 8548 10416 8560
rect 10371 8520 10416 8548
rect 10137 8511 10195 8517
rect 10410 8508 10416 8520
rect 10468 8508 10474 8560
rect 11149 8551 11207 8557
rect 11149 8517 11161 8551
rect 11195 8548 11207 8551
rect 11606 8548 11612 8560
rect 11195 8520 11612 8548
rect 11195 8517 11207 8520
rect 11149 8511 11207 8517
rect 11606 8508 11612 8520
rect 11664 8508 11670 8560
rect 12805 8551 12863 8557
rect 12805 8517 12817 8551
rect 12851 8548 12863 8551
rect 12894 8548 12900 8560
rect 12851 8520 12900 8548
rect 12851 8517 12863 8520
rect 12805 8511 12863 8517
rect 12894 8508 12900 8520
rect 12952 8508 12958 8560
rect 14016 8548 14044 8588
rect 14277 8585 14289 8619
rect 14323 8616 14335 8619
rect 16114 8616 16120 8628
rect 14323 8588 16120 8616
rect 14323 8585 14335 8588
rect 14277 8579 14335 8585
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 16758 8548 16764 8560
rect 14016 8534 14780 8548
rect 14030 8520 14780 8534
rect 16238 8520 16764 8548
rect 7331 8452 7512 8480
rect 8205 8483 8263 8489
rect 7331 8449 7343 8452
rect 7285 8443 7343 8449
rect 8205 8449 8217 8483
rect 8251 8480 8263 8483
rect 8665 8483 8723 8489
rect 8665 8480 8677 8483
rect 8251 8452 8677 8480
rect 8251 8449 8263 8452
rect 8205 8443 8263 8449
rect 8665 8449 8677 8452
rect 8711 8449 8723 8483
rect 8665 8443 8723 8449
rect 8757 8483 8815 8489
rect 8757 8449 8769 8483
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 5810 8412 5816 8424
rect 5123 8384 5816 8412
rect 5123 8381 5135 8384
rect 5077 8375 5135 8381
rect 4065 8347 4123 8353
rect 4065 8344 4077 8347
rect 3712 8316 4077 8344
rect 4065 8313 4077 8316
rect 4111 8344 4123 8347
rect 4706 8344 4712 8356
rect 4111 8316 4712 8344
rect 4111 8313 4123 8316
rect 4065 8307 4123 8313
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 4908 8344 4936 8375
rect 5810 8372 5816 8384
rect 5868 8372 5874 8424
rect 6733 8415 6791 8421
rect 6733 8381 6745 8415
rect 6779 8412 6791 8415
rect 7190 8412 7196 8424
rect 6779 8384 7196 8412
rect 6779 8381 6791 8384
rect 6733 8375 6791 8381
rect 7190 8372 7196 8384
rect 7248 8372 7254 8424
rect 7742 8372 7748 8424
rect 7800 8412 7806 8424
rect 8297 8415 8355 8421
rect 8297 8412 8309 8415
rect 7800 8384 8309 8412
rect 7800 8372 7806 8384
rect 8297 8381 8309 8384
rect 8343 8381 8355 8415
rect 8297 8375 8355 8381
rect 8481 8415 8539 8421
rect 8481 8381 8493 8415
rect 8527 8381 8539 8415
rect 8772 8412 8800 8443
rect 8846 8440 8852 8492
rect 8904 8480 8910 8492
rect 9677 8483 9735 8489
rect 9677 8480 9689 8483
rect 8904 8452 9689 8480
rect 8904 8440 8910 8452
rect 9677 8449 9689 8452
rect 9723 8449 9735 8483
rect 9950 8480 9956 8492
rect 9863 8452 9956 8480
rect 9677 8443 9735 8449
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 10226 8480 10232 8492
rect 10187 8452 10232 8480
rect 10226 8440 10232 8452
rect 10284 8440 10290 8492
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8449 10379 8483
rect 12526 8480 12532 8492
rect 12487 8452 12532 8480
rect 10321 8443 10379 8449
rect 9968 8412 9996 8440
rect 8772 8384 9996 8412
rect 8481 8375 8539 8381
rect 7760 8344 7788 8372
rect 4908 8316 7788 8344
rect 8496 8344 8524 8375
rect 8938 8344 8944 8356
rect 8496 8316 8944 8344
rect 8938 8304 8944 8316
rect 8996 8304 9002 8356
rect 9861 8347 9919 8353
rect 9861 8313 9873 8347
rect 9907 8344 9919 8347
rect 10042 8344 10048 8356
rect 9907 8316 10048 8344
rect 9907 8313 9919 8316
rect 9861 8307 9919 8313
rect 10042 8304 10048 8316
rect 10100 8344 10106 8356
rect 10336 8344 10364 8443
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 14366 8440 14372 8492
rect 14424 8480 14430 8492
rect 14461 8483 14519 8489
rect 14461 8480 14473 8483
rect 14424 8452 14473 8480
rect 14424 8440 14430 8452
rect 14461 8449 14473 8452
rect 14507 8449 14519 8483
rect 14461 8443 14519 8449
rect 14550 8440 14556 8492
rect 14608 8480 14614 8492
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 14608 8452 14657 8480
rect 14608 8440 14614 8452
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 14752 8480 14780 8520
rect 16758 8508 16764 8520
rect 16816 8508 16822 8560
rect 15286 8480 15292 8492
rect 14752 8452 15292 8480
rect 14645 8443 14703 8449
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 18233 8483 18291 8489
rect 18233 8449 18245 8483
rect 18279 8480 18291 8483
rect 18509 8483 18567 8489
rect 18509 8480 18521 8483
rect 18279 8452 18521 8480
rect 18279 8449 18291 8452
rect 18233 8443 18291 8449
rect 18509 8449 18521 8452
rect 18555 8480 18567 8483
rect 18598 8480 18604 8492
rect 18555 8452 18604 8480
rect 18555 8449 18567 8452
rect 18509 8443 18567 8449
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 11241 8415 11299 8421
rect 11241 8381 11253 8415
rect 11287 8381 11299 8415
rect 12544 8412 12572 8440
rect 13814 8412 13820 8424
rect 12544 8384 13820 8412
rect 11241 8375 11299 8381
rect 10100 8316 10364 8344
rect 10100 8304 10106 8316
rect 10686 8304 10692 8356
rect 10744 8344 10750 8356
rect 11256 8344 11284 8375
rect 13814 8372 13820 8384
rect 13872 8412 13878 8424
rect 14829 8415 14887 8421
rect 14829 8412 14841 8415
rect 13872 8384 14841 8412
rect 13872 8372 13878 8384
rect 14829 8381 14841 8384
rect 14875 8412 14887 8415
rect 15102 8412 15108 8424
rect 14875 8384 15108 8412
rect 14875 8381 14887 8384
rect 14829 8375 14887 8381
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 15197 8415 15255 8421
rect 15197 8381 15209 8415
rect 15243 8412 15255 8415
rect 15243 8384 18368 8412
rect 15243 8381 15255 8384
rect 15197 8375 15255 8381
rect 14642 8344 14648 8356
rect 10744 8316 11284 8344
rect 14603 8316 14648 8344
rect 10744 8304 10750 8316
rect 14642 8304 14648 8316
rect 14700 8304 14706 8356
rect 18340 8353 18368 8384
rect 18325 8347 18383 8353
rect 18325 8313 18337 8347
rect 18371 8313 18383 8347
rect 18325 8307 18383 8313
rect 2317 8279 2375 8285
rect 2317 8276 2329 8279
rect 1688 8248 2329 8276
rect 2317 8245 2329 8248
rect 2363 8276 2375 8279
rect 2590 8276 2596 8288
rect 2363 8248 2596 8276
rect 2363 8245 2375 8248
rect 2317 8239 2375 8245
rect 2590 8236 2596 8248
rect 2648 8236 2654 8288
rect 2958 8276 2964 8288
rect 2919 8248 2964 8276
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 7650 8236 7656 8288
rect 7708 8276 7714 8288
rect 7837 8279 7895 8285
rect 7837 8276 7849 8279
rect 7708 8248 7849 8276
rect 7708 8236 7714 8248
rect 7837 8245 7849 8248
rect 7883 8245 7895 8279
rect 7837 8239 7895 8245
rect 9950 8236 9956 8288
rect 10008 8276 10014 8288
rect 10778 8276 10784 8288
rect 10008 8248 10784 8276
rect 10008 8236 10014 8248
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 16574 8236 16580 8288
rect 16632 8285 16638 8288
rect 16632 8279 16681 8285
rect 16632 8245 16635 8279
rect 16669 8245 16681 8279
rect 16632 8239 16681 8245
rect 16632 8236 16638 8239
rect 0 8186 18860 8208
rect 0 8134 3110 8186
rect 3162 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 3302 8186
rect 3354 8134 3366 8186
rect 3418 8134 6210 8186
rect 6262 8134 6274 8186
rect 6326 8134 6338 8186
rect 6390 8134 6402 8186
rect 6454 8134 6466 8186
rect 6518 8134 9310 8186
rect 9362 8134 9374 8186
rect 9426 8134 9438 8186
rect 9490 8134 9502 8186
rect 9554 8134 9566 8186
rect 9618 8134 12410 8186
rect 12462 8134 12474 8186
rect 12526 8134 12538 8186
rect 12590 8134 12602 8186
rect 12654 8134 12666 8186
rect 12718 8134 15510 8186
rect 15562 8134 15574 8186
rect 15626 8134 15638 8186
rect 15690 8134 15702 8186
rect 15754 8134 15766 8186
rect 15818 8134 18860 8186
rect 0 8112 18860 8134
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 12802 8072 12808 8084
rect 4304 8044 12808 8072
rect 4304 8032 4310 8044
rect 12802 8032 12808 8044
rect 12860 8032 12866 8084
rect 14918 8032 14924 8084
rect 14976 8072 14982 8084
rect 15105 8075 15163 8081
rect 15105 8072 15117 8075
rect 14976 8044 15117 8072
rect 14976 8032 14982 8044
rect 15105 8041 15117 8044
rect 15151 8041 15163 8075
rect 15105 8035 15163 8041
rect 2774 8013 2780 8016
rect 1949 8007 2007 8013
rect 1949 7973 1961 8007
rect 1995 8004 2007 8007
rect 2731 8007 2780 8013
rect 2731 8004 2743 8007
rect 1995 7976 2743 8004
rect 1995 7973 2007 7976
rect 1949 7967 2007 7973
rect 2731 7973 2743 7976
rect 2777 7973 2780 8007
rect 2731 7967 2780 7973
rect 2774 7964 2780 7967
rect 2832 7964 2838 8016
rect 5350 8004 5356 8016
rect 4356 7976 5356 8004
rect 1765 7939 1823 7945
rect 1765 7905 1777 7939
rect 1811 7936 1823 7939
rect 2317 7939 2375 7945
rect 2317 7936 2329 7939
rect 1811 7908 2329 7936
rect 1811 7905 1823 7908
rect 1765 7899 1823 7905
rect 2317 7905 2329 7908
rect 2363 7905 2375 7939
rect 2317 7899 2375 7905
rect 2501 7939 2559 7945
rect 2501 7905 2513 7939
rect 2547 7936 2559 7939
rect 2958 7936 2964 7948
rect 2547 7908 2964 7936
rect 2547 7905 2559 7908
rect 2501 7899 2559 7905
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7837 2099 7871
rect 2041 7831 2099 7837
rect 2225 7871 2283 7877
rect 2225 7837 2237 7871
rect 2271 7837 2283 7871
rect 2406 7868 2412 7880
rect 2367 7840 2412 7868
rect 2225 7831 2283 7837
rect 566 7692 572 7744
rect 624 7732 630 7744
rect 1765 7735 1823 7741
rect 1765 7732 1777 7735
rect 624 7704 1777 7732
rect 624 7692 630 7704
rect 1765 7701 1777 7704
rect 1811 7701 1823 7735
rect 2056 7732 2084 7831
rect 2240 7800 2268 7831
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2516 7800 2544 7899
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 4062 7896 4068 7948
rect 4120 7936 4126 7948
rect 4356 7945 4384 7976
rect 5350 7964 5356 7976
rect 5408 7964 5414 8016
rect 7190 7964 7196 8016
rect 7248 8004 7254 8016
rect 7285 8007 7343 8013
rect 7285 8004 7297 8007
rect 7248 7976 7297 8004
rect 7248 7964 7254 7976
rect 7285 7973 7297 7976
rect 7331 7973 7343 8007
rect 9950 8004 9956 8016
rect 7285 7967 7343 7973
rect 9600 7976 9956 8004
rect 4341 7939 4399 7945
rect 4341 7936 4353 7939
rect 4120 7908 4353 7936
rect 4120 7896 4126 7908
rect 4341 7905 4353 7908
rect 4387 7905 4399 7939
rect 4341 7899 4399 7905
rect 4816 7908 5580 7936
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 4525 7871 4583 7877
rect 4525 7868 4537 7871
rect 4212 7840 4537 7868
rect 4212 7828 4218 7840
rect 4525 7837 4537 7840
rect 4571 7837 4583 7871
rect 4706 7868 4712 7880
rect 4667 7840 4712 7868
rect 4525 7831 4583 7837
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 4065 7803 4123 7809
rect 4065 7800 4077 7803
rect 2240 7772 2544 7800
rect 2608 7772 4077 7800
rect 2222 7732 2228 7744
rect 2056 7704 2228 7732
rect 1765 7695 1823 7701
rect 2222 7692 2228 7704
rect 2280 7732 2286 7744
rect 2608 7732 2636 7772
rect 4065 7769 4077 7772
rect 4111 7769 4123 7803
rect 4065 7763 4123 7769
rect 2280 7704 2636 7732
rect 2280 7692 2286 7704
rect 3050 7692 3056 7744
rect 3108 7732 3114 7744
rect 3697 7735 3755 7741
rect 3697 7732 3709 7735
rect 3108 7704 3709 7732
rect 3108 7692 3114 7704
rect 3697 7701 3709 7704
rect 3743 7701 3755 7735
rect 3697 7695 3755 7701
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 4816 7741 4844 7908
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 5000 7800 5028 7831
rect 5074 7828 5080 7880
rect 5132 7868 5138 7880
rect 5552 7877 5580 7908
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 7929 7939 7987 7945
rect 7929 7936 7941 7939
rect 6972 7908 7941 7936
rect 6972 7896 6978 7908
rect 7929 7905 7941 7908
rect 7975 7936 7987 7939
rect 8110 7936 8116 7948
rect 7975 7908 8116 7936
rect 7975 7905 7987 7908
rect 7929 7899 7987 7905
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 8386 7896 8392 7948
rect 8444 7936 8450 7948
rect 8444 7908 9536 7936
rect 8444 7896 8450 7908
rect 5445 7871 5503 7877
rect 5445 7868 5457 7871
rect 5132 7840 5177 7868
rect 5276 7840 5457 7868
rect 5132 7828 5138 7840
rect 5169 7803 5227 7809
rect 5169 7800 5181 7803
rect 5000 7772 5181 7800
rect 5169 7769 5181 7772
rect 5215 7769 5227 7803
rect 5169 7763 5227 7769
rect 4157 7735 4215 7741
rect 4157 7732 4169 7735
rect 4028 7704 4169 7732
rect 4028 7692 4034 7704
rect 4157 7701 4169 7704
rect 4203 7701 4215 7735
rect 4157 7695 4215 7701
rect 4801 7735 4859 7741
rect 4801 7701 4813 7735
rect 4847 7701 4859 7735
rect 4801 7695 4859 7701
rect 5074 7692 5080 7744
rect 5132 7732 5138 7744
rect 5184 7732 5212 7763
rect 5276 7741 5304 7840
rect 5445 7837 5457 7840
rect 5491 7837 5503 7871
rect 5445 7831 5503 7837
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7837 5595 7871
rect 5718 7868 5724 7880
rect 5679 7840 5724 7868
rect 5537 7831 5595 7837
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 6086 7828 6092 7880
rect 6144 7868 6150 7880
rect 6273 7871 6331 7877
rect 6273 7868 6285 7871
rect 6144 7840 6285 7868
rect 6144 7828 6150 7840
rect 6273 7837 6285 7840
rect 6319 7837 6331 7871
rect 7650 7868 7656 7880
rect 7611 7840 7656 7868
rect 6273 7831 6331 7837
rect 5350 7760 5356 7812
rect 5408 7800 5414 7812
rect 6288 7800 6316 7831
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 9508 7877 9536 7908
rect 9600 7877 9628 7976
rect 9950 7964 9956 7976
rect 10008 7964 10014 8016
rect 10045 8007 10103 8013
rect 10045 7973 10057 8007
rect 10091 8004 10103 8007
rect 10091 7976 10732 8004
rect 10091 7973 10103 7976
rect 10045 7967 10103 7973
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7837 9551 7871
rect 9493 7831 9551 7837
rect 9585 7871 9643 7877
rect 9585 7837 9597 7871
rect 9631 7837 9643 7871
rect 9858 7868 9864 7880
rect 9819 7840 9864 7868
rect 9585 7831 9643 7837
rect 6822 7800 6828 7812
rect 5408 7772 5453 7800
rect 6288 7772 6828 7800
rect 5408 7760 5414 7772
rect 6822 7760 6828 7772
rect 6880 7760 6886 7812
rect 7009 7803 7067 7809
rect 7009 7769 7021 7803
rect 7055 7800 7067 7803
rect 9122 7800 9128 7812
rect 7055 7772 9128 7800
rect 7055 7769 7067 7772
rect 7009 7763 7067 7769
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 9416 7800 9444 7831
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 10042 7868 10048 7880
rect 10003 7840 10048 7868
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10318 7868 10324 7880
rect 10279 7840 10324 7868
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 9769 7803 9827 7809
rect 9416 7772 9536 7800
rect 5132 7704 5212 7732
rect 5261 7735 5319 7741
rect 5132 7692 5138 7704
rect 5261 7701 5273 7735
rect 5307 7701 5319 7735
rect 5626 7732 5632 7744
rect 5587 7704 5632 7732
rect 5261 7695 5319 7701
rect 5626 7692 5632 7704
rect 5684 7692 5690 7744
rect 6178 7732 6184 7744
rect 6139 7704 6184 7732
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 7650 7692 7656 7744
rect 7708 7732 7714 7744
rect 7745 7735 7803 7741
rect 7745 7732 7757 7735
rect 7708 7704 7757 7732
rect 7708 7692 7714 7704
rect 7745 7701 7757 7704
rect 7791 7701 7803 7735
rect 9508 7732 9536 7772
rect 9769 7769 9781 7803
rect 9815 7800 9827 7803
rect 10428 7800 10456 7831
rect 10502 7828 10508 7880
rect 10560 7868 10566 7880
rect 10704 7877 10732 7976
rect 10778 7964 10784 8016
rect 10836 8004 10842 8016
rect 13633 8007 13691 8013
rect 10836 7976 12434 8004
rect 10836 7964 10842 7976
rect 12406 7936 12434 7976
rect 13633 7973 13645 8007
rect 13679 8004 13691 8007
rect 13814 8004 13820 8016
rect 13679 7976 13820 8004
rect 13679 7973 13691 7976
rect 13633 7967 13691 7973
rect 13814 7964 13820 7976
rect 13872 7964 13878 8016
rect 13265 7939 13323 7945
rect 13265 7936 13277 7939
rect 12406 7908 13277 7936
rect 13265 7905 13277 7908
rect 13311 7905 13323 7939
rect 13265 7899 13323 7905
rect 13722 7896 13728 7948
rect 13780 7936 13786 7948
rect 14001 7939 14059 7945
rect 14001 7936 14013 7939
rect 13780 7908 14013 7936
rect 13780 7896 13786 7908
rect 14001 7905 14013 7908
rect 14047 7905 14059 7939
rect 14458 7936 14464 7948
rect 14419 7908 14464 7936
rect 14001 7899 14059 7905
rect 14458 7896 14464 7908
rect 14516 7896 14522 7948
rect 15102 7896 15108 7948
rect 15160 7936 15166 7948
rect 15749 7939 15807 7945
rect 15749 7936 15761 7939
rect 15160 7908 15761 7936
rect 15160 7896 15166 7908
rect 15749 7905 15761 7908
rect 15795 7905 15807 7939
rect 15749 7899 15807 7905
rect 16117 7939 16175 7945
rect 16117 7905 16129 7939
rect 16163 7936 16175 7939
rect 16574 7936 16580 7948
rect 16163 7908 16580 7936
rect 16163 7905 16175 7908
rect 16117 7899 16175 7905
rect 10689 7871 10747 7877
rect 10560 7840 10605 7868
rect 10560 7828 10566 7840
rect 10689 7837 10701 7871
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 12618 7828 12624 7880
rect 12676 7868 12682 7880
rect 13449 7871 13507 7877
rect 13449 7868 13461 7871
rect 12676 7840 13461 7868
rect 12676 7828 12682 7840
rect 13449 7837 13461 7840
rect 13495 7837 13507 7871
rect 13449 7831 13507 7837
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7837 14151 7871
rect 14734 7868 14740 7880
rect 14695 7840 14740 7868
rect 14093 7831 14151 7837
rect 11330 7800 11336 7812
rect 9815 7772 10456 7800
rect 11291 7772 11336 7800
rect 9815 7769 9827 7772
rect 9769 7763 9827 7769
rect 11330 7760 11336 7772
rect 11388 7760 11394 7812
rect 14108 7800 14136 7831
rect 14734 7828 14740 7840
rect 14792 7828 14798 7880
rect 15764 7868 15792 7899
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 17494 7936 17500 7948
rect 17455 7908 17500 7936
rect 17494 7896 17500 7908
rect 17552 7936 17558 7948
rect 18046 7936 18052 7948
rect 17552 7908 18052 7936
rect 17552 7896 17558 7908
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 15838 7868 15844 7880
rect 15764 7840 15844 7868
rect 15838 7828 15844 7840
rect 15896 7828 15902 7880
rect 14366 7800 14372 7812
rect 14108 7772 14372 7800
rect 14366 7760 14372 7772
rect 14424 7760 14430 7812
rect 10042 7732 10048 7744
rect 9508 7704 10048 7732
rect 7745 7695 7803 7701
rect 10042 7692 10048 7704
rect 10100 7692 10106 7744
rect 10410 7732 10416 7744
rect 10371 7704 10416 7732
rect 10410 7692 10416 7704
rect 10468 7692 10474 7744
rect 10778 7692 10784 7744
rect 10836 7732 10842 7744
rect 11425 7735 11483 7741
rect 11425 7732 11437 7735
rect 10836 7704 11437 7732
rect 10836 7692 10842 7704
rect 11425 7701 11437 7704
rect 11471 7732 11483 7735
rect 12802 7732 12808 7744
rect 11471 7704 12808 7732
rect 11471 7701 11483 7704
rect 11425 7695 11483 7701
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 14645 7735 14703 7741
rect 14645 7701 14657 7735
rect 14691 7732 14703 7735
rect 14918 7732 14924 7744
rect 14691 7704 14924 7732
rect 14691 7701 14703 7704
rect 14645 7695 14703 7701
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 15286 7692 15292 7744
rect 15344 7732 15350 7744
rect 15473 7735 15531 7741
rect 15473 7732 15485 7735
rect 15344 7704 15485 7732
rect 15344 7692 15350 7704
rect 15473 7701 15485 7704
rect 15519 7732 15531 7735
rect 16500 7732 16528 7786
rect 16758 7732 16764 7744
rect 15519 7704 16764 7732
rect 15519 7701 15531 7704
rect 15473 7695 15531 7701
rect 16758 7692 16764 7704
rect 16816 7692 16822 7744
rect 0 7642 18860 7664
rect 0 7590 4660 7642
rect 4712 7590 4724 7642
rect 4776 7590 4788 7642
rect 4840 7590 4852 7642
rect 4904 7590 4916 7642
rect 4968 7590 7760 7642
rect 7812 7590 7824 7642
rect 7876 7590 7888 7642
rect 7940 7590 7952 7642
rect 8004 7590 8016 7642
rect 8068 7590 10860 7642
rect 10912 7590 10924 7642
rect 10976 7590 10988 7642
rect 11040 7590 11052 7642
rect 11104 7590 11116 7642
rect 11168 7590 13960 7642
rect 14012 7590 14024 7642
rect 14076 7590 14088 7642
rect 14140 7590 14152 7642
rect 14204 7590 14216 7642
rect 14268 7590 17060 7642
rect 17112 7590 17124 7642
rect 17176 7590 17188 7642
rect 17240 7590 17252 7642
rect 17304 7590 17316 7642
rect 17368 7590 18860 7642
rect 0 7568 18860 7590
rect 2222 7528 2228 7540
rect 2183 7500 2228 7528
rect 2222 7488 2228 7500
rect 2280 7488 2286 7540
rect 2406 7488 2412 7540
rect 2464 7528 2470 7540
rect 2685 7531 2743 7537
rect 2685 7528 2697 7531
rect 2464 7500 2697 7528
rect 2464 7488 2470 7500
rect 2685 7497 2697 7500
rect 2731 7497 2743 7531
rect 3050 7528 3056 7540
rect 3011 7500 3056 7528
rect 2685 7491 2743 7497
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 3145 7531 3203 7537
rect 3145 7497 3157 7531
rect 3191 7528 3203 7531
rect 3970 7528 3976 7540
rect 3191 7500 3976 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 3970 7488 3976 7500
rect 4028 7488 4034 7540
rect 6178 7528 6184 7540
rect 5184 7500 6184 7528
rect 566 7460 572 7472
rect 527 7432 572 7460
rect 566 7420 572 7432
rect 624 7420 630 7472
rect 2590 7460 2596 7472
rect 1794 7432 2596 7460
rect 2590 7420 2596 7432
rect 2648 7420 2654 7472
rect 2314 7392 2320 7404
rect 2056 7364 2320 7392
rect 2056 7333 2084 7364
rect 2314 7352 2320 7364
rect 2372 7352 2378 7404
rect 5184 7401 5212 7500
rect 6178 7488 6184 7500
rect 6236 7488 6242 7540
rect 9769 7531 9827 7537
rect 9769 7497 9781 7531
rect 9815 7528 9827 7531
rect 9953 7531 10011 7537
rect 9953 7528 9965 7531
rect 9815 7500 9965 7528
rect 9815 7497 9827 7500
rect 9769 7491 9827 7497
rect 9953 7497 9965 7500
rect 9999 7528 10011 7531
rect 12618 7528 12624 7540
rect 9999 7500 11468 7528
rect 12579 7500 12624 7528
rect 9999 7497 10011 7500
rect 9953 7491 10011 7497
rect 11440 7472 11468 7500
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 13170 7488 13176 7540
rect 13228 7528 13234 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 13228 7500 13461 7528
rect 13228 7488 13234 7500
rect 13449 7497 13461 7500
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 5902 7420 5908 7472
rect 5960 7420 5966 7472
rect 7484 7432 10180 7460
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7361 5227 7395
rect 5169 7355 5227 7361
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7392 5595 7395
rect 5626 7392 5632 7404
rect 5583 7364 5632 7392
rect 5583 7361 5595 7364
rect 5537 7355 5595 7361
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 7484 7401 7512 7432
rect 6963 7395 7021 7401
rect 6963 7361 6975 7395
rect 7009 7392 7021 7395
rect 7469 7395 7527 7401
rect 7469 7392 7481 7395
rect 7009 7364 7481 7392
rect 7009 7361 7021 7364
rect 6963 7355 7021 7361
rect 7469 7361 7481 7364
rect 7515 7361 7527 7395
rect 8754 7392 8760 7404
rect 8715 7364 8760 7392
rect 7469 7355 7527 7361
rect 8754 7352 8760 7364
rect 8812 7352 8818 7404
rect 293 7327 351 7333
rect 293 7293 305 7327
rect 339 7293 351 7327
rect 293 7287 351 7293
rect 2041 7327 2099 7333
rect 2041 7293 2053 7327
rect 2087 7293 2099 7327
rect 2041 7287 2099 7293
rect 3329 7327 3387 7333
rect 3329 7293 3341 7327
rect 3375 7324 3387 7327
rect 3786 7324 3792 7336
rect 3375 7296 3792 7324
rect 3375 7293 3387 7296
rect 3329 7287 3387 7293
rect 308 7188 336 7287
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 5074 7284 5080 7336
rect 5132 7324 5138 7336
rect 7377 7327 7435 7333
rect 7377 7324 7389 7327
rect 5132 7296 7389 7324
rect 5132 7284 5138 7296
rect 7377 7293 7389 7296
rect 7423 7293 7435 7327
rect 7377 7287 7435 7293
rect 8481 7327 8539 7333
rect 8481 7293 8493 7327
rect 8527 7324 8539 7327
rect 8846 7324 8852 7336
rect 8527 7296 8852 7324
rect 8527 7293 8539 7296
rect 8481 7287 8539 7293
rect 8846 7284 8852 7296
rect 8904 7284 8910 7336
rect 9674 7284 9680 7336
rect 9732 7324 9738 7336
rect 10045 7327 10103 7333
rect 10045 7324 10057 7327
rect 9732 7296 10057 7324
rect 9732 7284 9738 7296
rect 10045 7293 10057 7296
rect 10091 7293 10103 7327
rect 10152 7324 10180 7432
rect 11422 7420 11428 7472
rect 11480 7420 11486 7472
rect 13557 7469 13563 7472
rect 13541 7463 13563 7469
rect 13541 7429 13553 7463
rect 13541 7423 13563 7429
rect 13557 7420 13563 7423
rect 13615 7420 13621 7472
rect 14185 7463 14243 7469
rect 14185 7429 14197 7463
rect 14231 7460 14243 7463
rect 14550 7460 14556 7472
rect 14231 7432 14556 7460
rect 14231 7429 14243 7432
rect 14185 7423 14243 7429
rect 14550 7420 14556 7432
rect 14608 7420 14614 7472
rect 16758 7460 16764 7472
rect 15870 7432 16764 7460
rect 16758 7420 16764 7432
rect 16816 7420 16822 7472
rect 10410 7392 10416 7404
rect 10371 7364 10416 7392
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 11882 7401 11888 7404
rect 11839 7395 11888 7401
rect 11839 7392 11851 7395
rect 11795 7364 11851 7392
rect 11839 7361 11851 7364
rect 11885 7361 11888 7395
rect 11839 7355 11888 7361
rect 11882 7352 11888 7355
rect 11940 7392 11946 7404
rect 12253 7395 12311 7401
rect 12253 7392 12265 7395
rect 11940 7364 12265 7392
rect 11940 7352 11946 7364
rect 12253 7361 12265 7364
rect 12299 7361 12311 7395
rect 12894 7392 12900 7404
rect 12855 7364 12900 7392
rect 12253 7355 12311 7361
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 13170 7392 13176 7404
rect 13131 7364 13176 7392
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 13354 7392 13360 7404
rect 13315 7364 13360 7392
rect 13354 7352 13360 7364
rect 13412 7352 13418 7404
rect 13446 7352 13452 7404
rect 13504 7392 13510 7404
rect 13722 7395 13780 7401
rect 13504 7364 13549 7392
rect 13504 7352 13510 7364
rect 13722 7361 13734 7395
rect 13768 7390 13780 7395
rect 13998 7392 14004 7404
rect 13826 7390 14004 7392
rect 13768 7364 14004 7390
rect 13768 7362 13854 7364
rect 13768 7361 13780 7362
rect 13722 7355 13780 7361
rect 13998 7352 14004 7364
rect 14056 7352 14062 7404
rect 14274 7392 14280 7404
rect 14235 7364 14280 7392
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 16850 7352 16856 7404
rect 16908 7392 16914 7404
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 16908 7364 17049 7392
rect 16908 7352 16914 7364
rect 17037 7361 17049 7364
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 12161 7327 12219 7333
rect 12161 7324 12173 7327
rect 10152 7296 12173 7324
rect 10045 7287 10103 7293
rect 12161 7293 12173 7296
rect 12207 7293 12219 7327
rect 12161 7287 12219 7293
rect 8941 7259 8999 7265
rect 8941 7225 8953 7259
rect 8987 7256 8999 7259
rect 9950 7256 9956 7268
rect 8987 7228 9956 7256
rect 8987 7225 8999 7228
rect 8941 7219 8999 7225
rect 9950 7216 9956 7228
rect 10008 7216 10014 7268
rect 750 7188 756 7200
rect 308 7160 756 7188
rect 750 7148 756 7160
rect 808 7148 814 7200
rect 2590 7188 2596 7200
rect 2551 7160 2596 7188
rect 2590 7148 2596 7160
rect 2648 7148 2654 7200
rect 5077 7191 5135 7197
rect 5077 7157 5089 7191
rect 5123 7188 5135 7191
rect 5350 7188 5356 7200
rect 5123 7160 5356 7188
rect 5123 7157 5135 7160
rect 5077 7151 5135 7157
rect 5350 7148 5356 7160
rect 5408 7188 5414 7200
rect 5902 7188 5908 7200
rect 5408 7160 5908 7188
rect 5408 7148 5414 7160
rect 5902 7148 5908 7160
rect 5960 7148 5966 7200
rect 8570 7188 8576 7200
rect 8531 7160 8576 7188
rect 8570 7148 8576 7160
rect 8628 7148 8634 7200
rect 10060 7188 10088 7287
rect 12802 7284 12808 7336
rect 12860 7324 12866 7336
rect 14458 7324 14464 7336
rect 12860 7296 14464 7324
rect 12860 7284 12866 7296
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 14734 7284 14740 7336
rect 14792 7324 14798 7336
rect 14829 7327 14887 7333
rect 14829 7324 14841 7327
rect 14792 7296 14841 7324
rect 14792 7284 14798 7296
rect 14829 7293 14841 7296
rect 14875 7293 14887 7327
rect 14829 7287 14887 7293
rect 13262 7256 13268 7268
rect 13223 7228 13268 7256
rect 13262 7216 13268 7228
rect 13320 7216 13326 7268
rect 13630 7216 13636 7268
rect 13688 7256 13694 7268
rect 13817 7259 13875 7265
rect 13817 7256 13829 7259
rect 13688 7228 13829 7256
rect 13688 7216 13694 7228
rect 13817 7225 13829 7228
rect 13863 7225 13875 7259
rect 13817 7219 13875 7225
rect 10778 7188 10784 7200
rect 10060 7160 10784 7188
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 11146 7148 11152 7200
rect 11204 7188 11210 7200
rect 11330 7188 11336 7200
rect 11204 7160 11336 7188
rect 11204 7148 11210 7160
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 12989 7191 13047 7197
rect 12989 7157 13001 7191
rect 13035 7188 13047 7191
rect 13722 7188 13728 7200
rect 13035 7160 13728 7188
rect 13035 7157 13047 7160
rect 12989 7151 13047 7157
rect 13722 7148 13728 7160
rect 13780 7188 13786 7200
rect 14274 7188 14280 7200
rect 13780 7160 14280 7188
rect 13780 7148 13786 7160
rect 14274 7148 14280 7160
rect 14332 7148 14338 7200
rect 15286 7148 15292 7200
rect 15344 7188 15350 7200
rect 16255 7191 16313 7197
rect 16255 7188 16267 7191
rect 15344 7160 16267 7188
rect 15344 7148 15350 7160
rect 16255 7157 16267 7160
rect 16301 7157 16313 7191
rect 16255 7151 16313 7157
rect 16574 7148 16580 7200
rect 16632 7188 16638 7200
rect 16853 7191 16911 7197
rect 16853 7188 16865 7191
rect 16632 7160 16865 7188
rect 16632 7148 16638 7160
rect 16853 7157 16865 7160
rect 16899 7157 16911 7191
rect 16853 7151 16911 7157
rect 0 7098 18860 7120
rect 0 7046 3110 7098
rect 3162 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 3302 7098
rect 3354 7046 3366 7098
rect 3418 7046 6210 7098
rect 6262 7046 6274 7098
rect 6326 7046 6338 7098
rect 6390 7046 6402 7098
rect 6454 7046 6466 7098
rect 6518 7046 9310 7098
rect 9362 7046 9374 7098
rect 9426 7046 9438 7098
rect 9490 7046 9502 7098
rect 9554 7046 9566 7098
rect 9618 7046 12410 7098
rect 12462 7046 12474 7098
rect 12526 7046 12538 7098
rect 12590 7046 12602 7098
rect 12654 7046 12666 7098
rect 12718 7046 15510 7098
rect 15562 7046 15574 7098
rect 15626 7046 15638 7098
rect 15690 7046 15702 7098
rect 15754 7046 15766 7098
rect 15818 7046 18860 7098
rect 0 7024 18860 7046
rect 2133 6987 2191 6993
rect 2133 6953 2145 6987
rect 2179 6984 2191 6987
rect 2774 6984 2780 6996
rect 2179 6956 2780 6984
rect 2179 6953 2191 6956
rect 2133 6947 2191 6953
rect 2774 6944 2780 6956
rect 2832 6984 2838 6996
rect 2958 6984 2964 6996
rect 2832 6956 2964 6984
rect 2832 6944 2838 6956
rect 2958 6944 2964 6956
rect 3016 6944 3022 6996
rect 10318 6944 10324 6996
rect 10376 6984 10382 6996
rect 11609 6987 11667 6993
rect 11609 6984 11621 6987
rect 10376 6956 11621 6984
rect 10376 6944 10382 6956
rect 11609 6953 11621 6956
rect 11655 6953 11667 6987
rect 14366 6984 14372 6996
rect 14327 6956 14372 6984
rect 11609 6947 11667 6953
rect 14366 6944 14372 6956
rect 14424 6944 14430 6996
rect 16104 6987 16162 6993
rect 16104 6953 16116 6987
rect 16150 6984 16162 6987
rect 16666 6984 16672 6996
rect 16150 6956 16672 6984
rect 16150 6953 16162 6956
rect 16104 6947 16162 6953
rect 16666 6944 16672 6956
rect 16724 6944 16730 6996
rect 2593 6919 2651 6925
rect 2593 6885 2605 6919
rect 2639 6916 2651 6919
rect 7929 6919 7987 6925
rect 2639 6888 3188 6916
rect 2639 6885 2651 6888
rect 2593 6879 2651 6885
rect 1949 6851 2007 6857
rect 1949 6817 1961 6851
rect 1995 6848 2007 6851
rect 3053 6851 3111 6857
rect 3053 6848 3065 6851
rect 1995 6820 3065 6848
rect 1995 6817 2007 6820
rect 1949 6811 2007 6817
rect 3053 6817 3065 6820
rect 3099 6817 3111 6851
rect 3160 6848 3188 6888
rect 7929 6885 7941 6919
rect 7975 6885 7987 6919
rect 7929 6879 7987 6885
rect 4154 6848 4160 6860
rect 3160 6820 4160 6848
rect 3053 6811 3111 6817
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6848 4399 6851
rect 5442 6848 5448 6860
rect 4387 6820 5448 6848
rect 4387 6817 4399 6820
rect 4341 6811 4399 6817
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2593 6783 2651 6789
rect 2593 6780 2605 6783
rect 2271 6752 2605 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2593 6749 2605 6752
rect 2639 6780 2651 6783
rect 2777 6783 2835 6789
rect 2777 6780 2789 6783
rect 2639 6752 2789 6780
rect 2639 6749 2651 6752
rect 2593 6743 2651 6749
rect 2777 6749 2789 6752
rect 2823 6749 2835 6783
rect 2777 6743 2835 6749
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 2869 6743 2927 6749
rect 2314 6712 2320 6724
rect 2275 6684 2320 6712
rect 2314 6672 2320 6684
rect 2372 6672 2378 6724
rect 2406 6672 2412 6724
rect 2464 6712 2470 6724
rect 2501 6715 2559 6721
rect 2501 6712 2513 6715
rect 2464 6684 2513 6712
rect 2464 6672 2470 6684
rect 2501 6681 2513 6684
rect 2547 6681 2559 6715
rect 2501 6675 2559 6681
rect 1946 6644 1952 6656
rect 1907 6616 1952 6644
rect 1946 6604 1952 6616
rect 2004 6604 2010 6656
rect 2038 6604 2044 6656
rect 2096 6644 2102 6656
rect 2884 6644 2912 6743
rect 2958 6740 2964 6792
rect 3016 6780 3022 6792
rect 3145 6783 3203 6789
rect 3016 6752 3061 6780
rect 3016 6740 3022 6752
rect 3145 6749 3157 6783
rect 3191 6780 3203 6783
rect 3191 6752 3740 6780
rect 3191 6749 3203 6752
rect 3145 6743 3203 6749
rect 3712 6653 3740 6752
rect 3786 6740 3792 6792
rect 3844 6780 3850 6792
rect 4356 6780 4384 6811
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 7944 6848 7972 6879
rect 11146 6876 11152 6928
rect 11204 6876 11210 6928
rect 11514 6916 11520 6928
rect 11348 6888 11520 6916
rect 9122 6848 9128 6860
rect 7944 6820 8340 6848
rect 9035 6820 9128 6848
rect 3844 6752 4384 6780
rect 6549 6783 6607 6789
rect 3844 6740 3850 6752
rect 6549 6749 6561 6783
rect 6595 6780 6607 6783
rect 8113 6783 8171 6789
rect 6595 6752 8064 6780
rect 6595 6749 6607 6752
rect 6549 6743 6607 6749
rect 6730 6672 6736 6724
rect 6788 6721 6794 6724
rect 6788 6715 6852 6721
rect 6788 6681 6806 6715
rect 6840 6681 6852 6715
rect 8036 6712 8064 6752
rect 8113 6749 8125 6783
rect 8159 6780 8171 6783
rect 8202 6780 8208 6792
rect 8159 6752 8208 6780
rect 8159 6749 8171 6752
rect 8113 6743 8171 6749
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 8312 6789 8340 6820
rect 9122 6808 9128 6820
rect 9180 6848 9186 6860
rect 11164 6848 11192 6876
rect 11348 6857 11376 6888
rect 11514 6876 11520 6888
rect 11572 6876 11578 6928
rect 13998 6876 14004 6928
rect 14056 6916 14062 6928
rect 15289 6919 15347 6925
rect 15289 6916 15301 6919
rect 14056 6888 15301 6916
rect 14056 6876 14062 6888
rect 15289 6885 15301 6888
rect 15335 6885 15347 6919
rect 15289 6879 15347 6885
rect 9180 6820 11192 6848
rect 11333 6851 11391 6857
rect 9180 6808 9186 6820
rect 11333 6817 11345 6851
rect 11379 6817 11391 6851
rect 11333 6811 11391 6817
rect 13722 6808 13728 6860
rect 13780 6848 13786 6860
rect 14093 6851 14151 6857
rect 14093 6848 14105 6851
rect 13780 6820 14105 6848
rect 13780 6808 13786 6820
rect 14093 6817 14105 6820
rect 14139 6817 14151 6851
rect 14093 6811 14151 6817
rect 14458 6808 14464 6860
rect 14516 6848 14522 6860
rect 14829 6851 14887 6857
rect 14829 6848 14841 6851
rect 14516 6820 14841 6848
rect 14516 6808 14522 6820
rect 14829 6817 14841 6820
rect 14875 6817 14887 6851
rect 14829 6811 14887 6817
rect 14921 6851 14979 6857
rect 14921 6817 14933 6851
rect 14967 6817 14979 6851
rect 18414 6848 18420 6860
rect 14921 6811 14979 6817
rect 15488 6820 18420 6848
rect 8297 6783 8355 6789
rect 8297 6749 8309 6783
rect 8343 6780 8355 6783
rect 9306 6780 9312 6792
rect 8343 6752 9312 6780
rect 8343 6749 8355 6752
rect 8297 6743 8355 6749
rect 9306 6740 9312 6752
rect 9364 6740 9370 6792
rect 10778 6740 10784 6792
rect 10836 6780 10842 6792
rect 11057 6783 11115 6789
rect 11057 6780 11069 6783
rect 10836 6752 11069 6780
rect 10836 6740 10842 6752
rect 11057 6749 11069 6752
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6780 11299 6783
rect 11606 6780 11612 6792
rect 11287 6752 11612 6780
rect 11287 6749 11299 6752
rect 11241 6743 11299 6749
rect 11606 6740 11612 6752
rect 11664 6740 11670 6792
rect 11709 6783 11767 6789
rect 11709 6749 11721 6783
rect 11755 6780 11767 6783
rect 11882 6780 11888 6792
rect 11755 6752 11888 6780
rect 11755 6749 11767 6752
rect 11709 6743 11767 6749
rect 11882 6740 11888 6752
rect 11940 6740 11946 6792
rect 13814 6740 13820 6792
rect 13872 6780 13878 6792
rect 14001 6783 14059 6789
rect 14001 6780 14013 6783
rect 13872 6752 14013 6780
rect 13872 6740 13878 6752
rect 14001 6749 14013 6752
rect 14047 6749 14059 6783
rect 14001 6743 14059 6749
rect 14185 6783 14243 6789
rect 14185 6749 14197 6783
rect 14231 6780 14243 6783
rect 14366 6780 14372 6792
rect 14231 6752 14372 6780
rect 14231 6749 14243 6752
rect 14185 6743 14243 6749
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 14642 6740 14648 6792
rect 14700 6780 14706 6792
rect 14936 6780 14964 6811
rect 14700 6752 14964 6780
rect 14700 6740 14706 6752
rect 15286 6740 15292 6792
rect 15344 6780 15350 6792
rect 15381 6783 15439 6789
rect 15381 6780 15393 6783
rect 15344 6752 15393 6780
rect 15344 6740 15350 6752
rect 15381 6749 15393 6752
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 9674 6712 9680 6724
rect 8036 6684 9680 6712
rect 6788 6675 6852 6681
rect 6788 6672 6794 6675
rect 9674 6672 9680 6684
rect 9732 6672 9738 6724
rect 10689 6715 10747 6721
rect 10689 6681 10701 6715
rect 10735 6712 10747 6715
rect 11793 6715 11851 6721
rect 11793 6712 11805 6715
rect 10735 6684 11805 6712
rect 10735 6681 10747 6684
rect 10689 6675 10747 6681
rect 11793 6681 11805 6684
rect 11839 6712 11851 6715
rect 15488 6712 15516 6820
rect 18414 6808 18420 6820
rect 18472 6808 18478 6860
rect 15838 6780 15844 6792
rect 15799 6752 15844 6780
rect 15838 6740 15844 6752
rect 15896 6740 15902 6792
rect 18233 6783 18291 6789
rect 18233 6749 18245 6783
rect 18279 6780 18291 6783
rect 18506 6780 18512 6792
rect 18279 6752 18512 6780
rect 18279 6749 18291 6752
rect 18233 6743 18291 6749
rect 18506 6740 18512 6752
rect 18564 6740 18570 6792
rect 11839 6684 15516 6712
rect 15749 6715 15807 6721
rect 11839 6681 11851 6684
rect 11793 6675 11851 6681
rect 15749 6681 15761 6715
rect 15795 6712 15807 6715
rect 16206 6712 16212 6724
rect 15795 6684 16212 6712
rect 15795 6681 15807 6684
rect 15749 6675 15807 6681
rect 16206 6672 16212 6684
rect 16264 6672 16270 6724
rect 16758 6672 16764 6724
rect 16816 6672 16822 6724
rect 17402 6672 17408 6724
rect 17460 6712 17466 6724
rect 17865 6715 17923 6721
rect 17865 6712 17877 6715
rect 17460 6684 17877 6712
rect 17460 6672 17466 6684
rect 17865 6681 17877 6684
rect 17911 6681 17923 6715
rect 17865 6675 17923 6681
rect 2096 6616 2912 6644
rect 3697 6647 3755 6653
rect 2096 6604 2102 6616
rect 3697 6613 3709 6647
rect 3743 6613 3755 6647
rect 3697 6607 3755 6613
rect 3878 6604 3884 6656
rect 3936 6644 3942 6656
rect 4065 6647 4123 6653
rect 4065 6644 4077 6647
rect 3936 6616 4077 6644
rect 3936 6604 3942 6616
rect 4065 6613 4077 6616
rect 4111 6613 4123 6647
rect 4065 6607 4123 6613
rect 4157 6647 4215 6653
rect 4157 6613 4169 6647
rect 4203 6644 4215 6647
rect 4338 6644 4344 6656
rect 4203 6616 4344 6644
rect 4203 6613 4215 6616
rect 4157 6607 4215 6613
rect 4338 6604 4344 6616
rect 4396 6604 4402 6656
rect 8110 6604 8116 6656
rect 8168 6644 8174 6656
rect 8205 6647 8263 6653
rect 8205 6644 8217 6647
rect 8168 6616 8217 6644
rect 8168 6604 8174 6616
rect 8205 6613 8217 6616
rect 8251 6613 8263 6647
rect 8205 6607 8263 6613
rect 8386 6604 8392 6656
rect 8444 6644 8450 6656
rect 10873 6647 10931 6653
rect 10873 6644 10885 6647
rect 8444 6616 10885 6644
rect 8444 6604 8450 6616
rect 10873 6613 10885 6616
rect 10919 6613 10931 6647
rect 13630 6644 13636 6656
rect 13591 6616 13636 6644
rect 10873 6607 10931 6613
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 13817 6647 13875 6653
rect 13817 6613 13829 6647
rect 13863 6644 13875 6647
rect 14642 6644 14648 6656
rect 13863 6616 14648 6644
rect 13863 6613 13875 6616
rect 13817 6607 13875 6613
rect 14642 6604 14648 6616
rect 14700 6604 14706 6656
rect 14737 6647 14795 6653
rect 14737 6613 14749 6647
rect 14783 6644 14795 6647
rect 15194 6644 15200 6656
rect 14783 6616 15200 6644
rect 14783 6613 14795 6616
rect 14737 6607 14795 6613
rect 15194 6604 15200 6616
rect 15252 6604 15258 6656
rect 15838 6604 15844 6656
rect 15896 6644 15902 6656
rect 18325 6647 18383 6653
rect 18325 6644 18337 6647
rect 15896 6616 18337 6644
rect 15896 6604 15902 6616
rect 18325 6613 18337 6616
rect 18371 6613 18383 6647
rect 18325 6607 18383 6613
rect 0 6554 18860 6576
rect 0 6502 4660 6554
rect 4712 6502 4724 6554
rect 4776 6502 4788 6554
rect 4840 6502 4852 6554
rect 4904 6502 4916 6554
rect 4968 6502 7760 6554
rect 7812 6502 7824 6554
rect 7876 6502 7888 6554
rect 7940 6502 7952 6554
rect 8004 6502 8016 6554
rect 8068 6502 10860 6554
rect 10912 6502 10924 6554
rect 10976 6502 10988 6554
rect 11040 6502 11052 6554
rect 11104 6502 11116 6554
rect 11168 6502 13960 6554
rect 14012 6502 14024 6554
rect 14076 6502 14088 6554
rect 14140 6502 14152 6554
rect 14204 6502 14216 6554
rect 14268 6502 17060 6554
rect 17112 6502 17124 6554
rect 17176 6502 17188 6554
rect 17240 6502 17252 6554
rect 17304 6502 17316 6554
rect 17368 6502 18860 6554
rect 0 6480 18860 6502
rect 750 6400 756 6452
rect 808 6400 814 6452
rect 2958 6440 2964 6452
rect 2148 6412 2964 6440
rect 768 6372 796 6400
rect 1854 6372 1860 6384
rect 308 6344 796 6372
rect 1794 6344 1860 6372
rect 308 6313 336 6344
rect 1854 6332 1860 6344
rect 1912 6332 1918 6384
rect 2148 6313 2176 6412
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 3878 6440 3884 6452
rect 3839 6412 3884 6440
rect 3878 6400 3884 6412
rect 3936 6400 3942 6452
rect 4893 6443 4951 6449
rect 4893 6409 4905 6443
rect 4939 6409 4951 6443
rect 4893 6403 4951 6409
rect 4908 6372 4936 6403
rect 5166 6400 5172 6452
rect 5224 6440 5230 6452
rect 5353 6443 5411 6449
rect 5353 6440 5365 6443
rect 5224 6412 5365 6440
rect 5224 6400 5230 6412
rect 5353 6409 5365 6412
rect 5399 6409 5411 6443
rect 5353 6403 5411 6409
rect 8389 6443 8447 6449
rect 8389 6409 8401 6443
rect 8435 6440 8447 6443
rect 8570 6440 8576 6452
rect 8435 6412 8576 6440
rect 8435 6409 8447 6412
rect 8389 6403 8447 6409
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 11606 6440 11612 6452
rect 9232 6412 11612 6440
rect 5810 6372 5816 6384
rect 2332 6344 4936 6372
rect 5184 6344 5816 6372
rect 2332 6313 2360 6344
rect 293 6307 351 6313
rect 293 6273 305 6307
rect 339 6273 351 6307
rect 293 6267 351 6273
rect 2133 6307 2191 6313
rect 2133 6273 2145 6307
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6273 2375 6307
rect 2317 6267 2375 6273
rect 2406 6264 2412 6316
rect 2464 6304 2470 6316
rect 2777 6307 2835 6313
rect 2777 6304 2789 6307
rect 2464 6276 2789 6304
rect 2464 6264 2470 6276
rect 2777 6273 2789 6276
rect 2823 6273 2835 6307
rect 4246 6304 4252 6316
rect 4207 6276 4252 6304
rect 2777 6267 2835 6273
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 4338 6264 4344 6316
rect 4396 6304 4402 6316
rect 5184 6304 5212 6344
rect 5810 6332 5816 6344
rect 5868 6372 5874 6384
rect 6730 6372 6736 6384
rect 5868 6344 6736 6372
rect 5868 6332 5874 6344
rect 6730 6332 6736 6344
rect 6788 6372 6794 6384
rect 8202 6372 8208 6384
rect 6788 6344 8208 6372
rect 6788 6332 6794 6344
rect 8202 6332 8208 6344
rect 8260 6372 8266 6384
rect 9232 6372 9260 6412
rect 11606 6400 11612 6412
rect 11664 6400 11670 6452
rect 12710 6440 12716 6452
rect 12084 6412 12716 6440
rect 9950 6372 9956 6384
rect 8260 6344 9260 6372
rect 9911 6344 9956 6372
rect 8260 6332 8266 6344
rect 4396 6276 5212 6304
rect 5261 6307 5319 6313
rect 4396 6264 4402 6276
rect 5261 6273 5273 6307
rect 5307 6304 5319 6307
rect 5626 6304 5632 6316
rect 5307 6276 5632 6304
rect 5307 6273 5319 6276
rect 5261 6267 5319 6273
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 8110 6304 8116 6316
rect 8071 6276 8116 6304
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 8478 6304 8484 6316
rect 8439 6276 8484 6304
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 9232 6313 9260 6344
rect 9950 6332 9956 6344
rect 10008 6332 10014 6384
rect 9033 6307 9091 6313
rect 9033 6304 9045 6307
rect 8588 6276 9045 6304
rect 569 6239 627 6245
rect 569 6205 581 6239
rect 615 6236 627 6239
rect 1946 6236 1952 6248
rect 615 6208 1952 6236
rect 615 6205 627 6208
rect 569 6199 627 6205
rect 1946 6196 1952 6208
rect 2004 6196 2010 6248
rect 2225 6239 2283 6245
rect 2225 6205 2237 6239
rect 2271 6236 2283 6239
rect 2501 6239 2559 6245
rect 2501 6236 2513 6239
rect 2271 6208 2513 6236
rect 2271 6205 2283 6208
rect 2225 6199 2283 6205
rect 2501 6205 2513 6208
rect 2547 6205 2559 6239
rect 2501 6199 2559 6205
rect 2685 6239 2743 6245
rect 2685 6205 2697 6239
rect 2731 6236 2743 6239
rect 2958 6236 2964 6248
rect 2731 6208 2964 6236
rect 2731 6205 2743 6208
rect 2685 6199 2743 6205
rect 2958 6196 2964 6208
rect 3016 6196 3022 6248
rect 4433 6239 4491 6245
rect 4433 6205 4445 6239
rect 4479 6205 4491 6239
rect 4433 6199 4491 6205
rect 2593 6171 2651 6177
rect 2593 6168 2605 6171
rect 1596 6140 2605 6168
rect 934 6060 940 6112
rect 992 6100 998 6112
rect 1596 6100 1624 6140
rect 2593 6137 2605 6140
rect 2639 6137 2651 6171
rect 2593 6131 2651 6137
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 4448 6168 4476 6199
rect 5442 6196 5448 6248
rect 5500 6236 5506 6248
rect 6914 6236 6920 6248
rect 5500 6208 6920 6236
rect 5500 6196 5506 6208
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 8386 6236 8392 6248
rect 8347 6208 8392 6236
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 4120 6140 4476 6168
rect 8205 6171 8263 6177
rect 4120 6128 4126 6140
rect 8205 6137 8217 6171
rect 8251 6168 8263 6171
rect 8588 6168 8616 6276
rect 9033 6273 9045 6276
rect 9079 6273 9091 6307
rect 9033 6267 9091 6273
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 9306 6264 9312 6316
rect 9364 6304 9370 6316
rect 9674 6304 9680 6316
rect 9364 6276 9409 6304
rect 9635 6276 9680 6304
rect 9364 6264 9370 6276
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 11422 6304 11428 6316
rect 11086 6276 11428 6304
rect 11422 6264 11428 6276
rect 11480 6304 11486 6316
rect 12084 6313 12112 6412
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 15838 6440 15844 6452
rect 15212 6412 15844 6440
rect 15102 6372 15108 6384
rect 14936 6344 15108 6372
rect 12069 6307 12127 6313
rect 11480 6276 11928 6304
rect 11480 6264 11486 6276
rect 10686 6196 10692 6248
rect 10744 6236 10750 6248
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 10744 6208 11713 6236
rect 10744 6196 10750 6208
rect 11701 6205 11713 6208
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 8251 6140 8616 6168
rect 8772 6140 9076 6168
rect 8251 6137 8263 6140
rect 8205 6131 8263 6137
rect 2038 6100 2044 6112
rect 992 6072 1624 6100
rect 1999 6072 2044 6100
rect 992 6060 998 6072
rect 2038 6060 2044 6072
rect 2096 6060 2102 6112
rect 2682 6060 2688 6112
rect 2740 6100 2746 6112
rect 2869 6103 2927 6109
rect 2869 6100 2881 6103
rect 2740 6072 2881 6100
rect 2740 6060 2746 6072
rect 2869 6069 2881 6072
rect 2915 6069 2927 6103
rect 2869 6063 2927 6069
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 8772 6109 8800 6140
rect 8757 6103 8815 6109
rect 8757 6100 8769 6103
rect 7616 6072 8769 6100
rect 7616 6060 7622 6072
rect 8757 6069 8769 6072
rect 8803 6069 8815 6103
rect 8938 6100 8944 6112
rect 8899 6072 8944 6100
rect 8757 6063 8815 6069
rect 8938 6060 8944 6072
rect 8996 6060 9002 6112
rect 9048 6100 9076 6140
rect 11514 6100 11520 6112
rect 9048 6072 11520 6100
rect 11514 6060 11520 6072
rect 11572 6060 11578 6112
rect 11900 6109 11928 6276
rect 12069 6273 12081 6307
rect 12115 6273 12127 6307
rect 13630 6304 13636 6316
rect 13478 6276 13636 6304
rect 12069 6267 12127 6273
rect 13630 6264 13636 6276
rect 13688 6264 13694 6316
rect 14642 6304 14648 6316
rect 14603 6276 14648 6304
rect 14642 6264 14648 6276
rect 14700 6264 14706 6316
rect 14936 6313 14964 6344
rect 15102 6332 15108 6344
rect 15160 6332 15166 6384
rect 15212 6381 15240 6412
rect 15838 6400 15844 6412
rect 15896 6400 15902 6452
rect 16666 6440 16672 6452
rect 16627 6412 16672 6440
rect 16666 6400 16672 6412
rect 16724 6400 16730 6452
rect 16850 6440 16856 6452
rect 16811 6412 16856 6440
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 17221 6443 17279 6449
rect 17221 6409 17233 6443
rect 17267 6440 17279 6443
rect 17681 6443 17739 6449
rect 17681 6440 17693 6443
rect 17267 6412 17693 6440
rect 17267 6409 17279 6412
rect 17221 6403 17279 6409
rect 17681 6409 17693 6412
rect 17727 6409 17739 6443
rect 18046 6440 18052 6452
rect 18007 6412 18052 6440
rect 17681 6403 17739 6409
rect 18046 6400 18052 6412
rect 18104 6400 18110 6452
rect 15197 6375 15255 6381
rect 15197 6341 15209 6375
rect 15243 6341 15255 6375
rect 15197 6335 15255 6341
rect 14921 6307 14979 6313
rect 14921 6273 14933 6307
rect 14967 6273 14979 6307
rect 14921 6267 14979 6273
rect 16206 6264 16212 6316
rect 16264 6304 16270 6316
rect 16666 6304 16672 6316
rect 16264 6276 16672 6304
rect 16264 6264 16270 6276
rect 16666 6264 16672 6276
rect 16724 6264 16730 6316
rect 16942 6304 16948 6316
rect 16776 6276 16948 6304
rect 11974 6196 11980 6248
rect 12032 6236 12038 6248
rect 12345 6239 12403 6245
rect 12345 6236 12357 6239
rect 12032 6208 12357 6236
rect 12032 6196 12038 6208
rect 12345 6205 12357 6208
rect 12391 6205 12403 6239
rect 12345 6199 12403 6205
rect 13648 6168 13676 6264
rect 14366 6196 14372 6248
rect 14424 6236 14430 6248
rect 16776 6236 16804 6276
rect 16942 6264 16948 6276
rect 17000 6304 17006 6316
rect 17313 6307 17371 6313
rect 17313 6304 17325 6307
rect 17000 6276 17325 6304
rect 17000 6264 17006 6276
rect 17313 6273 17325 6276
rect 17359 6273 17371 6307
rect 17313 6267 17371 6273
rect 17402 6236 17408 6248
rect 14424 6208 16804 6236
rect 17363 6208 17408 6236
rect 14424 6196 14430 6208
rect 17402 6196 17408 6208
rect 17460 6196 17466 6248
rect 17494 6196 17500 6248
rect 17552 6236 17558 6248
rect 18141 6239 18199 6245
rect 18141 6236 18153 6239
rect 17552 6208 18153 6236
rect 17552 6196 17558 6208
rect 18141 6205 18153 6208
rect 18187 6205 18199 6239
rect 18141 6199 18199 6205
rect 18233 6239 18291 6245
rect 18233 6205 18245 6239
rect 18279 6205 18291 6239
rect 18233 6199 18291 6205
rect 13648 6140 14044 6168
rect 11885 6103 11943 6109
rect 11885 6069 11897 6103
rect 11931 6100 11943 6103
rect 13648 6100 13676 6140
rect 11931 6072 13676 6100
rect 11931 6069 11943 6072
rect 11885 6063 11943 6069
rect 13722 6060 13728 6112
rect 13780 6100 13786 6112
rect 13817 6103 13875 6109
rect 13817 6100 13829 6103
rect 13780 6072 13829 6100
rect 13780 6060 13786 6072
rect 13817 6069 13829 6072
rect 13863 6069 13875 6103
rect 14016 6100 14044 6140
rect 14550 6100 14556 6112
rect 14016 6072 14556 6100
rect 13817 6063 13875 6069
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 14737 6103 14795 6109
rect 14737 6069 14749 6103
rect 14783 6100 14795 6103
rect 15286 6100 15292 6112
rect 14783 6072 15292 6100
rect 14783 6069 14795 6072
rect 14737 6063 14795 6069
rect 15286 6060 15292 6072
rect 15344 6100 15350 6112
rect 18248 6100 18276 6199
rect 15344 6072 18276 6100
rect 15344 6060 15350 6072
rect 0 6010 18860 6032
rect 0 5958 3110 6010
rect 3162 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 3302 6010
rect 3354 5958 3366 6010
rect 3418 5958 6210 6010
rect 6262 5958 6274 6010
rect 6326 5958 6338 6010
rect 6390 5958 6402 6010
rect 6454 5958 6466 6010
rect 6518 5958 9310 6010
rect 9362 5958 9374 6010
rect 9426 5958 9438 6010
rect 9490 5958 9502 6010
rect 9554 5958 9566 6010
rect 9618 5958 12410 6010
rect 12462 5958 12474 6010
rect 12526 5958 12538 6010
rect 12590 5958 12602 6010
rect 12654 5958 12666 6010
rect 12718 5958 15510 6010
rect 15562 5958 15574 6010
rect 15626 5958 15638 6010
rect 15690 5958 15702 6010
rect 15754 5958 15766 6010
rect 15818 5958 18860 6010
rect 0 5936 18860 5958
rect 2406 5896 2412 5908
rect 2367 5868 2412 5896
rect 2406 5856 2412 5868
rect 2464 5856 2470 5908
rect 3237 5899 3295 5905
rect 3237 5865 3249 5899
rect 3283 5896 3295 5899
rect 4246 5896 4252 5908
rect 3283 5868 4252 5896
rect 3283 5865 3295 5868
rect 3237 5859 3295 5865
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 5626 5896 5632 5908
rect 5587 5868 5632 5896
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 7469 5899 7527 5905
rect 7469 5865 7481 5899
rect 7515 5896 7527 5899
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 7515 5868 7849 5896
rect 7515 5865 7527 5868
rect 7469 5859 7527 5865
rect 7837 5865 7849 5868
rect 7883 5896 7895 5899
rect 8478 5896 8484 5908
rect 7883 5868 8484 5896
rect 7883 5865 7895 5868
rect 7837 5859 7895 5865
rect 8478 5856 8484 5868
rect 8536 5856 8542 5908
rect 10597 5899 10655 5905
rect 10597 5865 10609 5899
rect 10643 5896 10655 5899
rect 15378 5896 15384 5908
rect 10643 5868 15384 5896
rect 10643 5865 10655 5868
rect 10597 5859 10655 5865
rect 2038 5788 2044 5840
rect 2096 5828 2102 5840
rect 2096 5800 3740 5828
rect 2096 5788 2102 5800
rect 750 5692 756 5704
rect 711 5664 756 5692
rect 750 5652 756 5664
rect 808 5652 814 5704
rect 2314 5692 2320 5704
rect 2275 5664 2320 5692
rect 2314 5652 2320 5664
rect 2372 5652 2378 5704
rect 2884 5701 2912 5800
rect 2961 5763 3019 5769
rect 2961 5729 2973 5763
rect 3007 5760 3019 5763
rect 3421 5763 3479 5769
rect 3421 5760 3433 5763
rect 3007 5732 3433 5760
rect 3007 5729 3019 5732
rect 2961 5723 3019 5729
rect 3421 5729 3433 5732
rect 3467 5729 3479 5763
rect 3421 5723 3479 5729
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 3050 5652 3056 5704
rect 3108 5692 3114 5704
rect 3712 5701 3740 5800
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 4120 5800 5028 5828
rect 4120 5788 4126 5800
rect 5000 5769 5028 5800
rect 4985 5763 5043 5769
rect 4985 5729 4997 5763
rect 5031 5729 5043 5763
rect 4985 5723 5043 5729
rect 3329 5695 3387 5701
rect 3329 5692 3341 5695
rect 3108 5664 3341 5692
rect 3108 5652 3114 5664
rect 3329 5661 3341 5664
rect 3375 5661 3387 5695
rect 3329 5655 3387 5661
rect 3513 5695 3571 5701
rect 3513 5661 3525 5695
rect 3559 5661 3571 5695
rect 3513 5655 3571 5661
rect 3697 5695 3755 5701
rect 3697 5661 3709 5695
rect 3743 5661 3755 5695
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3697 5655 3755 5661
rect 3804 5664 3985 5692
rect 2332 5624 2360 5652
rect 3528 5624 3556 5655
rect 3804 5624 3832 5664
rect 3973 5661 3985 5664
rect 4019 5692 4031 5695
rect 4062 5692 4068 5704
rect 4019 5664 4068 5692
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 6089 5695 6147 5701
rect 6089 5661 6101 5695
rect 6135 5692 6147 5695
rect 6822 5692 6828 5704
rect 6135 5664 6828 5692
rect 6135 5661 6147 5664
rect 6089 5655 6147 5661
rect 2332 5596 3832 5624
rect 3878 5584 3884 5636
rect 3936 5624 3942 5636
rect 4540 5624 4568 5655
rect 6822 5652 6828 5664
rect 6880 5692 6886 5704
rect 7466 5692 7472 5704
rect 6880 5664 7472 5692
rect 6880 5652 6886 5664
rect 7466 5652 7472 5664
rect 7524 5652 7530 5704
rect 7558 5652 7564 5704
rect 7616 5692 7622 5704
rect 10413 5695 10471 5701
rect 7616 5664 7661 5692
rect 7616 5652 7622 5664
rect 10413 5661 10425 5695
rect 10459 5692 10471 5695
rect 10612 5692 10640 5859
rect 15378 5856 15384 5868
rect 15436 5856 15442 5908
rect 16942 5856 16948 5908
rect 17000 5896 17006 5908
rect 17819 5899 17877 5905
rect 17819 5896 17831 5899
rect 17000 5868 17831 5896
rect 17000 5856 17006 5868
rect 17819 5865 17831 5868
rect 17865 5865 17877 5899
rect 17819 5859 17877 5865
rect 11149 5831 11207 5837
rect 11149 5797 11161 5831
rect 11195 5828 11207 5831
rect 11238 5828 11244 5840
rect 11195 5800 11244 5828
rect 11195 5797 11207 5800
rect 11149 5791 11207 5797
rect 11238 5788 11244 5800
rect 11296 5788 11302 5840
rect 11974 5828 11980 5840
rect 11935 5800 11980 5828
rect 11974 5788 11980 5800
rect 12032 5788 12038 5840
rect 12253 5831 12311 5837
rect 12253 5797 12265 5831
rect 12299 5797 12311 5831
rect 12253 5791 12311 5797
rect 13081 5831 13139 5837
rect 13081 5797 13093 5831
rect 13127 5828 13139 5831
rect 14645 5831 14703 5837
rect 14645 5828 14657 5831
rect 13127 5800 14657 5828
rect 13127 5797 13139 5800
rect 13081 5791 13139 5797
rect 14645 5797 14657 5800
rect 14691 5797 14703 5831
rect 14645 5791 14703 5797
rect 10459 5664 10640 5692
rect 11793 5695 11851 5701
rect 10459 5661 10471 5664
rect 10413 5655 10471 5661
rect 11793 5661 11805 5695
rect 11839 5692 11851 5695
rect 12268 5692 12296 5791
rect 12805 5763 12863 5769
rect 12805 5760 12817 5763
rect 11839 5664 12296 5692
rect 12544 5732 12817 5760
rect 11839 5661 11851 5664
rect 11793 5655 11851 5661
rect 5166 5624 5172 5636
rect 3936 5596 4568 5624
rect 5079 5596 5172 5624
rect 3936 5584 3942 5596
rect 5166 5584 5172 5596
rect 5224 5624 5230 5636
rect 6356 5627 6414 5633
rect 6356 5624 6368 5627
rect 5224 5596 6368 5624
rect 5224 5584 5230 5596
rect 6356 5593 6368 5596
rect 6402 5624 6414 5627
rect 7576 5624 7604 5652
rect 8662 5624 8668 5636
rect 6402 5596 7604 5624
rect 8623 5596 8668 5624
rect 6402 5593 6414 5596
rect 6356 5587 6414 5593
rect 8662 5584 8668 5596
rect 8720 5624 8726 5636
rect 10965 5627 11023 5633
rect 10965 5624 10977 5627
rect 8720 5596 10977 5624
rect 8720 5584 8726 5596
rect 10965 5593 10977 5596
rect 11011 5593 11023 5627
rect 10965 5587 11023 5593
rect 474 5516 480 5568
rect 532 5556 538 5568
rect 661 5559 719 5565
rect 661 5556 673 5559
rect 532 5528 673 5556
rect 532 5516 538 5528
rect 661 5525 673 5528
rect 707 5525 719 5559
rect 661 5519 719 5525
rect 2406 5516 2412 5568
rect 2464 5556 2470 5568
rect 2866 5556 2872 5568
rect 2464 5528 2872 5556
rect 2464 5516 2470 5528
rect 2866 5516 2872 5528
rect 2924 5516 2930 5568
rect 3970 5556 3976 5568
rect 3931 5528 3976 5556
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 5258 5516 5264 5568
rect 5316 5556 5322 5568
rect 8021 5559 8079 5565
rect 5316 5528 5361 5556
rect 5316 5516 5322 5528
rect 8021 5525 8033 5559
rect 8067 5556 8079 5559
rect 9030 5556 9036 5568
rect 8067 5528 9036 5556
rect 8067 5525 8079 5528
rect 8021 5519 8079 5525
rect 9030 5516 9036 5528
rect 9088 5516 9094 5568
rect 10778 5516 10784 5568
rect 10836 5556 10842 5568
rect 12544 5556 12572 5732
rect 12805 5729 12817 5732
rect 12851 5760 12863 5763
rect 12894 5760 12900 5772
rect 12851 5732 12900 5760
rect 12851 5729 12863 5732
rect 12805 5723 12863 5729
rect 12894 5720 12900 5732
rect 12952 5760 12958 5772
rect 13722 5760 13728 5772
rect 12952 5732 13728 5760
rect 12952 5720 12958 5732
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 14277 5763 14335 5769
rect 14277 5760 14289 5763
rect 13832 5732 14289 5760
rect 12713 5695 12771 5701
rect 12713 5661 12725 5695
rect 12759 5692 12771 5695
rect 13541 5695 13599 5701
rect 13541 5692 13553 5695
rect 12759 5664 13553 5692
rect 12759 5661 12771 5664
rect 12713 5655 12771 5661
rect 13541 5661 13553 5664
rect 13587 5692 13599 5695
rect 13630 5692 13636 5704
rect 13587 5664 13636 5692
rect 13587 5661 13599 5664
rect 13541 5655 13599 5661
rect 13630 5652 13636 5664
rect 13688 5652 13694 5704
rect 13832 5701 13860 5732
rect 14277 5729 14289 5732
rect 14323 5760 14335 5763
rect 14366 5760 14372 5772
rect 14323 5732 14372 5760
rect 14323 5729 14335 5732
rect 14277 5723 14335 5729
rect 14366 5720 14372 5732
rect 14424 5720 14430 5772
rect 15286 5760 15292 5772
rect 15247 5732 15292 5760
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 16393 5763 16451 5769
rect 16393 5729 16405 5763
rect 16439 5760 16451 5763
rect 16574 5760 16580 5772
rect 16439 5732 16580 5760
rect 16439 5729 16451 5732
rect 16393 5723 16451 5729
rect 16574 5720 16580 5732
rect 16632 5720 16638 5772
rect 13811 5695 13869 5701
rect 13811 5661 13823 5695
rect 13857 5661 13869 5695
rect 14158 5695 14216 5701
rect 14158 5692 14170 5695
rect 13811 5655 13869 5661
rect 13924 5664 14170 5692
rect 12621 5627 12679 5633
rect 12621 5593 12633 5627
rect 12667 5624 12679 5627
rect 13081 5627 13139 5633
rect 13081 5624 13093 5627
rect 12667 5596 13093 5624
rect 12667 5593 12679 5596
rect 12621 5587 12679 5593
rect 13081 5593 13093 5596
rect 13127 5593 13139 5627
rect 13648 5624 13676 5652
rect 13924 5624 13952 5664
rect 14158 5661 14170 5664
rect 14204 5661 14216 5695
rect 14158 5655 14216 5661
rect 14458 5652 14464 5704
rect 14516 5692 14522 5704
rect 15378 5692 15384 5704
rect 14516 5664 15384 5692
rect 14516 5652 14522 5664
rect 15378 5652 15384 5664
rect 15436 5692 15442 5704
rect 16025 5695 16083 5701
rect 16025 5692 16037 5695
rect 15436 5664 16037 5692
rect 15436 5652 15442 5664
rect 16025 5661 16037 5664
rect 16071 5661 16083 5695
rect 16025 5655 16083 5661
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5692 18291 5695
rect 18506 5692 18512 5704
rect 18279 5664 18512 5692
rect 18279 5661 18291 5664
rect 18233 5655 18291 5661
rect 18506 5652 18512 5664
rect 18564 5652 18570 5704
rect 15105 5627 15163 5633
rect 15105 5624 15117 5627
rect 13648 5596 13952 5624
rect 14568 5596 15117 5624
rect 13081 5587 13139 5593
rect 10836 5528 12572 5556
rect 10836 5516 10842 5528
rect 13630 5516 13636 5568
rect 13688 5556 13694 5568
rect 14568 5565 14596 5596
rect 15105 5593 15117 5596
rect 15151 5593 15163 5627
rect 15105 5587 15163 5593
rect 13817 5559 13875 5565
rect 13817 5556 13829 5559
rect 13688 5528 13829 5556
rect 13688 5516 13694 5528
rect 13817 5525 13829 5528
rect 13863 5525 13875 5559
rect 13817 5519 13875 5525
rect 14553 5559 14611 5565
rect 14553 5525 14565 5559
rect 14599 5525 14611 5559
rect 15010 5556 15016 5568
rect 14971 5528 15016 5556
rect 14553 5519 14611 5525
rect 15010 5516 15016 5528
rect 15068 5516 15074 5568
rect 15654 5516 15660 5568
rect 15712 5556 15718 5568
rect 15841 5559 15899 5565
rect 15841 5556 15853 5559
rect 15712 5528 15853 5556
rect 15712 5516 15718 5528
rect 15841 5525 15853 5528
rect 15887 5556 15899 5559
rect 16666 5556 16672 5568
rect 15887 5528 16672 5556
rect 15887 5525 15899 5528
rect 15841 5519 15899 5525
rect 16666 5516 16672 5528
rect 16724 5556 16730 5568
rect 16776 5556 16804 5610
rect 18322 5556 18328 5568
rect 16724 5528 16804 5556
rect 18283 5528 18328 5556
rect 16724 5516 16730 5528
rect 18322 5516 18328 5528
rect 18380 5516 18386 5568
rect 0 5466 18860 5488
rect 0 5414 4660 5466
rect 4712 5414 4724 5466
rect 4776 5414 4788 5466
rect 4840 5414 4852 5466
rect 4904 5414 4916 5466
rect 4968 5414 7760 5466
rect 7812 5414 7824 5466
rect 7876 5414 7888 5466
rect 7940 5414 7952 5466
rect 8004 5414 8016 5466
rect 8068 5414 10860 5466
rect 10912 5414 10924 5466
rect 10976 5414 10988 5466
rect 11040 5414 11052 5466
rect 11104 5414 11116 5466
rect 11168 5414 13960 5466
rect 14012 5414 14024 5466
rect 14076 5414 14088 5466
rect 14140 5414 14152 5466
rect 14204 5414 14216 5466
rect 14268 5414 17060 5466
rect 17112 5414 17124 5466
rect 17176 5414 17188 5466
rect 17240 5414 17252 5466
rect 17304 5414 17316 5466
rect 17368 5414 18860 5466
rect 0 5392 18860 5414
rect 2314 5361 2320 5364
rect 2271 5355 2320 5361
rect 2271 5321 2283 5355
rect 2317 5321 2320 5355
rect 2271 5315 2320 5321
rect 2314 5312 2320 5315
rect 2372 5312 2378 5364
rect 4433 5355 4491 5361
rect 4433 5321 4445 5355
rect 4479 5352 4491 5355
rect 5258 5352 5264 5364
rect 4479 5324 5264 5352
rect 4479 5321 4491 5324
rect 4433 5315 4491 5321
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 8849 5355 8907 5361
rect 8849 5321 8861 5355
rect 8895 5352 8907 5355
rect 10778 5352 10784 5364
rect 8895 5324 9352 5352
rect 8895 5321 8907 5324
rect 8849 5315 8907 5321
rect 1854 5244 1860 5296
rect 1912 5284 1918 5296
rect 2590 5284 2596 5296
rect 1912 5256 2596 5284
rect 1912 5244 1918 5256
rect 2590 5244 2596 5256
rect 2648 5244 2654 5296
rect 7650 5244 7656 5296
rect 7708 5244 7714 5296
rect 8938 5244 8944 5296
rect 8996 5284 9002 5296
rect 9324 5293 9352 5324
rect 9416 5324 10784 5352
rect 9125 5287 9183 5293
rect 9125 5284 9137 5287
rect 8996 5256 9137 5284
rect 8996 5244 9002 5256
rect 9125 5253 9137 5256
rect 9171 5253 9183 5287
rect 9125 5247 9183 5253
rect 9309 5287 9367 5293
rect 9309 5253 9321 5287
rect 9355 5253 9367 5287
rect 9309 5247 9367 5253
rect 474 5216 480 5228
rect 435 5188 480 5216
rect 474 5176 480 5188
rect 532 5176 538 5228
rect 845 5219 903 5225
rect 845 5185 857 5219
rect 891 5216 903 5219
rect 934 5216 940 5228
rect 891 5188 940 5216
rect 891 5185 903 5188
rect 845 5179 903 5185
rect 934 5176 940 5188
rect 992 5176 998 5228
rect 4062 5216 4068 5228
rect 4023 5188 4068 5216
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 7466 5216 7472 5228
rect 7427 5188 7472 5216
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 7668 5216 7696 5244
rect 7736 5219 7794 5225
rect 7736 5216 7748 5219
rect 7668 5188 7748 5216
rect 7736 5185 7748 5188
rect 7782 5216 7794 5219
rect 9030 5216 9036 5228
rect 7782 5188 8524 5216
rect 8991 5188 9036 5216
rect 7782 5185 7794 5188
rect 7736 5179 7794 5185
rect 3050 5108 3056 5160
rect 3108 5148 3114 5160
rect 3878 5148 3884 5160
rect 3108 5120 3884 5148
rect 3108 5108 3114 5120
rect 3878 5108 3884 5120
rect 3936 5148 3942 5160
rect 3973 5151 4031 5157
rect 3973 5148 3985 5151
rect 3936 5120 3985 5148
rect 3936 5108 3942 5120
rect 3973 5117 3985 5120
rect 4019 5117 4031 5151
rect 8496 5148 8524 5188
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 9416 5148 9444 5324
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 15654 5284 15660 5296
rect 8496 5120 9444 5148
rect 9692 5256 10626 5284
rect 14752 5256 15660 5284
rect 3973 5111 4031 5117
rect 8846 5040 8852 5092
rect 8904 5080 8910 5092
rect 9033 5083 9091 5089
rect 9033 5080 9045 5083
rect 8904 5052 9045 5080
rect 8904 5040 8910 5052
rect 9033 5049 9045 5052
rect 9079 5049 9091 5083
rect 9033 5043 9091 5049
rect 2590 5012 2596 5024
rect 2551 4984 2596 5012
rect 2590 4972 2596 4984
rect 2648 4972 2654 5024
rect 9214 4972 9220 5024
rect 9272 5012 9278 5024
rect 9692 5021 9720 5256
rect 13449 5219 13507 5225
rect 13449 5185 13461 5219
rect 13495 5216 13507 5219
rect 13814 5216 13820 5228
rect 13495 5188 13820 5216
rect 13495 5185 13507 5188
rect 13449 5179 13507 5185
rect 13814 5176 13820 5188
rect 13872 5176 13878 5228
rect 9861 5151 9919 5157
rect 9861 5117 9873 5151
rect 9907 5148 9919 5151
rect 10137 5151 10195 5157
rect 9907 5120 9996 5148
rect 9907 5117 9919 5120
rect 9861 5111 9919 5117
rect 9968 5024 9996 5120
rect 10137 5117 10149 5151
rect 10183 5148 10195 5151
rect 11146 5148 11152 5160
rect 10183 5120 11152 5148
rect 10183 5117 10195 5120
rect 10137 5111 10195 5117
rect 11146 5108 11152 5120
rect 11204 5108 11210 5160
rect 13541 5151 13599 5157
rect 13541 5117 13553 5151
rect 13587 5148 13599 5151
rect 13630 5148 13636 5160
rect 13587 5120 13636 5148
rect 13587 5117 13599 5120
rect 13541 5111 13599 5117
rect 13630 5108 13636 5120
rect 13688 5108 13694 5160
rect 9677 5015 9735 5021
rect 9677 5012 9689 5015
rect 9272 4984 9689 5012
rect 9272 4972 9278 4984
rect 9677 4981 9689 4984
rect 9723 4981 9735 5015
rect 9950 5012 9956 5024
rect 9863 4984 9956 5012
rect 9677 4975 9735 4981
rect 9950 4972 9956 4984
rect 10008 5012 10014 5024
rect 11238 5012 11244 5024
rect 10008 4984 11244 5012
rect 10008 4972 10014 4984
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 11514 4972 11520 5024
rect 11572 5012 11578 5024
rect 11609 5015 11667 5021
rect 11609 5012 11621 5015
rect 11572 4984 11621 5012
rect 11572 4972 11578 4984
rect 11609 4981 11621 4984
rect 11655 4981 11667 5015
rect 13814 5012 13820 5024
rect 13775 4984 13820 5012
rect 11609 4975 11667 4981
rect 13814 4972 13820 4984
rect 13872 4972 13878 5024
rect 14550 4972 14556 5024
rect 14608 5012 14614 5024
rect 14752 5021 14780 5256
rect 15654 5244 15660 5256
rect 15712 5244 15718 5296
rect 17221 5287 17279 5293
rect 17221 5253 17233 5287
rect 17267 5284 17279 5287
rect 17494 5284 17500 5296
rect 17267 5256 17500 5284
rect 17267 5253 17279 5256
rect 17221 5247 17279 5253
rect 17494 5244 17500 5256
rect 17552 5244 17558 5296
rect 14918 5216 14924 5228
rect 14879 5188 14924 5216
rect 14918 5176 14924 5188
rect 14976 5176 14982 5228
rect 16942 5216 16948 5228
rect 16903 5188 16948 5216
rect 16942 5176 16948 5188
rect 17000 5176 17006 5228
rect 15197 5151 15255 5157
rect 15197 5117 15209 5151
rect 15243 5148 15255 5151
rect 18322 5148 18328 5160
rect 15243 5120 18328 5148
rect 15243 5117 15255 5120
rect 15197 5111 15255 5117
rect 18322 5108 18328 5120
rect 18380 5108 18386 5160
rect 14737 5015 14795 5021
rect 14737 5012 14749 5015
rect 14608 4984 14749 5012
rect 14608 4972 14614 4984
rect 14737 4981 14749 4984
rect 14783 4981 14795 5015
rect 14737 4975 14795 4981
rect 16669 5015 16727 5021
rect 16669 4981 16681 5015
rect 16715 5012 16727 5015
rect 16850 5012 16856 5024
rect 16715 4984 16856 5012
rect 16715 4981 16727 4984
rect 16669 4975 16727 4981
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 0 4922 18860 4944
rect 0 4870 3110 4922
rect 3162 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 3302 4922
rect 3354 4870 3366 4922
rect 3418 4870 6210 4922
rect 6262 4870 6274 4922
rect 6326 4870 6338 4922
rect 6390 4870 6402 4922
rect 6454 4870 6466 4922
rect 6518 4870 9310 4922
rect 9362 4870 9374 4922
rect 9426 4870 9438 4922
rect 9490 4870 9502 4922
rect 9554 4870 9566 4922
rect 9618 4870 12410 4922
rect 12462 4870 12474 4922
rect 12526 4870 12538 4922
rect 12590 4870 12602 4922
rect 12654 4870 12666 4922
rect 12718 4870 15510 4922
rect 15562 4870 15574 4922
rect 15626 4870 15638 4922
rect 15690 4870 15702 4922
rect 15754 4870 15766 4922
rect 15818 4870 18860 4922
rect 0 4848 18860 4870
rect 11146 4808 11152 4820
rect 11107 4780 11152 4808
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 13725 4811 13783 4817
rect 13725 4777 13737 4811
rect 13771 4808 13783 4811
rect 13906 4808 13912 4820
rect 13771 4780 13912 4808
rect 13771 4777 13783 4780
rect 13725 4771 13783 4777
rect 13906 4768 13912 4780
rect 13964 4768 13970 4820
rect 11793 4743 11851 4749
rect 11793 4740 11805 4743
rect 11624 4712 11805 4740
rect 2958 4672 2964 4684
rect 2746 4644 2964 4672
rect 753 4607 811 4613
rect 753 4573 765 4607
rect 799 4604 811 4607
rect 2746 4604 2774 4644
rect 2958 4632 2964 4644
rect 3016 4672 3022 4684
rect 3697 4675 3755 4681
rect 3697 4672 3709 4675
rect 3016 4644 3709 4672
rect 3016 4632 3022 4644
rect 3697 4641 3709 4644
rect 3743 4672 3755 4675
rect 6089 4675 6147 4681
rect 6089 4672 6101 4675
rect 3743 4644 6101 4672
rect 3743 4641 3755 4644
rect 3697 4635 3755 4641
rect 6089 4641 6101 4644
rect 6135 4672 6147 4675
rect 6914 4672 6920 4684
rect 6135 4644 6920 4672
rect 6135 4641 6147 4644
rect 6089 4635 6147 4641
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 8481 4675 8539 4681
rect 8481 4641 8493 4675
rect 8527 4672 8539 4675
rect 9950 4672 9956 4684
rect 8527 4644 9956 4672
rect 8527 4641 8539 4644
rect 8481 4635 8539 4641
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 11624 4681 11652 4712
rect 11793 4709 11805 4712
rect 11839 4709 11851 4743
rect 11793 4703 11851 4709
rect 11609 4675 11667 4681
rect 11609 4641 11621 4675
rect 11655 4641 11667 4675
rect 11609 4635 11667 4641
rect 11716 4644 12388 4672
rect 6454 4604 6460 4616
rect 799 4576 2774 4604
rect 6415 4576 6460 4604
rect 799 4573 811 4576
rect 753 4567 811 4573
rect 6454 4564 6460 4576
rect 6512 4564 6518 4616
rect 7650 4564 7656 4616
rect 7708 4604 7714 4616
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7708 4576 7941 4604
rect 7708 4564 7714 4576
rect 7929 4573 7941 4576
rect 7975 4604 7987 4607
rect 8021 4607 8079 4613
rect 8021 4604 8033 4607
rect 7975 4576 8033 4604
rect 7975 4573 7987 4576
rect 7929 4567 7987 4573
rect 8021 4573 8033 4576
rect 8067 4573 8079 4607
rect 11514 4604 11520 4616
rect 11475 4576 11520 4604
rect 8021 4567 8079 4573
rect 11514 4564 11520 4576
rect 11572 4604 11578 4616
rect 11716 4604 11744 4644
rect 12360 4613 12388 4644
rect 13814 4632 13820 4684
rect 13872 4672 13878 4684
rect 15197 4675 15255 4681
rect 15197 4672 15209 4675
rect 13872 4644 15209 4672
rect 13872 4632 13878 4644
rect 15197 4641 15209 4644
rect 15243 4641 15255 4675
rect 15470 4672 15476 4684
rect 15431 4644 15476 4672
rect 15197 4635 15255 4641
rect 15470 4632 15476 4644
rect 15528 4632 15534 4684
rect 16850 4632 16856 4684
rect 16908 4672 16914 4684
rect 17589 4675 17647 4681
rect 17589 4672 17601 4675
rect 16908 4644 17601 4672
rect 16908 4632 16914 4644
rect 17589 4641 17601 4644
rect 17635 4641 17647 4675
rect 17589 4635 17647 4641
rect 11572 4576 11744 4604
rect 11793 4607 11851 4613
rect 11572 4564 11578 4576
rect 11793 4573 11805 4607
rect 11839 4573 11851 4607
rect 11793 4567 11851 4573
rect 11885 4607 11943 4613
rect 11885 4573 11897 4607
rect 11931 4604 11943 4607
rect 12161 4607 12219 4613
rect 12161 4604 12173 4607
rect 11931 4576 12173 4604
rect 11931 4573 11943 4576
rect 11885 4567 11943 4573
rect 12161 4573 12173 4576
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 12345 4607 12403 4613
rect 12345 4573 12357 4607
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 3510 4496 3516 4548
rect 3568 4536 3574 4548
rect 3973 4539 4031 4545
rect 3973 4536 3985 4539
rect 3568 4508 3985 4536
rect 3568 4496 3574 4508
rect 3973 4505 3985 4508
rect 4019 4505 4031 4539
rect 8386 4536 8392 4548
rect 5198 4522 5948 4536
rect 7498 4522 8392 4536
rect 3973 4499 4031 4505
rect 5184 4508 5948 4522
rect 474 4428 480 4480
rect 532 4468 538 4480
rect 661 4471 719 4477
rect 661 4468 673 4471
rect 532 4440 673 4468
rect 532 4428 538 4440
rect 661 4437 673 4440
rect 707 4437 719 4471
rect 661 4431 719 4437
rect 2501 4471 2559 4477
rect 2501 4437 2513 4471
rect 2547 4468 2559 4471
rect 2590 4468 2596 4480
rect 2547 4440 2596 4468
rect 2547 4437 2559 4440
rect 2501 4431 2559 4437
rect 2590 4428 2596 4440
rect 2648 4468 2654 4480
rect 3421 4471 3479 4477
rect 3421 4468 3433 4471
rect 2648 4440 3433 4468
rect 2648 4428 2654 4440
rect 3421 4437 3433 4440
rect 3467 4468 3479 4471
rect 5184 4468 5212 4508
rect 5442 4468 5448 4480
rect 3467 4440 5212 4468
rect 5403 4440 5448 4468
rect 3467 4437 3479 4440
rect 3421 4431 3479 4437
rect 5442 4428 5448 4440
rect 5500 4428 5506 4480
rect 5920 4477 5948 4508
rect 7484 4508 8392 4522
rect 5905 4471 5963 4477
rect 5905 4437 5917 4471
rect 5951 4468 5963 4471
rect 7484 4468 7512 4508
rect 8386 4496 8392 4508
rect 8444 4536 8450 4548
rect 8757 4539 8815 4545
rect 8444 4508 8708 4536
rect 8444 4496 8450 4508
rect 5951 4440 7512 4468
rect 8205 4471 8263 4477
rect 5951 4437 5963 4440
rect 5905 4431 5963 4437
rect 8205 4437 8217 4471
rect 8251 4468 8263 4471
rect 8570 4468 8576 4480
rect 8251 4440 8576 4468
rect 8251 4437 8263 4440
rect 8205 4431 8263 4437
rect 8570 4428 8576 4440
rect 8628 4428 8634 4480
rect 8680 4468 8708 4508
rect 8757 4505 8769 4539
rect 8803 4536 8815 4539
rect 8846 4536 8852 4548
rect 8803 4508 8852 4536
rect 8803 4505 8815 4508
rect 8757 4499 8815 4505
rect 8846 4496 8852 4508
rect 8904 4496 8910 4548
rect 9214 4496 9220 4548
rect 9272 4496 9278 4548
rect 11606 4496 11612 4548
rect 11664 4536 11670 4548
rect 11808 4536 11836 4567
rect 11664 4508 11836 4536
rect 11664 4496 11670 4508
rect 9232 4468 9260 4496
rect 8680 4440 9260 4468
rect 9766 4428 9772 4480
rect 9824 4468 9830 4480
rect 10229 4471 10287 4477
rect 10229 4468 10241 4471
rect 9824 4440 10241 4468
rect 9824 4428 9830 4440
rect 10229 4437 10241 4440
rect 10275 4468 10287 4471
rect 11900 4468 11928 4567
rect 17862 4564 17868 4616
rect 17920 4604 17926 4616
rect 17920 4576 17965 4604
rect 17920 4564 17926 4576
rect 11974 4496 11980 4548
rect 12032 4536 12038 4548
rect 12069 4539 12127 4545
rect 12069 4536 12081 4539
rect 12032 4508 12081 4536
rect 12032 4496 12038 4508
rect 12069 4505 12081 4508
rect 12115 4505 12127 4539
rect 12069 4499 12127 4505
rect 12250 4468 12256 4480
rect 10275 4440 11928 4468
rect 12211 4440 12256 4468
rect 10275 4437 10287 4440
rect 10229 4431 10287 4437
rect 12250 4428 12256 4440
rect 12308 4428 12314 4480
rect 13170 4428 13176 4480
rect 13228 4468 13234 4480
rect 13541 4471 13599 4477
rect 13541 4468 13553 4471
rect 13228 4440 13553 4468
rect 13228 4428 13234 4440
rect 13541 4437 13553 4440
rect 13587 4468 13599 4471
rect 14016 4468 14044 4522
rect 15194 4496 15200 4548
rect 15252 4536 15258 4548
rect 15841 4539 15899 4545
rect 15841 4536 15853 4539
rect 15252 4508 15853 4536
rect 15252 4496 15258 4508
rect 15841 4505 15853 4508
rect 15887 4505 15899 4539
rect 15841 4499 15899 4505
rect 14550 4468 14556 4480
rect 13587 4440 14556 4468
rect 13587 4437 13599 4440
rect 13541 4431 13599 4437
rect 14550 4428 14556 4440
rect 14608 4468 14614 4480
rect 15657 4471 15715 4477
rect 15657 4468 15669 4471
rect 14608 4440 15669 4468
rect 14608 4428 14614 4440
rect 15657 4437 15669 4440
rect 15703 4468 15715 4471
rect 16408 4468 16436 4522
rect 15703 4440 16436 4468
rect 15703 4437 15715 4440
rect 15657 4431 15715 4437
rect 0 4378 18860 4400
rect 0 4326 4660 4378
rect 4712 4326 4724 4378
rect 4776 4326 4788 4378
rect 4840 4326 4852 4378
rect 4904 4326 4916 4378
rect 4968 4326 7760 4378
rect 7812 4326 7824 4378
rect 7876 4326 7888 4378
rect 7940 4326 7952 4378
rect 8004 4326 8016 4378
rect 8068 4326 10860 4378
rect 10912 4326 10924 4378
rect 10976 4326 10988 4378
rect 11040 4326 11052 4378
rect 11104 4326 11116 4378
rect 11168 4326 13960 4378
rect 14012 4326 14024 4378
rect 14076 4326 14088 4378
rect 14140 4326 14152 4378
rect 14204 4326 14216 4378
rect 14268 4326 17060 4378
rect 17112 4326 17124 4378
rect 17176 4326 17188 4378
rect 17240 4326 17252 4378
rect 17304 4326 17316 4378
rect 17368 4326 18860 4378
rect 0 4304 18860 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 2501 4267 2559 4273
rect 2501 4264 2513 4267
rect 2464 4236 2513 4264
rect 2464 4224 2470 4236
rect 2501 4233 2513 4236
rect 2547 4233 2559 4267
rect 3510 4264 3516 4276
rect 3471 4236 3516 4264
rect 2501 4227 2559 4233
rect 3510 4224 3516 4236
rect 3568 4224 3574 4276
rect 3973 4267 4031 4273
rect 3973 4233 3985 4267
rect 4019 4264 4031 4267
rect 4338 4264 4344 4276
rect 4019 4236 4344 4264
rect 4019 4233 4031 4236
rect 3973 4227 4031 4233
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 6273 4267 6331 4273
rect 6273 4233 6285 4267
rect 6319 4264 6331 4267
rect 6454 4264 6460 4276
rect 6319 4236 6460 4264
rect 6319 4233 6331 4236
rect 6273 4227 6331 4233
rect 6454 4224 6460 4236
rect 6512 4224 6518 4276
rect 7653 4267 7711 4273
rect 7653 4233 7665 4267
rect 7699 4264 7711 4267
rect 8113 4267 8171 4273
rect 8113 4264 8125 4267
rect 7699 4236 8125 4264
rect 7699 4233 7711 4236
rect 7653 4227 7711 4233
rect 8113 4233 8125 4236
rect 8159 4233 8171 4267
rect 8113 4227 8171 4233
rect 8481 4267 8539 4273
rect 8481 4233 8493 4267
rect 8527 4264 8539 4267
rect 8527 4236 8800 4264
rect 8527 4233 8539 4236
rect 8481 4227 8539 4233
rect 2590 4196 2596 4208
rect 1886 4168 2596 4196
rect 2590 4156 2596 4168
rect 2648 4156 2654 4208
rect 2866 4196 2872 4208
rect 2700 4168 2872 4196
rect 474 4128 480 4140
rect 435 4100 480 4128
rect 474 4088 480 4100
rect 532 4088 538 4140
rect 845 4063 903 4069
rect 845 4029 857 4063
rect 891 4060 903 4063
rect 2406 4060 2412 4072
rect 891 4032 2412 4060
rect 891 4029 903 4032
rect 845 4023 903 4029
rect 2406 4020 2412 4032
rect 2464 4020 2470 4072
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4060 2559 4063
rect 2700 4060 2728 4168
rect 2866 4156 2872 4168
rect 2924 4196 2930 4208
rect 3329 4199 3387 4205
rect 3329 4196 3341 4199
rect 2924 4168 3341 4196
rect 2924 4156 2930 4168
rect 3329 4165 3341 4168
rect 3375 4165 3387 4199
rect 7009 4199 7067 4205
rect 3329 4159 3387 4165
rect 3528 4168 5212 4196
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4097 2835 4131
rect 2777 4091 2835 4097
rect 2547 4032 2728 4060
rect 2792 4060 2820 4091
rect 3050 4088 3056 4140
rect 3108 4128 3114 4140
rect 3237 4131 3295 4137
rect 3108 4100 3153 4128
rect 3108 4088 3114 4100
rect 3237 4097 3249 4131
rect 3283 4126 3295 4131
rect 3528 4128 3556 4168
rect 3786 4128 3792 4140
rect 3344 4126 3556 4128
rect 3283 4100 3556 4126
rect 3747 4100 3792 4128
rect 3283 4098 3372 4100
rect 3283 4097 3295 4098
rect 3237 4091 3295 4097
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 3896 4137 3924 4168
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4097 3939 4131
rect 3881 4091 3939 4097
rect 3988 4118 4108 4128
rect 4157 4121 4215 4127
rect 4157 4118 4169 4121
rect 3988 4100 4169 4118
rect 2961 4063 3019 4069
rect 2961 4060 2973 4063
rect 2792 4032 2973 4060
rect 2547 4029 2559 4032
rect 2501 4023 2559 4029
rect 2961 4029 2973 4032
rect 3007 4060 3019 4063
rect 3988 4060 4016 4100
rect 4080 4090 4169 4100
rect 4157 4087 4169 4090
rect 4203 4087 4215 4121
rect 4338 4088 4344 4140
rect 4396 4128 4402 4140
rect 4982 4128 4988 4140
rect 4396 4100 4441 4128
rect 4943 4100 4988 4128
rect 4396 4088 4402 4100
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 5184 4137 5212 4168
rect 7009 4165 7021 4199
rect 7055 4196 7067 4199
rect 8662 4196 8668 4208
rect 7055 4168 8668 4196
rect 7055 4165 7067 4168
rect 7009 4159 7067 4165
rect 8662 4156 8668 4168
rect 8720 4156 8726 4208
rect 8772 4196 8800 4236
rect 8846 4224 8852 4276
rect 8904 4264 8910 4276
rect 8941 4267 8999 4273
rect 8941 4264 8953 4267
rect 8904 4236 8953 4264
rect 8904 4224 8910 4236
rect 8941 4233 8953 4236
rect 8987 4233 8999 4267
rect 8941 4227 8999 4233
rect 10045 4267 10103 4273
rect 10045 4233 10057 4267
rect 10091 4264 10103 4267
rect 10505 4267 10563 4273
rect 10505 4264 10517 4267
rect 10091 4236 10517 4264
rect 10091 4233 10103 4236
rect 10045 4227 10103 4233
rect 10505 4233 10517 4236
rect 10551 4233 10563 4267
rect 14734 4264 14740 4276
rect 10505 4227 10563 4233
rect 10612 4236 14740 4264
rect 10612 4196 10640 4236
rect 14734 4224 14740 4236
rect 14792 4224 14798 4276
rect 8772 4168 10640 4196
rect 10704 4168 11100 4196
rect 10060 4140 10088 4168
rect 5169 4131 5227 4137
rect 5169 4097 5181 4131
rect 5215 4128 5227 4131
rect 5442 4128 5448 4140
rect 5215 4100 5448 4128
rect 5215 4097 5227 4100
rect 5169 4091 5227 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 6457 4131 6515 4137
rect 6457 4097 6469 4131
rect 6503 4128 6515 4131
rect 6503 4100 7328 4128
rect 6503 4097 6515 4100
rect 6457 4091 6515 4097
rect 4157 4081 4215 4087
rect 3007 4032 4016 4060
rect 3007 4029 3019 4032
rect 2961 4023 3019 4029
rect 2271 3995 2329 4001
rect 2271 3961 2283 3995
rect 2317 3992 2329 3995
rect 6825 3995 6883 4001
rect 2317 3964 2912 3992
rect 2317 3961 2329 3964
rect 2271 3955 2329 3961
rect 2685 3927 2743 3933
rect 2685 3893 2697 3927
rect 2731 3924 2743 3927
rect 2774 3924 2780 3936
rect 2731 3896 2780 3924
rect 2731 3893 2743 3896
rect 2685 3887 2743 3893
rect 2774 3884 2780 3896
rect 2832 3884 2838 3936
rect 2884 3924 2912 3964
rect 6825 3961 6837 3995
rect 6871 3992 6883 3995
rect 6914 3992 6920 4004
rect 6871 3964 6920 3992
rect 6871 3961 6883 3964
rect 6825 3955 6883 3961
rect 6914 3952 6920 3964
rect 6972 3952 6978 4004
rect 7300 4001 7328 4100
rect 7650 4088 7656 4140
rect 7708 4128 7714 4140
rect 7745 4131 7803 4137
rect 7745 4128 7757 4131
rect 7708 4100 7757 4128
rect 7708 4088 7714 4100
rect 7745 4097 7757 4100
rect 7791 4097 7803 4131
rect 7745 4091 7803 4097
rect 8570 4088 8576 4140
rect 8628 4128 8634 4140
rect 9125 4131 9183 4137
rect 8628 4100 8673 4128
rect 8628 4088 8634 4100
rect 9125 4097 9137 4131
rect 9171 4128 9183 4131
rect 9171 4100 9720 4128
rect 9171 4097 9183 4100
rect 9125 4091 9183 4097
rect 7558 4020 7564 4072
rect 7616 4060 7622 4072
rect 7837 4063 7895 4069
rect 7837 4060 7849 4063
rect 7616 4032 7849 4060
rect 7616 4020 7622 4032
rect 7837 4029 7849 4032
rect 7883 4029 7895 4063
rect 7837 4023 7895 4029
rect 8757 4063 8815 4069
rect 8757 4029 8769 4063
rect 8803 4029 8815 4063
rect 8757 4023 8815 4029
rect 7285 3995 7343 4001
rect 7285 3961 7297 3995
rect 7331 3961 7343 3995
rect 7285 3955 7343 3961
rect 3510 3924 3516 3936
rect 2884 3896 3516 3924
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 3697 3927 3755 3933
rect 3697 3893 3709 3927
rect 3743 3924 3755 3927
rect 4249 3927 4307 3933
rect 4249 3924 4261 3927
rect 3743 3896 4261 3924
rect 3743 3893 3755 3896
rect 3697 3887 3755 3893
rect 4249 3893 4261 3896
rect 4295 3924 4307 3927
rect 4614 3924 4620 3936
rect 4295 3896 4620 3924
rect 4295 3893 4307 3896
rect 4249 3887 4307 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4982 3924 4988 3936
rect 4943 3896 4988 3924
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 8772 3924 8800 4023
rect 9692 4001 9720 4100
rect 10042 4088 10048 4140
rect 10100 4088 10106 4140
rect 10704 4128 10732 4168
rect 10244 4100 10732 4128
rect 9766 4020 9772 4072
rect 9824 4060 9830 4072
rect 10244 4069 10272 4100
rect 10778 4088 10784 4140
rect 10836 4128 10842 4140
rect 10873 4131 10931 4137
rect 10873 4128 10885 4131
rect 10836 4100 10885 4128
rect 10836 4088 10842 4100
rect 10873 4097 10885 4100
rect 10919 4097 10931 4131
rect 11072 4128 11100 4168
rect 11238 4156 11244 4208
rect 11296 4196 11302 4208
rect 12158 4196 12164 4208
rect 11296 4168 12164 4196
rect 11296 4156 11302 4168
rect 12158 4156 12164 4168
rect 12216 4196 12222 4208
rect 12216 4168 12480 4196
rect 12216 4156 12222 4168
rect 11422 4128 11428 4140
rect 11072 4100 11428 4128
rect 10873 4091 10931 4097
rect 11422 4088 11428 4100
rect 11480 4137 11486 4140
rect 11480 4131 11539 4137
rect 11480 4097 11493 4131
rect 11527 4097 11539 4131
rect 11606 4128 11612 4140
rect 11567 4100 11612 4128
rect 11480 4091 11539 4097
rect 11480 4088 11486 4091
rect 11606 4088 11612 4100
rect 11664 4088 11670 4140
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 10137 4063 10195 4069
rect 10137 4060 10149 4063
rect 9824 4032 10149 4060
rect 9824 4020 9830 4032
rect 10137 4029 10149 4032
rect 10183 4029 10195 4063
rect 10137 4023 10195 4029
rect 10229 4063 10287 4069
rect 10229 4029 10241 4063
rect 10275 4029 10287 4063
rect 10962 4060 10968 4072
rect 10923 4032 10968 4060
rect 10229 4023 10287 4029
rect 9677 3995 9735 4001
rect 9677 3961 9689 3995
rect 9723 3961 9735 3995
rect 9677 3955 9735 3961
rect 9950 3952 9956 4004
rect 10008 3992 10014 4004
rect 10244 3992 10272 4023
rect 10962 4020 10968 4032
rect 11020 4020 11026 4072
rect 11057 4063 11115 4069
rect 11057 4029 11069 4063
rect 11103 4029 11115 4063
rect 11716 4060 11744 4091
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 12069 4131 12127 4137
rect 12069 4128 12081 4131
rect 11848 4100 12081 4128
rect 11848 4088 11854 4100
rect 12069 4097 12081 4100
rect 12115 4097 12127 4131
rect 12250 4128 12256 4140
rect 12211 4100 12256 4128
rect 12069 4091 12127 4097
rect 12250 4088 12256 4100
rect 12308 4088 12314 4140
rect 12452 4128 12480 4168
rect 13170 4156 13176 4208
rect 13228 4156 13234 4208
rect 14550 4196 14556 4208
rect 14511 4168 14556 4196
rect 14550 4156 14556 4168
rect 14608 4196 14614 4208
rect 14608 4168 15042 4196
rect 14608 4156 14614 4168
rect 18233 4131 18291 4137
rect 12452 4100 12940 4128
rect 12268 4060 12296 4088
rect 12452 4069 12480 4100
rect 11716 4032 12296 4060
rect 12437 4063 12495 4069
rect 11057 4023 11115 4029
rect 12437 4029 12449 4063
rect 12483 4029 12495 4063
rect 12802 4060 12808 4072
rect 12763 4032 12808 4060
rect 12437 4023 12495 4029
rect 11072 3992 11100 4023
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 12912 4060 12940 4100
rect 18233 4097 18245 4131
rect 18279 4128 18291 4131
rect 18506 4128 18512 4140
rect 18279 4100 18512 4128
rect 18279 4097 18291 4100
rect 18233 4091 18291 4097
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 13814 4060 13820 4072
rect 12912 4032 13820 4060
rect 13814 4020 13820 4032
rect 13872 4020 13878 4072
rect 14737 4063 14795 4069
rect 14737 4029 14749 4063
rect 14783 4060 14795 4063
rect 14826 4060 14832 4072
rect 14783 4032 14832 4060
rect 14783 4029 14795 4032
rect 14737 4023 14795 4029
rect 14826 4020 14832 4032
rect 14884 4020 14890 4072
rect 15470 4020 15476 4072
rect 15528 4060 15534 4072
rect 16485 4063 16543 4069
rect 16485 4060 16497 4063
rect 15528 4032 16497 4060
rect 15528 4020 15534 4032
rect 16485 4029 16497 4032
rect 16531 4029 16543 4063
rect 16485 4023 16543 4029
rect 12161 3995 12219 4001
rect 12161 3992 12173 3995
rect 10008 3964 10272 3992
rect 10980 3964 12173 3992
rect 10008 3952 10014 3964
rect 10980 3924 11008 3964
rect 12161 3961 12173 3964
rect 12207 3961 12219 3995
rect 12161 3955 12219 3961
rect 11882 3924 11888 3936
rect 8772 3896 11008 3924
rect 11843 3896 11888 3924
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 13722 3884 13728 3936
rect 13780 3924 13786 3936
rect 14231 3927 14289 3933
rect 14231 3924 14243 3927
rect 13780 3896 14243 3924
rect 13780 3884 13786 3896
rect 14231 3893 14243 3896
rect 14277 3893 14289 3927
rect 14231 3887 14289 3893
rect 16227 3927 16285 3933
rect 16227 3893 16239 3927
rect 16273 3924 16285 3927
rect 17770 3924 17776 3936
rect 16273 3896 17776 3924
rect 16273 3893 16285 3896
rect 16227 3887 16285 3893
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 18322 3924 18328 3936
rect 18283 3896 18328 3924
rect 18322 3884 18328 3896
rect 18380 3884 18386 3936
rect 0 3834 18860 3856
rect 0 3782 3110 3834
rect 3162 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 3302 3834
rect 3354 3782 3366 3834
rect 3418 3782 6210 3834
rect 6262 3782 6274 3834
rect 6326 3782 6338 3834
rect 6390 3782 6402 3834
rect 6454 3782 6466 3834
rect 6518 3782 9310 3834
rect 9362 3782 9374 3834
rect 9426 3782 9438 3834
rect 9490 3782 9502 3834
rect 9554 3782 9566 3834
rect 9618 3782 12410 3834
rect 12462 3782 12474 3834
rect 12526 3782 12538 3834
rect 12590 3782 12602 3834
rect 12654 3782 12666 3834
rect 12718 3782 15510 3834
rect 15562 3782 15574 3834
rect 15626 3782 15638 3834
rect 15690 3782 15702 3834
rect 15754 3782 15766 3834
rect 15818 3782 18860 3834
rect 0 3760 18860 3782
rect 2774 3680 2780 3732
rect 2832 3720 2838 3732
rect 9950 3720 9956 3732
rect 2832 3692 2877 3720
rect 7576 3692 9956 3720
rect 2832 3680 2838 3692
rect 7576 3664 7604 3692
rect 9950 3680 9956 3692
rect 10008 3680 10014 3732
rect 10045 3723 10103 3729
rect 10045 3689 10057 3723
rect 10091 3720 10103 3723
rect 10962 3720 10968 3732
rect 10091 3692 10968 3720
rect 10091 3689 10103 3692
rect 10045 3683 10103 3689
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 12802 3680 12808 3732
rect 12860 3720 12866 3732
rect 12897 3723 12955 3729
rect 12897 3720 12909 3723
rect 12860 3692 12909 3720
rect 12860 3680 12866 3692
rect 12897 3689 12909 3692
rect 12943 3689 12955 3723
rect 12897 3683 12955 3689
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 18141 3723 18199 3729
rect 18141 3720 18153 3723
rect 14792 3692 18153 3720
rect 14792 3680 14798 3692
rect 18141 3689 18153 3692
rect 18187 3689 18199 3723
rect 18141 3683 18199 3689
rect 2682 3652 2688 3664
rect 2595 3624 2688 3652
rect 2682 3612 2688 3624
rect 2740 3652 2746 3664
rect 4341 3655 4399 3661
rect 4341 3652 4353 3655
rect 2740 3624 4353 3652
rect 2740 3612 2746 3624
rect 4341 3621 4353 3624
rect 4387 3621 4399 3655
rect 4341 3615 4399 3621
rect 5626 3612 5632 3664
rect 5684 3652 5690 3664
rect 7558 3652 7564 3664
rect 5684 3624 7564 3652
rect 5684 3612 5690 3624
rect 2225 3587 2283 3593
rect 2225 3553 2237 3587
rect 2271 3584 2283 3587
rect 3697 3587 3755 3593
rect 3697 3584 3709 3587
rect 2271 3556 3709 3584
rect 2271 3553 2283 3556
rect 2225 3547 2283 3553
rect 3697 3553 3709 3556
rect 3743 3584 3755 3587
rect 3786 3584 3792 3596
rect 3743 3556 3792 3584
rect 3743 3553 3755 3556
rect 3697 3547 3755 3553
rect 3786 3544 3792 3556
rect 3844 3544 3850 3596
rect 4246 3584 4252 3596
rect 3896 3556 4252 3584
rect 1765 3519 1823 3525
rect 1765 3485 1777 3519
rect 1811 3485 1823 3519
rect 1765 3479 1823 3485
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 2590 3516 2596 3528
rect 1903 3488 2596 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 1780 3448 1808 3479
rect 2590 3476 2596 3488
rect 2648 3516 2654 3528
rect 2869 3519 2927 3525
rect 2869 3516 2881 3519
rect 2648 3488 2881 3516
rect 2648 3476 2654 3488
rect 2869 3485 2881 3488
rect 2915 3485 2927 3519
rect 3142 3516 3148 3528
rect 3103 3488 3148 3516
rect 2869 3479 2927 3485
rect 3142 3476 3148 3488
rect 3200 3476 3206 3528
rect 3896 3525 3924 3556
rect 4246 3544 4252 3556
rect 4304 3544 4310 3596
rect 4982 3544 4988 3596
rect 5040 3584 5046 3596
rect 6288 3593 6316 3624
rect 7558 3612 7564 3624
rect 7616 3612 7622 3664
rect 7650 3612 7656 3664
rect 7708 3652 7714 3664
rect 11606 3652 11612 3664
rect 7708 3624 11612 3652
rect 7708 3612 7714 3624
rect 6181 3587 6239 3593
rect 6181 3584 6193 3587
rect 5040 3556 6193 3584
rect 5040 3544 5046 3556
rect 6181 3553 6193 3556
rect 6227 3553 6239 3587
rect 6181 3547 6239 3553
rect 6273 3587 6331 3593
rect 6273 3553 6285 3587
rect 6319 3553 6331 3587
rect 6273 3547 6331 3553
rect 6457 3587 6515 3593
rect 6457 3553 6469 3587
rect 6503 3584 6515 3587
rect 6730 3584 6736 3596
rect 6503 3556 6736 3584
rect 6503 3553 6515 3556
rect 6457 3547 6515 3553
rect 6730 3544 6736 3556
rect 6788 3584 6794 3596
rect 9692 3593 9720 3624
rect 11606 3612 11612 3624
rect 11664 3612 11670 3664
rect 14277 3655 14335 3661
rect 14277 3621 14289 3655
rect 14323 3652 14335 3655
rect 14553 3655 14611 3661
rect 14553 3652 14565 3655
rect 14323 3624 14565 3652
rect 14323 3621 14335 3624
rect 14277 3615 14335 3621
rect 14553 3621 14565 3624
rect 14599 3621 14611 3655
rect 14553 3615 14611 3621
rect 14918 3612 14924 3664
rect 14976 3652 14982 3664
rect 15657 3655 15715 3661
rect 15657 3652 15669 3655
rect 14976 3624 15669 3652
rect 14976 3612 14982 3624
rect 15657 3621 15669 3624
rect 15703 3621 15715 3655
rect 15657 3615 15715 3621
rect 9677 3587 9735 3593
rect 6788 3556 8156 3584
rect 6788 3544 6794 3556
rect 3329 3519 3387 3525
rect 3329 3485 3341 3519
rect 3375 3485 3387 3519
rect 3329 3479 3387 3485
rect 3881 3519 3939 3525
rect 3881 3485 3893 3519
rect 3927 3485 3939 3519
rect 3881 3479 3939 3485
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 2314 3448 2320 3460
rect 1780 3420 2320 3448
rect 2314 3408 2320 3420
rect 2372 3408 2378 3460
rect 566 3340 572 3392
rect 624 3380 630 3392
rect 1581 3383 1639 3389
rect 1581 3380 1593 3383
rect 624 3352 1593 3380
rect 624 3340 630 3352
rect 1581 3349 1593 3352
rect 1627 3349 1639 3383
rect 1581 3343 1639 3349
rect 2866 3340 2872 3392
rect 2924 3380 2930 3392
rect 3053 3383 3111 3389
rect 3053 3380 3065 3383
rect 2924 3352 3065 3380
rect 2924 3340 2930 3352
rect 3053 3349 3065 3352
rect 3099 3349 3111 3383
rect 3344 3380 3372 3479
rect 3988 3448 4016 3479
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 4525 3519 4583 3525
rect 4120 3488 4165 3516
rect 4120 3476 4126 3488
rect 4525 3485 4537 3519
rect 4571 3485 4583 3519
rect 4525 3479 4583 3485
rect 4540 3448 4568 3479
rect 4614 3476 4620 3528
rect 4672 3516 4678 3528
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 4672 3488 5733 3516
rect 4672 3476 4678 3488
rect 5721 3485 5733 3488
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 6549 3519 6607 3525
rect 6549 3485 6561 3519
rect 6595 3516 6607 3519
rect 6638 3516 6644 3528
rect 6595 3488 6644 3516
rect 6595 3485 6607 3488
rect 6549 3479 6607 3485
rect 5442 3448 5448 3460
rect 3988 3420 5448 3448
rect 5442 3408 5448 3420
rect 5500 3408 5506 3460
rect 5920 3448 5948 3479
rect 6638 3476 6644 3488
rect 6696 3476 6702 3528
rect 8128 3525 8156 3556
rect 9677 3553 9689 3587
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 11882 3544 11888 3596
rect 11940 3584 11946 3596
rect 12529 3587 12587 3593
rect 12529 3584 12541 3587
rect 11940 3556 12541 3584
rect 11940 3544 11946 3556
rect 12529 3553 12541 3556
rect 12575 3553 12587 3587
rect 12529 3547 12587 3553
rect 13630 3544 13636 3596
rect 13688 3584 13694 3596
rect 13909 3587 13967 3593
rect 13909 3584 13921 3587
rect 13688 3556 13921 3584
rect 13688 3544 13694 3556
rect 13909 3553 13921 3556
rect 13955 3553 13967 3587
rect 13909 3547 13967 3553
rect 14642 3544 14648 3596
rect 14700 3584 14706 3596
rect 15105 3587 15163 3593
rect 15105 3584 15117 3587
rect 14700 3556 15117 3584
rect 14700 3544 14706 3556
rect 15105 3553 15117 3556
rect 15151 3553 15163 3587
rect 15105 3547 15163 3553
rect 7837 3519 7895 3525
rect 7837 3516 7849 3519
rect 7392 3488 7849 3516
rect 7392 3460 7420 3488
rect 7837 3485 7849 3488
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3485 8171 3519
rect 8113 3479 8171 3485
rect 8297 3519 8355 3525
rect 8297 3485 8309 3519
rect 8343 3485 8355 3519
rect 9766 3516 9772 3528
rect 9727 3488 9772 3516
rect 8297 3479 8355 3485
rect 7374 3448 7380 3460
rect 5920 3420 7380 3448
rect 7374 3408 7380 3420
rect 7432 3408 7438 3460
rect 7558 3408 7564 3460
rect 7616 3448 7622 3460
rect 7745 3451 7803 3457
rect 7745 3448 7757 3451
rect 7616 3420 7757 3448
rect 7616 3408 7622 3420
rect 7745 3417 7757 3420
rect 7791 3417 7803 3451
rect 7852 3448 7880 3479
rect 8202 3448 8208 3460
rect 7852 3420 8208 3448
rect 7745 3411 7803 3417
rect 8202 3408 8208 3420
rect 8260 3408 8266 3460
rect 8312 3448 8340 3479
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 12621 3519 12679 3525
rect 12621 3485 12633 3519
rect 12667 3516 12679 3519
rect 13722 3516 13728 3528
rect 12667 3488 13728 3516
rect 12667 3485 12679 3488
rect 12621 3479 12679 3485
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 15013 3519 15071 3525
rect 15013 3516 15025 3519
rect 13872 3488 15025 3516
rect 13872 3476 13878 3488
rect 15013 3485 15025 3488
rect 15059 3516 15071 3519
rect 15286 3516 15292 3528
rect 15059 3488 15292 3516
rect 15059 3485 15071 3488
rect 15013 3479 15071 3485
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 15657 3519 15715 3525
rect 15657 3485 15669 3519
rect 15703 3516 15715 3519
rect 15746 3516 15752 3528
rect 15703 3488 15752 3516
rect 15703 3485 15715 3488
rect 15657 3479 15715 3485
rect 15746 3476 15752 3488
rect 15804 3476 15810 3528
rect 15838 3476 15844 3528
rect 15896 3516 15902 3528
rect 16117 3519 16175 3525
rect 16117 3516 16129 3519
rect 15896 3488 16129 3516
rect 15896 3476 15902 3488
rect 16117 3485 16129 3488
rect 16163 3485 16175 3519
rect 16117 3479 16175 3485
rect 18138 3476 18144 3528
rect 18196 3476 18202 3528
rect 10778 3448 10784 3460
rect 8312 3420 10784 3448
rect 4154 3380 4160 3392
rect 3344 3352 4160 3380
rect 3053 3343 3111 3349
rect 4154 3340 4160 3352
rect 4212 3380 4218 3392
rect 5718 3380 5724 3392
rect 4212 3352 5724 3380
rect 4212 3340 4218 3352
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 5813 3383 5871 3389
rect 5813 3349 5825 3383
rect 5859 3380 5871 3383
rect 5994 3380 6000 3392
rect 5859 3352 6000 3380
rect 5859 3349 5871 3352
rect 5813 3343 5871 3349
rect 5994 3340 6000 3352
rect 6052 3340 6058 3392
rect 6181 3383 6239 3389
rect 6181 3349 6193 3383
rect 6227 3380 6239 3383
rect 6546 3380 6552 3392
rect 6227 3352 6552 3380
rect 6227 3349 6239 3352
rect 6181 3343 6239 3349
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 6638 3340 6644 3392
rect 6696 3380 6702 3392
rect 8312 3380 8340 3420
rect 10778 3408 10784 3420
rect 10836 3408 10842 3460
rect 11422 3408 11428 3460
rect 11480 3448 11486 3460
rect 11974 3448 11980 3460
rect 11480 3420 11980 3448
rect 11480 3408 11486 3420
rect 11974 3408 11980 3420
rect 12032 3448 12038 3460
rect 13630 3448 13636 3460
rect 12032 3420 13636 3448
rect 12032 3408 12038 3420
rect 13630 3408 13636 3420
rect 13688 3408 13694 3460
rect 6696 3352 8340 3380
rect 6696 3340 6702 3352
rect 8386 3340 8392 3392
rect 8444 3380 8450 3392
rect 8573 3383 8631 3389
rect 8573 3380 8585 3383
rect 8444 3352 8585 3380
rect 8444 3340 8450 3352
rect 8573 3349 8585 3352
rect 8619 3380 8631 3383
rect 9030 3380 9036 3392
rect 8619 3352 9036 3380
rect 8619 3349 8631 3352
rect 8573 3343 8631 3349
rect 9030 3340 9036 3352
rect 9088 3340 9094 3392
rect 11330 3340 11336 3392
rect 11388 3380 11394 3392
rect 12253 3383 12311 3389
rect 12253 3380 12265 3383
rect 11388 3352 12265 3380
rect 11388 3340 11394 3352
rect 12253 3349 12265 3352
rect 12299 3380 12311 3383
rect 13170 3380 13176 3392
rect 12299 3352 13176 3380
rect 12299 3349 12311 3352
rect 12253 3343 12311 3349
rect 13170 3340 13176 3352
rect 13228 3340 13234 3392
rect 13740 3380 13768 3476
rect 14921 3451 14979 3457
rect 14921 3448 14933 3451
rect 14016 3420 14933 3448
rect 14016 3380 14044 3420
rect 14921 3417 14933 3420
rect 14967 3417 14979 3451
rect 17865 3451 17923 3457
rect 14921 3411 14979 3417
rect 14366 3380 14372 3392
rect 13740 3352 14044 3380
rect 14327 3352 14372 3380
rect 14366 3340 14372 3352
rect 14424 3340 14430 3392
rect 15102 3340 15108 3392
rect 15160 3380 15166 3392
rect 15473 3383 15531 3389
rect 15473 3380 15485 3383
rect 15160 3352 15485 3380
rect 15160 3340 15166 3352
rect 15473 3349 15485 3352
rect 15519 3380 15531 3383
rect 16500 3380 16528 3434
rect 17865 3417 17877 3451
rect 17911 3448 17923 3451
rect 18156 3448 18184 3476
rect 18233 3451 18291 3457
rect 18233 3448 18245 3451
rect 17911 3420 18245 3448
rect 17911 3417 17923 3420
rect 17865 3411 17923 3417
rect 18233 3417 18245 3420
rect 18279 3417 18291 3451
rect 18233 3411 18291 3417
rect 15519 3352 16528 3380
rect 15519 3349 15531 3352
rect 15473 3343 15531 3349
rect 0 3290 18860 3312
rect 0 3238 4660 3290
rect 4712 3238 4724 3290
rect 4776 3238 4788 3290
rect 4840 3238 4852 3290
rect 4904 3238 4916 3290
rect 4968 3238 7760 3290
rect 7812 3238 7824 3290
rect 7876 3238 7888 3290
rect 7940 3238 7952 3290
rect 8004 3238 8016 3290
rect 8068 3238 10860 3290
rect 10912 3238 10924 3290
rect 10976 3238 10988 3290
rect 11040 3238 11052 3290
rect 11104 3238 11116 3290
rect 11168 3238 13960 3290
rect 14012 3238 14024 3290
rect 14076 3238 14088 3290
rect 14140 3238 14152 3290
rect 14204 3238 14216 3290
rect 14268 3238 17060 3290
rect 17112 3238 17124 3290
rect 17176 3238 17188 3290
rect 17240 3238 17252 3290
rect 17304 3238 17316 3290
rect 17368 3238 18860 3290
rect 0 3216 18860 3238
rect 2041 3179 2099 3185
rect 2041 3145 2053 3179
rect 2087 3145 2099 3179
rect 2590 3176 2596 3188
rect 2551 3148 2596 3176
rect 2041 3139 2099 3145
rect 566 3108 572 3120
rect 527 3080 572 3108
rect 566 3068 572 3080
rect 624 3068 630 3120
rect 2056 3108 2084 3139
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 3142 3176 3148 3188
rect 3103 3148 3148 3176
rect 3142 3136 3148 3148
rect 3200 3136 3206 3188
rect 4062 3176 4068 3188
rect 3252 3148 4068 3176
rect 2314 3108 2320 3120
rect 2056 3080 2320 3108
rect 2314 3068 2320 3080
rect 2372 3108 2378 3120
rect 3252 3108 3280 3148
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 5442 3176 5448 3188
rect 5403 3148 5448 3176
rect 5442 3136 5448 3148
rect 5500 3136 5506 3188
rect 5718 3136 5724 3188
rect 5776 3176 5782 3188
rect 5905 3179 5963 3185
rect 5905 3176 5917 3179
rect 5776 3148 5917 3176
rect 5776 3136 5782 3148
rect 5905 3145 5917 3148
rect 5951 3145 5963 3179
rect 5905 3139 5963 3145
rect 9030 3136 9036 3188
rect 9088 3176 9094 3188
rect 11330 3176 11336 3188
rect 9088 3148 11336 3176
rect 9088 3136 9094 3148
rect 4525 3111 4583 3117
rect 4525 3108 4537 3111
rect 2372 3080 3280 3108
rect 2372 3068 2378 3080
rect 2682 3040 2688 3052
rect 1702 3012 2268 3040
rect 2643 3012 2688 3040
rect 290 2972 296 2984
rect 251 2944 296 2972
rect 290 2932 296 2944
rect 348 2932 354 2984
rect 2240 2845 2268 3012
rect 2682 3000 2688 3012
rect 2740 3000 2746 3052
rect 3252 3049 3280 3080
rect 3712 3080 4537 3108
rect 3712 3052 3740 3080
rect 4525 3077 4537 3080
rect 4571 3077 4583 3111
rect 6546 3108 6552 3120
rect 4525 3071 4583 3077
rect 4632 3080 6552 3108
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 3694 3040 3700 3052
rect 3607 3012 3700 3040
rect 3237 3003 3295 3009
rect 3068 2972 3096 3003
rect 3694 3000 3700 3012
rect 3752 3000 3758 3052
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3040 3939 3043
rect 3973 3043 4031 3049
rect 3973 3040 3985 3043
rect 3927 3012 3985 3040
rect 3927 3009 3939 3012
rect 3881 3003 3939 3009
rect 3973 3009 3985 3012
rect 4019 3009 4031 3043
rect 4154 3040 4160 3052
rect 4115 3012 4160 3040
rect 3973 3003 4031 3009
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 4246 3000 4252 3052
rect 4304 3040 4310 3052
rect 4632 3049 4660 3080
rect 6546 3068 6552 3080
rect 6604 3068 6610 3120
rect 7098 3068 7104 3120
rect 7156 3108 7162 3120
rect 7377 3111 7435 3117
rect 7377 3108 7389 3111
rect 7156 3080 7389 3108
rect 7156 3068 7162 3080
rect 7377 3077 7389 3080
rect 7423 3077 7435 3111
rect 7377 3071 7435 3077
rect 7561 3111 7619 3117
rect 7561 3077 7573 3111
rect 7607 3108 7619 3111
rect 7929 3111 7987 3117
rect 7929 3108 7941 3111
rect 7607 3080 7941 3108
rect 7607 3077 7619 3080
rect 7561 3071 7619 3077
rect 7929 3077 7941 3080
rect 7975 3108 7987 3111
rect 9214 3108 9220 3120
rect 7975 3080 9220 3108
rect 7975 3077 7987 3080
rect 7929 3071 7987 3077
rect 9214 3068 9220 3080
rect 9272 3068 9278 3120
rect 9858 3068 9864 3120
rect 9916 3108 9922 3120
rect 9916 3080 10088 3108
rect 10796 3094 10824 3148
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 12986 3176 12992 3188
rect 11532 3148 12992 3176
rect 9916 3068 9922 3080
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 4304 3012 4445 3040
rect 4304 3000 4310 3012
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 4433 3003 4491 3009
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 7282 3040 7288 3052
rect 5859 3012 7288 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 3510 2972 3516 2984
rect 3068 2944 3516 2972
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 4448 2904 4476 3003
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 7650 3040 7656 3052
rect 7611 3012 7656 3040
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 8202 3040 8208 3052
rect 7800 3012 7845 3040
rect 8163 3012 8208 3040
rect 7800 3000 7806 3012
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 10060 3049 10088 3080
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3009 10011 3043
rect 9953 3003 10011 3009
rect 10045 3043 10103 3049
rect 10045 3009 10057 3043
rect 10091 3009 10103 3043
rect 10045 3003 10103 3009
rect 5994 2932 6000 2984
rect 6052 2972 6058 2984
rect 6273 2975 6331 2981
rect 6273 2972 6285 2975
rect 6052 2944 6285 2972
rect 6052 2932 6058 2944
rect 6273 2941 6285 2944
rect 6319 2941 6331 2975
rect 6273 2935 6331 2941
rect 7466 2932 7472 2984
rect 7524 2972 7530 2984
rect 9861 2975 9919 2981
rect 9861 2972 9873 2975
rect 7524 2944 9873 2972
rect 7524 2932 7530 2944
rect 9861 2941 9873 2944
rect 9907 2941 9919 2975
rect 9968 2972 9996 3003
rect 10413 2975 10471 2981
rect 9968 2944 10088 2972
rect 9861 2935 9919 2941
rect 7098 2904 7104 2916
rect 4448 2876 7104 2904
rect 7098 2864 7104 2876
rect 7156 2864 7162 2916
rect 8389 2907 8447 2913
rect 8389 2873 8401 2907
rect 8435 2904 8447 2907
rect 9122 2904 9128 2916
rect 8435 2876 9128 2904
rect 8435 2873 8447 2876
rect 8389 2867 8447 2873
rect 9122 2864 9128 2876
rect 9180 2864 9186 2916
rect 2225 2839 2283 2845
rect 2225 2805 2237 2839
rect 2271 2836 2283 2839
rect 2498 2836 2504 2848
rect 2271 2808 2504 2836
rect 2271 2805 2283 2808
rect 2225 2799 2283 2805
rect 2498 2796 2504 2808
rect 2556 2796 2562 2848
rect 3786 2836 3792 2848
rect 3747 2808 3792 2836
rect 3786 2796 3792 2808
rect 3844 2796 3850 2848
rect 3973 2839 4031 2845
rect 3973 2805 3985 2839
rect 4019 2836 4031 2839
rect 4338 2836 4344 2848
rect 4019 2808 4344 2836
rect 4019 2805 4031 2808
rect 3973 2799 4031 2805
rect 4338 2796 4344 2808
rect 4396 2796 4402 2848
rect 6733 2839 6791 2845
rect 6733 2805 6745 2839
rect 6779 2836 6791 2839
rect 7190 2836 7196 2848
rect 6779 2808 7196 2836
rect 6779 2805 6791 2808
rect 6733 2799 6791 2805
rect 7190 2796 7196 2808
rect 7248 2796 7254 2848
rect 7837 2839 7895 2845
rect 7837 2805 7849 2839
rect 7883 2836 7895 2839
rect 8846 2836 8852 2848
rect 7883 2808 8852 2836
rect 7883 2805 7895 2808
rect 7837 2799 7895 2805
rect 8846 2796 8852 2808
rect 8904 2796 8910 2848
rect 9030 2796 9036 2848
rect 9088 2836 9094 2848
rect 9401 2839 9459 2845
rect 9401 2836 9413 2839
rect 9088 2808 9413 2836
rect 9088 2796 9094 2808
rect 9401 2805 9413 2808
rect 9447 2805 9459 2839
rect 10060 2836 10088 2944
rect 10413 2941 10425 2975
rect 10459 2972 10471 2975
rect 11532 2972 11560 3148
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 14642 3176 14648 3188
rect 14603 3148 14648 3176
rect 14642 3136 14648 3148
rect 14700 3136 14706 3188
rect 14875 3179 14933 3185
rect 14875 3145 14887 3179
rect 14921 3176 14933 3179
rect 15838 3176 15844 3188
rect 14921 3148 15844 3176
rect 14921 3145 14933 3148
rect 14875 3139 14933 3145
rect 15838 3136 15844 3148
rect 15896 3136 15902 3188
rect 15102 3068 15108 3120
rect 15160 3108 15166 3120
rect 15160 3094 15318 3108
rect 15160 3080 15332 3094
rect 15160 3068 15166 3080
rect 11839 3043 11897 3049
rect 11839 3009 11851 3043
rect 11885 3040 11897 3043
rect 12437 3043 12495 3049
rect 12437 3040 12449 3043
rect 11885 3012 12449 3040
rect 11885 3009 11897 3012
rect 11839 3003 11897 3009
rect 12437 3009 12449 3012
rect 12483 3040 12495 3043
rect 12802 3040 12808 3052
rect 12483 3012 12808 3040
rect 12483 3009 12495 3012
rect 12437 3003 12495 3009
rect 12802 3000 12808 3012
rect 12860 3000 12866 3052
rect 13538 3040 13544 3052
rect 13499 3012 13544 3040
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 14277 3043 14335 3049
rect 14277 3009 14289 3043
rect 14323 3040 14335 3043
rect 14366 3040 14372 3052
rect 14323 3012 14372 3040
rect 14323 3009 14335 3012
rect 14277 3003 14335 3009
rect 10459 2944 11560 2972
rect 12345 2975 12403 2981
rect 10459 2941 10471 2944
rect 10413 2935 10471 2941
rect 12345 2941 12357 2975
rect 12391 2941 12403 2975
rect 12345 2935 12403 2941
rect 10318 2836 10324 2848
rect 10060 2808 10324 2836
rect 9401 2799 9459 2805
rect 10318 2796 10324 2808
rect 10376 2836 10382 2848
rect 12360 2836 12388 2935
rect 12805 2907 12863 2913
rect 12805 2873 12817 2907
rect 12851 2904 12863 2907
rect 13740 2904 13768 3003
rect 14366 3000 14372 3012
rect 14424 3000 14430 3052
rect 14550 3040 14556 3052
rect 14511 3012 14556 3040
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 14734 3040 14740 3052
rect 14695 3012 14740 3040
rect 14734 3000 14740 3012
rect 14792 3040 14798 3052
rect 15304 3040 15332 3080
rect 15378 3040 15384 3052
rect 14792 3012 15148 3040
rect 15304 3012 15384 3040
rect 14792 3000 14798 3012
rect 15120 2984 15148 3012
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 16301 3043 16359 3049
rect 16301 3009 16313 3043
rect 16347 3040 16359 3043
rect 18322 3040 18328 3052
rect 16347 3012 18328 3040
rect 16347 3009 16359 3012
rect 16301 3003 16359 3009
rect 18322 3000 18328 3012
rect 18380 3000 18386 3052
rect 14093 2975 14151 2981
rect 14093 2941 14105 2975
rect 14139 2972 14151 2975
rect 14918 2972 14924 2984
rect 14139 2944 14924 2972
rect 14139 2941 14151 2944
rect 14093 2935 14151 2941
rect 14918 2932 14924 2944
rect 14976 2932 14982 2984
rect 15102 2932 15108 2984
rect 15160 2932 15166 2984
rect 15838 2932 15844 2984
rect 15896 2972 15902 2984
rect 16669 2975 16727 2981
rect 16669 2972 16681 2975
rect 15896 2944 16681 2972
rect 15896 2932 15902 2944
rect 16669 2941 16681 2944
rect 16715 2972 16727 2975
rect 17862 2972 17868 2984
rect 16715 2944 17868 2972
rect 16715 2941 16727 2944
rect 16669 2935 16727 2941
rect 17862 2932 17868 2944
rect 17920 2932 17926 2984
rect 12851 2876 13768 2904
rect 12851 2873 12863 2876
rect 12805 2867 12863 2873
rect 10376 2808 12388 2836
rect 10376 2796 10382 2808
rect 0 2746 18860 2768
rect 0 2694 3110 2746
rect 3162 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 3302 2746
rect 3354 2694 3366 2746
rect 3418 2694 6210 2746
rect 6262 2694 6274 2746
rect 6326 2694 6338 2746
rect 6390 2694 6402 2746
rect 6454 2694 6466 2746
rect 6518 2694 9310 2746
rect 9362 2694 9374 2746
rect 9426 2694 9438 2746
rect 9490 2694 9502 2746
rect 9554 2694 9566 2746
rect 9618 2694 12410 2746
rect 12462 2694 12474 2746
rect 12526 2694 12538 2746
rect 12590 2694 12602 2746
rect 12654 2694 12666 2746
rect 12718 2694 15510 2746
rect 15562 2694 15574 2746
rect 15626 2694 15638 2746
rect 15690 2694 15702 2746
rect 15754 2694 15766 2746
rect 15818 2694 18860 2746
rect 0 2672 18860 2694
rect 3237 2635 3295 2641
rect 3237 2601 3249 2635
rect 3283 2632 3295 2635
rect 3510 2632 3516 2644
rect 3283 2604 3516 2632
rect 3283 2601 3295 2604
rect 3237 2595 3295 2601
rect 3510 2592 3516 2604
rect 3568 2632 3574 2644
rect 6733 2635 6791 2641
rect 3568 2604 4016 2632
rect 3568 2592 3574 2604
rect 3786 2564 3792 2576
rect 3068 2536 3792 2564
rect 3068 2505 3096 2536
rect 3786 2524 3792 2536
rect 3844 2524 3850 2576
rect 3053 2499 3111 2505
rect 3053 2465 3065 2499
rect 3099 2465 3111 2499
rect 3694 2496 3700 2508
rect 3655 2468 3700 2496
rect 3053 2459 3111 2465
rect 3694 2456 3700 2468
rect 3752 2456 3758 2508
rect 3988 2505 4016 2604
rect 6733 2601 6745 2635
rect 6779 2632 6791 2635
rect 7466 2632 7472 2644
rect 6779 2604 7472 2632
rect 6779 2601 6791 2604
rect 6733 2595 6791 2601
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 7561 2635 7619 2641
rect 7561 2601 7573 2635
rect 7607 2632 7619 2635
rect 7650 2632 7656 2644
rect 7607 2604 7656 2632
rect 7607 2601 7619 2604
rect 7561 2595 7619 2601
rect 7650 2592 7656 2604
rect 7708 2592 7714 2644
rect 10318 2641 10324 2644
rect 10275 2635 10324 2641
rect 10275 2601 10287 2635
rect 10321 2601 10324 2635
rect 10275 2595 10324 2601
rect 10318 2592 10324 2595
rect 10376 2592 10382 2644
rect 14550 2632 14556 2644
rect 11348 2604 14556 2632
rect 6457 2567 6515 2573
rect 6457 2533 6469 2567
rect 6503 2564 6515 2567
rect 7742 2564 7748 2576
rect 6503 2536 7748 2564
rect 6503 2533 6515 2536
rect 6457 2527 6515 2533
rect 7742 2524 7748 2536
rect 7800 2524 7806 2576
rect 3973 2499 4031 2505
rect 3973 2465 3985 2499
rect 4019 2465 4031 2499
rect 3973 2459 4031 2465
rect 4801 2499 4859 2505
rect 4801 2465 4813 2499
rect 4847 2496 4859 2499
rect 5442 2496 5448 2508
rect 4847 2468 5448 2496
rect 4847 2465 4859 2468
rect 4801 2459 4859 2465
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 7006 2456 7012 2508
rect 7064 2496 7070 2508
rect 8846 2496 8852 2508
rect 7064 2468 8156 2496
rect 8807 2468 8852 2496
rect 7064 2456 7070 2468
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2428 3387 2431
rect 3375 2400 3832 2428
rect 3375 2397 3387 2400
rect 3329 2391 3387 2397
rect 3804 2304 3832 2400
rect 5534 2388 5540 2440
rect 5592 2428 5598 2440
rect 6273 2431 6331 2437
rect 6273 2428 6285 2431
rect 5592 2400 6285 2428
rect 5592 2388 5598 2400
rect 6273 2397 6285 2400
rect 6319 2397 6331 2431
rect 6273 2391 6331 2397
rect 6457 2431 6515 2437
rect 6457 2397 6469 2431
rect 6503 2428 6515 2431
rect 6546 2428 6552 2440
rect 6503 2400 6552 2428
rect 6503 2397 6515 2400
rect 6457 2391 6515 2397
rect 6546 2388 6552 2400
rect 6604 2388 6610 2440
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2397 6975 2431
rect 7098 2428 7104 2440
rect 7059 2400 7104 2428
rect 6917 2391 6975 2397
rect 4893 2363 4951 2369
rect 4893 2329 4905 2363
rect 4939 2360 4951 2363
rect 5626 2360 5632 2372
rect 4939 2332 5632 2360
rect 4939 2329 4951 2332
rect 4893 2323 4951 2329
rect 5626 2320 5632 2332
rect 5684 2320 5690 2372
rect 6822 2360 6828 2372
rect 6783 2332 6828 2360
rect 6822 2320 6828 2332
rect 6880 2320 6886 2372
rect 842 2252 848 2304
rect 900 2292 906 2304
rect 3053 2295 3111 2301
rect 3053 2292 3065 2295
rect 900 2264 3065 2292
rect 900 2252 906 2264
rect 3053 2261 3065 2264
rect 3099 2261 3111 2295
rect 3053 2255 3111 2261
rect 3786 2252 3792 2304
rect 3844 2292 3850 2304
rect 4985 2295 5043 2301
rect 4985 2292 4997 2295
rect 3844 2264 4997 2292
rect 3844 2252 3850 2264
rect 4985 2261 4997 2264
rect 5031 2261 5043 2295
rect 4985 2255 5043 2261
rect 5258 2252 5264 2304
rect 5316 2292 5322 2304
rect 5353 2295 5411 2301
rect 5353 2292 5365 2295
rect 5316 2264 5365 2292
rect 5316 2252 5322 2264
rect 5353 2261 5365 2264
rect 5399 2261 5411 2295
rect 6932 2292 6960 2391
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 8128 2437 8156 2468
rect 8846 2456 8852 2468
rect 8904 2456 8910 2508
rect 9122 2496 9128 2508
rect 8956 2468 9128 2496
rect 8956 2440 8984 2468
rect 9122 2456 9128 2468
rect 9180 2456 9186 2508
rect 7561 2431 7619 2437
rect 7561 2428 7573 2431
rect 7248 2400 7573 2428
rect 7248 2388 7254 2400
rect 7561 2397 7573 2400
rect 7607 2397 7619 2431
rect 7561 2391 7619 2397
rect 8113 2431 8171 2437
rect 8113 2397 8125 2431
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2428 8263 2431
rect 8481 2431 8539 2437
rect 8481 2428 8493 2431
rect 8251 2400 8493 2428
rect 8251 2397 8263 2400
rect 8205 2391 8263 2397
rect 8481 2397 8493 2400
rect 8527 2397 8539 2431
rect 8481 2391 8539 2397
rect 8938 2388 8944 2440
rect 8996 2388 9002 2440
rect 7006 2320 7012 2372
rect 7064 2360 7070 2372
rect 7285 2363 7343 2369
rect 7285 2360 7297 2363
rect 7064 2332 7297 2360
rect 7064 2320 7070 2332
rect 7285 2329 7297 2332
rect 7331 2329 7343 2363
rect 7466 2360 7472 2372
rect 7427 2332 7472 2360
rect 7285 2323 7343 2329
rect 7466 2320 7472 2332
rect 7524 2320 7530 2372
rect 9214 2320 9220 2372
rect 9272 2320 9278 2372
rect 10594 2320 10600 2372
rect 10652 2360 10658 2372
rect 10778 2360 10784 2372
rect 10652 2332 10784 2360
rect 10652 2320 10658 2332
rect 10778 2320 10784 2332
rect 10836 2360 10842 2372
rect 11348 2369 11376 2604
rect 14550 2592 14556 2604
rect 14608 2632 14614 2644
rect 15194 2632 15200 2644
rect 14608 2604 15200 2632
rect 14608 2592 14614 2604
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 11882 2524 11888 2576
rect 11940 2564 11946 2576
rect 12894 2564 12900 2576
rect 11940 2536 12900 2564
rect 11940 2524 11946 2536
rect 12894 2524 12900 2536
rect 12952 2524 12958 2576
rect 12986 2524 12992 2576
rect 13044 2564 13050 2576
rect 13044 2536 13089 2564
rect 13044 2524 13050 2536
rect 11514 2496 11520 2508
rect 11475 2468 11520 2496
rect 11514 2456 11520 2468
rect 11572 2456 11578 2508
rect 12250 2456 12256 2508
rect 12308 2496 12314 2508
rect 13265 2499 13323 2505
rect 13265 2496 13277 2499
rect 12308 2468 12480 2496
rect 12308 2456 12314 2468
rect 12342 2428 12348 2440
rect 12303 2400 12348 2428
rect 12342 2388 12348 2400
rect 12400 2388 12406 2440
rect 12452 2437 12480 2468
rect 12544 2468 13277 2496
rect 12544 2437 12572 2468
rect 13265 2465 13277 2468
rect 13311 2465 13323 2499
rect 13814 2496 13820 2508
rect 13775 2468 13820 2496
rect 13265 2459 13323 2465
rect 13814 2456 13820 2468
rect 13872 2456 13878 2508
rect 15841 2499 15899 2505
rect 15841 2465 15853 2499
rect 15887 2496 15899 2499
rect 16942 2496 16948 2508
rect 15887 2468 16948 2496
rect 15887 2465 15899 2468
rect 15841 2459 15899 2465
rect 16942 2456 16948 2468
rect 17000 2456 17006 2508
rect 17862 2496 17868 2508
rect 17823 2468 17868 2496
rect 17862 2456 17868 2468
rect 17920 2456 17926 2508
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2397 12495 2431
rect 12437 2391 12495 2397
rect 12529 2431 12587 2437
rect 12529 2397 12541 2431
rect 12575 2428 12587 2431
rect 12618 2428 12624 2440
rect 12575 2400 12624 2428
rect 12575 2397 12587 2400
rect 12529 2391 12587 2397
rect 12618 2388 12624 2400
rect 12676 2388 12682 2440
rect 12713 2431 12771 2437
rect 12713 2397 12725 2431
rect 12759 2428 12771 2431
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 12759 2400 12817 2428
rect 12759 2397 12771 2400
rect 12713 2391 12771 2397
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 13541 2431 13599 2437
rect 13541 2428 13553 2431
rect 12805 2391 12863 2397
rect 13004 2400 13553 2428
rect 11333 2363 11391 2369
rect 11333 2360 11345 2363
rect 10836 2332 11345 2360
rect 10836 2320 10842 2332
rect 11333 2329 11345 2332
rect 11379 2329 11391 2363
rect 11333 2323 11391 2329
rect 11606 2320 11612 2372
rect 11664 2360 11670 2372
rect 12897 2363 12955 2369
rect 12897 2360 12909 2363
rect 11664 2332 12909 2360
rect 11664 2320 11670 2332
rect 12897 2329 12909 2332
rect 12943 2329 12955 2363
rect 12897 2323 12955 2329
rect 7374 2292 7380 2304
rect 6932 2264 7380 2292
rect 5353 2255 5411 2261
rect 7374 2252 7380 2264
rect 7432 2252 7438 2304
rect 7650 2252 7656 2304
rect 7708 2292 7714 2304
rect 7929 2295 7987 2301
rect 7929 2292 7941 2295
rect 7708 2264 7941 2292
rect 7708 2252 7714 2264
rect 7929 2261 7941 2264
rect 7975 2261 7987 2295
rect 7929 2255 7987 2261
rect 8754 2252 8760 2304
rect 8812 2292 8818 2304
rect 10873 2295 10931 2301
rect 10873 2292 10885 2295
rect 8812 2264 10885 2292
rect 8812 2252 8818 2264
rect 10873 2261 10885 2264
rect 10919 2261 10931 2295
rect 11238 2292 11244 2304
rect 11199 2264 11244 2292
rect 10873 2255 10931 2261
rect 11238 2252 11244 2264
rect 11296 2252 11302 2304
rect 11974 2252 11980 2304
rect 12032 2292 12038 2304
rect 12342 2292 12348 2304
rect 12032 2264 12348 2292
rect 12032 2252 12038 2264
rect 12342 2252 12348 2264
rect 12400 2292 12406 2304
rect 13004 2292 13032 2400
rect 13541 2397 13553 2400
rect 13587 2397 13599 2431
rect 13541 2391 13599 2397
rect 13630 2388 13636 2440
rect 13688 2437 13694 2440
rect 13688 2431 13737 2437
rect 13688 2397 13691 2431
rect 13725 2397 13737 2431
rect 13688 2391 13737 2397
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2428 18291 2431
rect 18506 2428 18512 2440
rect 18279 2400 18512 2428
rect 18279 2397 18291 2400
rect 18233 2391 18291 2397
rect 13688 2388 13694 2391
rect 18506 2388 18512 2400
rect 18564 2388 18570 2440
rect 13081 2363 13139 2369
rect 13081 2329 13093 2363
rect 13127 2329 13139 2363
rect 13081 2323 13139 2329
rect 12400 2264 13032 2292
rect 13096 2292 13124 2323
rect 13170 2320 13176 2372
rect 13228 2360 13234 2372
rect 13648 2360 13676 2388
rect 13228 2332 13676 2360
rect 14084 2363 14142 2369
rect 13228 2320 13234 2332
rect 14084 2329 14096 2363
rect 14130 2360 14142 2363
rect 14550 2360 14556 2372
rect 14130 2332 14556 2360
rect 14130 2329 14142 2332
rect 14084 2323 14142 2329
rect 14550 2320 14556 2332
rect 14608 2320 14614 2372
rect 17586 2360 17592 2372
rect 15672 2332 16422 2360
rect 17547 2332 17592 2360
rect 13449 2295 13507 2301
rect 13449 2292 13461 2295
rect 13096 2264 13461 2292
rect 12400 2252 12406 2264
rect 13449 2261 13461 2264
rect 13495 2261 13507 2295
rect 13449 2255 13507 2261
rect 14642 2252 14648 2304
rect 14700 2292 14706 2304
rect 15197 2295 15255 2301
rect 15197 2292 15209 2295
rect 14700 2264 15209 2292
rect 14700 2252 14706 2264
rect 15197 2261 15209 2264
rect 15243 2261 15255 2295
rect 15378 2292 15384 2304
rect 15339 2264 15384 2292
rect 15197 2255 15255 2261
rect 15378 2252 15384 2264
rect 15436 2292 15442 2304
rect 15672 2301 15700 2332
rect 17586 2320 17592 2332
rect 17644 2320 17650 2372
rect 15657 2295 15715 2301
rect 15657 2292 15669 2295
rect 15436 2264 15669 2292
rect 15436 2252 15442 2264
rect 15657 2261 15669 2264
rect 15703 2261 15715 2295
rect 15657 2255 15715 2261
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 16172 2264 18337 2292
rect 16172 2252 16178 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 0 2202 18860 2224
rect 0 2150 4660 2202
rect 4712 2150 4724 2202
rect 4776 2150 4788 2202
rect 4840 2150 4852 2202
rect 4904 2150 4916 2202
rect 4968 2150 7760 2202
rect 7812 2150 7824 2202
rect 7876 2150 7888 2202
rect 7940 2150 7952 2202
rect 8004 2150 8016 2202
rect 8068 2150 10860 2202
rect 10912 2150 10924 2202
rect 10976 2150 10988 2202
rect 11040 2150 11052 2202
rect 11104 2150 11116 2202
rect 11168 2150 13960 2202
rect 14012 2150 14024 2202
rect 14076 2150 14088 2202
rect 14140 2150 14152 2202
rect 14204 2150 14216 2202
rect 14268 2150 17060 2202
rect 17112 2150 17124 2202
rect 17176 2150 17188 2202
rect 17240 2150 17252 2202
rect 17304 2150 17316 2202
rect 17368 2150 18860 2202
rect 0 2128 18860 2150
rect 1210 2048 1216 2100
rect 1268 2088 1274 2100
rect 2958 2088 2964 2100
rect 1268 2060 2964 2088
rect 1268 2048 1274 2060
rect 2958 2048 2964 2060
rect 3016 2088 3022 2100
rect 3786 2088 3792 2100
rect 3016 2060 3372 2088
rect 3747 2060 3792 2088
rect 3016 2048 3022 2060
rect 842 2020 848 2032
rect 803 1992 848 2020
rect 842 1980 848 1992
rect 900 1980 906 2032
rect 2774 2020 2780 2032
rect 2332 1992 2780 2020
rect 290 1844 296 1896
rect 348 1884 354 1896
rect 569 1887 627 1893
rect 569 1884 581 1887
rect 348 1856 581 1884
rect 348 1844 354 1856
rect 569 1853 581 1856
rect 615 1884 627 1887
rect 1210 1884 1216 1896
rect 615 1856 1216 1884
rect 615 1853 627 1856
rect 569 1847 627 1853
rect 1210 1844 1216 1856
rect 1268 1844 1274 1896
rect 1964 1816 1992 1938
rect 2332 1893 2360 1992
rect 2774 1980 2780 1992
rect 2832 1980 2838 2032
rect 2958 1912 2964 1964
rect 3016 1952 3022 1964
rect 3344 1961 3372 2060
rect 3786 2048 3792 2060
rect 3844 2048 3850 2100
rect 4338 2048 4344 2100
rect 4396 2088 4402 2100
rect 4893 2091 4951 2097
rect 4893 2088 4905 2091
rect 4396 2060 4905 2088
rect 4396 2048 4402 2060
rect 4893 2057 4905 2060
rect 4939 2057 4951 2091
rect 5258 2088 5264 2100
rect 5219 2060 5264 2088
rect 4893 2051 4951 2057
rect 5258 2048 5264 2060
rect 5316 2048 5322 2100
rect 5353 2091 5411 2097
rect 5353 2057 5365 2091
rect 5399 2088 5411 2091
rect 5626 2088 5632 2100
rect 5399 2060 5632 2088
rect 5399 2057 5411 2060
rect 5353 2051 5411 2057
rect 5626 2048 5632 2060
rect 5684 2048 5690 2100
rect 6365 2091 6423 2097
rect 6365 2057 6377 2091
rect 6411 2088 6423 2091
rect 6638 2088 6644 2100
rect 6411 2060 6644 2088
rect 6411 2057 6423 2060
rect 6365 2051 6423 2057
rect 6638 2048 6644 2060
rect 6696 2048 6702 2100
rect 6822 2048 6828 2100
rect 6880 2088 6886 2100
rect 7282 2088 7288 2100
rect 6880 2060 7288 2088
rect 6880 2048 6886 2060
rect 7282 2048 7288 2060
rect 7340 2048 7346 2100
rect 9033 2091 9091 2097
rect 9033 2057 9045 2091
rect 9079 2057 9091 2091
rect 10594 2088 10600 2100
rect 10555 2060 10600 2088
rect 9033 2051 9091 2057
rect 3510 1980 3516 2032
rect 3568 1980 3574 2032
rect 7098 1980 7104 2032
rect 7156 2020 7162 2032
rect 7650 2020 7656 2032
rect 7156 1992 7656 2020
rect 7156 1980 7162 1992
rect 7650 1980 7656 1992
rect 7708 2020 7714 2032
rect 9048 2020 9076 2051
rect 10594 2048 10600 2060
rect 10652 2048 10658 2100
rect 11057 2091 11115 2097
rect 11057 2057 11069 2091
rect 11103 2088 11115 2091
rect 11238 2088 11244 2100
rect 11103 2060 11244 2088
rect 11103 2057 11115 2060
rect 11057 2051 11115 2057
rect 11238 2048 11244 2060
rect 11296 2048 11302 2100
rect 12618 2088 12624 2100
rect 12579 2060 12624 2088
rect 12618 2048 12624 2060
rect 12676 2048 12682 2100
rect 14550 2048 14556 2100
rect 14608 2088 14614 2100
rect 16942 2088 16948 2100
rect 14608 2060 14872 2088
rect 14608 2048 14614 2060
rect 9217 2023 9275 2029
rect 9217 2020 9229 2023
rect 7708 1992 8050 2020
rect 9048 1992 9229 2020
rect 7708 1980 7714 1992
rect 9217 1989 9229 1992
rect 9263 2020 9275 2023
rect 9263 1992 11192 2020
rect 9263 1989 9275 1992
rect 9217 1983 9275 1989
rect 3053 1955 3111 1961
rect 3053 1952 3065 1955
rect 3016 1924 3065 1952
rect 3016 1912 3022 1924
rect 3053 1921 3065 1924
rect 3099 1921 3111 1955
rect 3053 1915 3111 1921
rect 3329 1955 3387 1961
rect 3329 1921 3341 1955
rect 3375 1921 3387 1955
rect 3329 1915 3387 1921
rect 3421 1955 3479 1961
rect 3421 1921 3433 1955
rect 3467 1952 3479 1955
rect 3528 1952 3556 1980
rect 3467 1924 3556 1952
rect 3605 1955 3663 1961
rect 3467 1921 3479 1924
rect 3421 1915 3479 1921
rect 3605 1921 3617 1955
rect 3651 1921 3663 1955
rect 3878 1952 3884 1964
rect 3839 1924 3884 1952
rect 3605 1915 3663 1921
rect 2317 1887 2375 1893
rect 2317 1853 2329 1887
rect 2363 1853 2375 1887
rect 2317 1847 2375 1853
rect 2777 1887 2835 1893
rect 2777 1853 2789 1887
rect 2823 1884 2835 1887
rect 3513 1887 3571 1893
rect 3513 1884 3525 1887
rect 2823 1856 3525 1884
rect 2823 1853 2835 1856
rect 2777 1847 2835 1853
rect 3513 1853 3525 1856
rect 3559 1853 3571 1887
rect 3513 1847 3571 1853
rect 1964 1788 2544 1816
rect 2516 1760 2544 1788
rect 2590 1776 2596 1828
rect 2648 1816 2654 1828
rect 3237 1819 3295 1825
rect 3237 1816 3249 1819
rect 2648 1788 3249 1816
rect 2648 1776 2654 1788
rect 3237 1785 3249 1788
rect 3283 1785 3295 1819
rect 3620 1816 3648 1915
rect 3878 1912 3884 1924
rect 3936 1912 3942 1964
rect 5902 1912 5908 1964
rect 5960 1952 5966 1964
rect 6457 1955 6515 1961
rect 6457 1952 6469 1955
rect 5960 1924 6469 1952
rect 5960 1912 5966 1924
rect 6457 1921 6469 1924
rect 6503 1921 6515 1955
rect 6457 1915 6515 1921
rect 6914 1912 6920 1964
rect 6972 1952 6978 1964
rect 7282 1952 7288 1964
rect 6972 1924 7288 1952
rect 6972 1912 6978 1924
rect 7282 1912 7288 1924
rect 7340 1912 7346 1964
rect 9030 1912 9036 1964
rect 9088 1952 9094 1964
rect 9125 1955 9183 1961
rect 9125 1952 9137 1955
rect 9088 1924 9137 1952
rect 9088 1912 9094 1924
rect 9125 1921 9137 1924
rect 9171 1921 9183 1955
rect 9125 1915 9183 1921
rect 9306 1912 9312 1964
rect 9364 1952 9370 1964
rect 9401 1955 9459 1961
rect 9401 1952 9413 1955
rect 9364 1924 9413 1952
rect 9364 1912 9370 1924
rect 9401 1921 9413 1924
rect 9447 1952 9459 1955
rect 9582 1952 9588 1964
rect 9447 1924 9588 1952
rect 9447 1921 9459 1924
rect 9401 1915 9459 1921
rect 9582 1912 9588 1924
rect 9640 1912 9646 1964
rect 9876 1961 9904 1992
rect 11164 1961 11192 1992
rect 11974 1980 11980 2032
rect 12032 2020 12038 2032
rect 14737 2023 14795 2029
rect 14737 2020 14749 2023
rect 12032 1992 13032 2020
rect 12032 1980 12038 1992
rect 9861 1955 9919 1961
rect 9861 1921 9873 1955
rect 9907 1921 9919 1955
rect 10689 1955 10747 1961
rect 10689 1952 10701 1955
rect 9861 1915 9919 1921
rect 10244 1924 10701 1952
rect 5537 1887 5595 1893
rect 5537 1853 5549 1887
rect 5583 1884 5595 1887
rect 5718 1884 5724 1896
rect 5583 1856 5724 1884
rect 5583 1853 5595 1856
rect 5537 1847 5595 1853
rect 5718 1844 5724 1856
rect 5776 1884 5782 1896
rect 5994 1884 6000 1896
rect 5776 1856 6000 1884
rect 5776 1844 5782 1856
rect 5994 1844 6000 1856
rect 6052 1844 6058 1896
rect 6273 1887 6331 1893
rect 6273 1853 6285 1887
rect 6319 1884 6331 1887
rect 6546 1884 6552 1896
rect 6319 1856 6552 1884
rect 6319 1853 6331 1856
rect 6273 1847 6331 1853
rect 6546 1844 6552 1856
rect 6604 1884 6610 1896
rect 7006 1884 7012 1896
rect 6604 1856 7012 1884
rect 6604 1844 6610 1856
rect 7006 1844 7012 1856
rect 7064 1844 7070 1896
rect 7561 1887 7619 1893
rect 7561 1853 7573 1887
rect 7607 1884 7619 1887
rect 8294 1884 8300 1896
rect 7607 1856 8300 1884
rect 7607 1853 7619 1856
rect 7561 1847 7619 1853
rect 8294 1844 8300 1856
rect 8352 1844 8358 1896
rect 9950 1884 9956 1896
rect 9911 1856 9956 1884
rect 9950 1844 9956 1856
rect 10008 1844 10014 1896
rect 10244 1893 10272 1924
rect 10689 1921 10701 1924
rect 10735 1921 10747 1955
rect 10689 1915 10747 1921
rect 11149 1955 11207 1961
rect 11149 1921 11161 1955
rect 11195 1921 11207 1955
rect 11149 1915 11207 1921
rect 12529 1955 12587 1961
rect 12529 1921 12541 1955
rect 12575 1952 12587 1955
rect 12802 1952 12808 1964
rect 12575 1924 12808 1952
rect 12575 1921 12587 1924
rect 12529 1915 12587 1921
rect 12802 1912 12808 1924
rect 12860 1912 12866 1964
rect 13004 1961 13032 1992
rect 14016 1992 14749 2020
rect 12989 1955 13047 1961
rect 12989 1921 13001 1955
rect 13035 1921 13047 1955
rect 12989 1915 13047 1921
rect 10229 1887 10287 1893
rect 10229 1853 10241 1887
rect 10275 1853 10287 1887
rect 10229 1847 10287 1853
rect 10505 1887 10563 1893
rect 10505 1853 10517 1887
rect 10551 1853 10563 1887
rect 10505 1847 10563 1853
rect 6086 1816 6092 1828
rect 3620 1788 6092 1816
rect 3237 1779 3295 1785
rect 6086 1776 6092 1788
rect 6144 1776 6150 1828
rect 10520 1816 10548 1847
rect 12250 1844 12256 1896
rect 12308 1884 12314 1896
rect 14016 1893 14044 1992
rect 14737 1989 14749 1992
rect 14783 1989 14795 2023
rect 14737 1983 14795 1989
rect 14277 1955 14335 1961
rect 14277 1921 14289 1955
rect 14323 1921 14335 1955
rect 14458 1952 14464 1964
rect 14419 1924 14464 1952
rect 14277 1915 14335 1921
rect 14001 1887 14059 1893
rect 14001 1884 14013 1887
rect 12308 1856 14013 1884
rect 12308 1844 12314 1856
rect 14001 1853 14013 1856
rect 14047 1853 14059 1887
rect 14292 1884 14320 1915
rect 14458 1912 14464 1924
rect 14516 1912 14522 1964
rect 14642 1952 14648 1964
rect 14603 1924 14648 1952
rect 14642 1912 14648 1924
rect 14700 1912 14706 1964
rect 14553 1887 14611 1893
rect 14553 1884 14565 1887
rect 14292 1856 14565 1884
rect 14001 1847 14059 1853
rect 14553 1853 14565 1856
rect 14599 1853 14611 1887
rect 14844 1884 14872 2060
rect 14936 2060 16948 2088
rect 14936 1964 14964 2060
rect 16942 2048 16948 2060
rect 17000 2048 17006 2100
rect 14918 1912 14924 1964
rect 14976 1952 14982 1964
rect 15286 1952 15292 1964
rect 14976 1924 15069 1952
rect 15247 1924 15292 1952
rect 14976 1912 14982 1924
rect 15286 1912 15292 1924
rect 15344 1912 15350 1964
rect 15556 1955 15614 1961
rect 15556 1952 15568 1955
rect 15396 1924 15568 1952
rect 15194 1884 15200 1896
rect 14844 1856 15200 1884
rect 14553 1847 14611 1853
rect 15194 1844 15200 1856
rect 15252 1844 15258 1896
rect 15396 1884 15424 1924
rect 15556 1921 15568 1924
rect 15602 1952 15614 1955
rect 16482 1952 16488 1964
rect 15602 1924 16488 1952
rect 15602 1921 15614 1924
rect 15556 1915 15614 1921
rect 16482 1912 16488 1924
rect 16540 1912 16546 1964
rect 15304 1856 15424 1884
rect 10778 1816 10784 1828
rect 10520 1788 10784 1816
rect 10778 1776 10784 1788
rect 10836 1816 10842 1828
rect 14093 1819 14151 1825
rect 10836 1788 12940 1816
rect 10836 1776 10842 1788
rect 2498 1748 2504 1760
rect 2459 1720 2504 1748
rect 2498 1708 2504 1720
rect 2556 1708 2562 1760
rect 2866 1748 2872 1760
rect 2827 1720 2872 1748
rect 2866 1708 2872 1720
rect 2924 1708 2930 1760
rect 2961 1751 3019 1757
rect 2961 1717 2973 1751
rect 3007 1748 3019 1751
rect 3510 1748 3516 1760
rect 3007 1720 3516 1748
rect 3007 1717 3019 1720
rect 2961 1711 3019 1717
rect 3510 1708 3516 1720
rect 3568 1708 3574 1760
rect 6822 1748 6828 1760
rect 6783 1720 6828 1748
rect 6822 1708 6828 1720
rect 6880 1708 6886 1760
rect 7098 1748 7104 1760
rect 7059 1720 7104 1748
rect 7098 1708 7104 1720
rect 7156 1708 7162 1760
rect 9122 1708 9128 1760
rect 9180 1748 9186 1760
rect 9180 1720 9225 1748
rect 9180 1708 9186 1720
rect 11146 1708 11152 1760
rect 11204 1748 11210 1760
rect 12912 1757 12940 1788
rect 14093 1785 14105 1819
rect 14139 1816 14151 1819
rect 14642 1816 14648 1828
rect 14139 1788 14648 1816
rect 14139 1785 14151 1788
rect 14093 1779 14151 1785
rect 14642 1776 14648 1788
rect 14700 1776 14706 1828
rect 15102 1816 15108 1828
rect 15015 1788 15108 1816
rect 15102 1776 15108 1788
rect 15160 1816 15166 1828
rect 15304 1816 15332 1856
rect 15160 1788 15332 1816
rect 15160 1776 15166 1788
rect 11241 1751 11299 1757
rect 11241 1748 11253 1751
rect 11204 1720 11253 1748
rect 11204 1708 11210 1720
rect 11241 1717 11253 1720
rect 11287 1717 11299 1751
rect 11241 1711 11299 1717
rect 12897 1751 12955 1757
rect 12897 1717 12909 1751
rect 12943 1748 12955 1751
rect 12986 1748 12992 1760
rect 12943 1720 12992 1748
rect 12943 1717 12955 1720
rect 12897 1711 12955 1717
rect 12986 1708 12992 1720
rect 13044 1708 13050 1760
rect 14182 1708 14188 1760
rect 14240 1748 14246 1760
rect 16666 1748 16672 1760
rect 14240 1720 14285 1748
rect 16627 1720 16672 1748
rect 14240 1708 14246 1720
rect 16666 1708 16672 1720
rect 16724 1708 16730 1760
rect 0 1658 18860 1680
rect 0 1606 3110 1658
rect 3162 1606 3174 1658
rect 3226 1606 3238 1658
rect 3290 1606 3302 1658
rect 3354 1606 3366 1658
rect 3418 1606 6210 1658
rect 6262 1606 6274 1658
rect 6326 1606 6338 1658
rect 6390 1606 6402 1658
rect 6454 1606 6466 1658
rect 6518 1606 9310 1658
rect 9362 1606 9374 1658
rect 9426 1606 9438 1658
rect 9490 1606 9502 1658
rect 9554 1606 9566 1658
rect 9618 1606 12410 1658
rect 12462 1606 12474 1658
rect 12526 1606 12538 1658
rect 12590 1606 12602 1658
rect 12654 1606 12666 1658
rect 12718 1606 15510 1658
rect 15562 1606 15574 1658
rect 15626 1606 15638 1658
rect 15690 1606 15702 1658
rect 15754 1606 15766 1658
rect 15818 1606 18860 1658
rect 0 1584 18860 1606
rect 2958 1504 2964 1556
rect 3016 1544 3022 1556
rect 3694 1544 3700 1556
rect 3016 1516 3700 1544
rect 3016 1504 3022 1516
rect 3694 1504 3700 1516
rect 3752 1544 3758 1556
rect 3789 1547 3847 1553
rect 3789 1544 3801 1547
rect 3752 1516 3801 1544
rect 3752 1504 3758 1516
rect 3789 1513 3801 1516
rect 3835 1513 3847 1547
rect 5902 1544 5908 1556
rect 5863 1516 5908 1544
rect 3789 1507 3847 1513
rect 5902 1504 5908 1516
rect 5960 1504 5966 1556
rect 6086 1544 6092 1556
rect 6047 1516 6092 1544
rect 6086 1504 6092 1516
rect 6144 1504 6150 1556
rect 9950 1504 9956 1556
rect 10008 1544 10014 1556
rect 10229 1547 10287 1553
rect 10229 1544 10241 1547
rect 10008 1516 10241 1544
rect 10008 1504 10014 1516
rect 10229 1513 10241 1516
rect 10275 1513 10287 1547
rect 10229 1507 10287 1513
rect 11149 1547 11207 1553
rect 11149 1513 11161 1547
rect 11195 1544 11207 1547
rect 11974 1544 11980 1556
rect 11195 1516 11980 1544
rect 11195 1513 11207 1516
rect 11149 1507 11207 1513
rect 11974 1504 11980 1516
rect 12032 1504 12038 1556
rect 14182 1504 14188 1556
rect 14240 1544 14246 1556
rect 14829 1547 14887 1553
rect 14829 1544 14841 1547
rect 14240 1516 14841 1544
rect 14240 1504 14246 1516
rect 14829 1513 14841 1516
rect 14875 1513 14887 1547
rect 17586 1544 17592 1556
rect 17547 1516 17592 1544
rect 14829 1507 14887 1513
rect 17586 1504 17592 1516
rect 17644 1504 17650 1556
rect 2774 1436 2780 1488
rect 2832 1476 2838 1488
rect 3878 1476 3884 1488
rect 2832 1448 3884 1476
rect 2832 1436 2838 1448
rect 3878 1436 3884 1448
rect 3936 1436 3942 1488
rect 14458 1476 14464 1488
rect 6748 1448 11560 1476
rect 1210 1368 1216 1420
rect 1268 1408 1274 1420
rect 1305 1411 1363 1417
rect 1305 1408 1317 1411
rect 1268 1380 1317 1408
rect 1268 1368 1274 1380
rect 1305 1377 1317 1380
rect 1351 1377 1363 1411
rect 1305 1371 1363 1377
rect 1581 1411 1639 1417
rect 1581 1377 1593 1411
rect 1627 1408 1639 1411
rect 2866 1408 2872 1420
rect 1627 1380 2872 1408
rect 1627 1377 1639 1380
rect 1581 1371 1639 1377
rect 2866 1368 2872 1380
rect 2924 1368 2930 1420
rect 3053 1411 3111 1417
rect 3053 1377 3065 1411
rect 3099 1408 3111 1411
rect 5626 1408 5632 1420
rect 3099 1380 3924 1408
rect 5587 1380 5632 1408
rect 3099 1377 3111 1380
rect 3053 1371 3111 1377
rect 3421 1343 3479 1349
rect 3421 1340 3433 1343
rect 3344 1312 3433 1340
rect 3344 1284 3372 1312
rect 3421 1309 3433 1312
rect 3467 1309 3479 1343
rect 3421 1303 3479 1309
rect 3513 1343 3571 1349
rect 3513 1309 3525 1343
rect 3559 1340 3571 1343
rect 3694 1340 3700 1352
rect 3559 1312 3700 1340
rect 3559 1309 3571 1312
rect 3513 1303 3571 1309
rect 3694 1300 3700 1312
rect 3752 1300 3758 1352
rect 3896 1349 3924 1380
rect 5626 1368 5632 1380
rect 5684 1368 5690 1420
rect 5994 1368 6000 1420
rect 6052 1408 6058 1420
rect 6748 1417 6776 1448
rect 6733 1411 6791 1417
rect 6733 1408 6745 1411
rect 6052 1380 6745 1408
rect 6052 1368 6058 1380
rect 6733 1377 6745 1380
rect 6779 1377 6791 1411
rect 6733 1371 6791 1377
rect 7374 1368 7380 1420
rect 7432 1408 7438 1420
rect 9122 1408 9128 1420
rect 7432 1380 8708 1408
rect 9083 1380 9128 1408
rect 7432 1368 7438 1380
rect 8680 1352 8708 1380
rect 9122 1368 9128 1380
rect 9180 1368 9186 1420
rect 9968 1417 9996 1448
rect 11532 1420 11560 1448
rect 12912 1448 14464 1476
rect 9953 1411 10011 1417
rect 9953 1377 9965 1411
rect 9999 1377 10011 1411
rect 9953 1371 10011 1377
rect 10980 1380 11284 1408
rect 3881 1343 3939 1349
rect 3881 1309 3893 1343
rect 3927 1340 3939 1343
rect 4982 1340 4988 1352
rect 3927 1312 4988 1340
rect 3927 1309 3939 1312
rect 3881 1303 3939 1309
rect 4982 1300 4988 1312
rect 5040 1340 5046 1352
rect 5537 1343 5595 1349
rect 5537 1340 5549 1343
rect 5040 1312 5549 1340
rect 5040 1300 5046 1312
rect 5537 1309 5549 1312
rect 5583 1309 5595 1343
rect 5537 1303 5595 1309
rect 6457 1343 6515 1349
rect 6457 1309 6469 1343
rect 6503 1340 6515 1343
rect 6822 1340 6828 1352
rect 6503 1312 6828 1340
rect 6503 1309 6515 1312
rect 6457 1303 6515 1309
rect 6822 1300 6828 1312
rect 6880 1300 6886 1352
rect 8294 1300 8300 1352
rect 8352 1340 8358 1352
rect 8481 1343 8539 1349
rect 8481 1340 8493 1343
rect 8352 1312 8493 1340
rect 8352 1300 8358 1312
rect 8481 1309 8493 1312
rect 8527 1309 8539 1343
rect 8662 1340 8668 1352
rect 8623 1312 8668 1340
rect 8481 1303 8539 1309
rect 8662 1300 8668 1312
rect 8720 1300 8726 1352
rect 8754 1300 8760 1352
rect 8812 1340 8818 1352
rect 9861 1343 9919 1349
rect 8812 1312 8857 1340
rect 8812 1300 8818 1312
rect 9861 1309 9873 1343
rect 9907 1340 9919 1343
rect 10042 1340 10048 1352
rect 9907 1312 10048 1340
rect 9907 1309 9919 1312
rect 9861 1303 9919 1309
rect 10042 1300 10048 1312
rect 10100 1300 10106 1352
rect 10229 1343 10287 1349
rect 10229 1309 10241 1343
rect 10275 1309 10287 1343
rect 10229 1303 10287 1309
rect 2498 1164 2504 1216
rect 2556 1204 2562 1216
rect 2792 1204 2820 1258
rect 2866 1232 2872 1284
rect 2924 1272 2930 1284
rect 3237 1275 3295 1281
rect 3237 1272 3249 1275
rect 2924 1244 3249 1272
rect 2924 1232 2930 1244
rect 3237 1241 3249 1244
rect 3283 1241 3295 1275
rect 3237 1235 3295 1241
rect 3326 1232 3332 1284
rect 3384 1232 3390 1284
rect 6549 1275 6607 1281
rect 3436 1244 4108 1272
rect 3436 1204 3464 1244
rect 4080 1216 4108 1244
rect 6549 1241 6561 1275
rect 6595 1272 6607 1275
rect 6638 1272 6644 1284
rect 6595 1244 6644 1272
rect 6595 1241 6607 1244
rect 6549 1235 6607 1241
rect 6638 1232 6644 1244
rect 6696 1232 6702 1284
rect 10134 1232 10140 1284
rect 10192 1272 10198 1284
rect 10244 1272 10272 1303
rect 10410 1300 10416 1352
rect 10468 1340 10474 1352
rect 10980 1340 11008 1380
rect 11146 1340 11152 1352
rect 10468 1312 11008 1340
rect 11107 1312 11152 1340
rect 10468 1300 10474 1312
rect 11146 1300 11152 1312
rect 11204 1300 11210 1352
rect 11256 1349 11284 1380
rect 11514 1368 11520 1420
rect 11572 1408 11578 1420
rect 12912 1417 12940 1448
rect 14458 1436 14464 1448
rect 14516 1436 14522 1488
rect 12897 1411 12955 1417
rect 12897 1408 12909 1411
rect 11572 1380 12909 1408
rect 11572 1368 11578 1380
rect 12897 1377 12909 1380
rect 12943 1377 12955 1411
rect 12897 1371 12955 1377
rect 12986 1368 12992 1420
rect 13044 1408 13050 1420
rect 13817 1411 13875 1417
rect 13817 1408 13829 1411
rect 13044 1380 13829 1408
rect 13044 1368 13050 1380
rect 13817 1377 13829 1380
rect 13863 1377 13875 1411
rect 14918 1408 14924 1420
rect 13817 1371 13875 1377
rect 13924 1380 14924 1408
rect 11241 1343 11299 1349
rect 11241 1309 11253 1343
rect 11287 1309 11299 1343
rect 11241 1303 11299 1309
rect 12805 1343 12863 1349
rect 12805 1309 12817 1343
rect 12851 1340 12863 1343
rect 13722 1340 13728 1352
rect 12851 1312 13728 1340
rect 12851 1309 12863 1312
rect 12805 1303 12863 1309
rect 13722 1300 13728 1312
rect 13780 1340 13786 1352
rect 13924 1340 13952 1380
rect 14918 1368 14924 1380
rect 14976 1368 14982 1420
rect 15194 1408 15200 1420
rect 15155 1380 15200 1408
rect 15194 1368 15200 1380
rect 15252 1368 15258 1420
rect 16114 1408 16120 1420
rect 16075 1380 16120 1408
rect 16114 1368 16120 1380
rect 16172 1368 16178 1420
rect 13780 1312 13952 1340
rect 13780 1300 13786 1312
rect 14734 1300 14740 1352
rect 14792 1340 14798 1352
rect 15013 1343 15071 1349
rect 15013 1340 15025 1343
rect 14792 1312 15025 1340
rect 14792 1300 14798 1312
rect 15013 1309 15025 1312
rect 15059 1309 15071 1343
rect 15838 1340 15844 1352
rect 15799 1312 15844 1340
rect 15013 1303 15071 1309
rect 15838 1300 15844 1312
rect 15896 1300 15902 1352
rect 17770 1340 17776 1352
rect 17731 1312 17776 1340
rect 17770 1300 17776 1312
rect 17828 1300 17834 1352
rect 17862 1300 17868 1352
rect 17920 1340 17926 1352
rect 18046 1340 18052 1352
rect 17920 1312 17965 1340
rect 18007 1312 18052 1340
rect 17920 1300 17926 1312
rect 18046 1300 18052 1312
rect 18104 1300 18110 1352
rect 18141 1343 18199 1349
rect 18141 1309 18153 1343
rect 18187 1340 18199 1343
rect 18414 1340 18420 1352
rect 18187 1312 18420 1340
rect 18187 1309 18199 1312
rect 18141 1303 18199 1309
rect 18414 1300 18420 1312
rect 18472 1300 18478 1352
rect 10873 1275 10931 1281
rect 10873 1272 10885 1275
rect 10192 1244 10885 1272
rect 10192 1232 10198 1244
rect 10873 1241 10885 1244
rect 10919 1241 10931 1275
rect 10873 1235 10931 1241
rect 11057 1275 11115 1281
rect 11057 1241 11069 1275
rect 11103 1272 11115 1275
rect 11333 1275 11391 1281
rect 11333 1272 11345 1275
rect 11103 1244 11345 1272
rect 11103 1241 11115 1244
rect 11057 1235 11115 1241
rect 11333 1241 11345 1244
rect 11379 1241 11391 1275
rect 11333 1235 11391 1241
rect 12713 1275 12771 1281
rect 12713 1241 12725 1275
rect 12759 1272 12771 1275
rect 12759 1244 13308 1272
rect 12759 1241 12771 1244
rect 12713 1235 12771 1241
rect 2556 1176 3464 1204
rect 3513 1207 3571 1213
rect 2556 1164 2562 1176
rect 3513 1173 3525 1207
rect 3559 1204 3571 1207
rect 3602 1204 3608 1216
rect 3559 1176 3608 1204
rect 3559 1173 3571 1176
rect 3513 1167 3571 1173
rect 3602 1164 3608 1176
rect 3660 1164 3666 1216
rect 4062 1204 4068 1216
rect 3975 1176 4068 1204
rect 4062 1164 4068 1176
rect 4120 1204 4126 1216
rect 7098 1204 7104 1216
rect 4120 1176 7104 1204
rect 4120 1164 4126 1176
rect 7098 1164 7104 1176
rect 7156 1164 7162 1216
rect 8754 1164 8760 1216
rect 8812 1204 8818 1216
rect 9401 1207 9459 1213
rect 9401 1204 9413 1207
rect 8812 1176 9413 1204
rect 8812 1164 8818 1176
rect 9401 1173 9413 1176
rect 9447 1173 9459 1207
rect 9401 1167 9459 1173
rect 9769 1207 9827 1213
rect 9769 1173 9781 1207
rect 9815 1204 9827 1207
rect 10318 1204 10324 1216
rect 9815 1176 10324 1204
rect 9815 1173 9827 1176
rect 9769 1167 9827 1173
rect 10318 1164 10324 1176
rect 10376 1164 10382 1216
rect 10888 1204 10916 1235
rect 11790 1204 11796 1216
rect 10888 1176 11796 1204
rect 11790 1164 11796 1176
rect 11848 1164 11854 1216
rect 12250 1164 12256 1216
rect 12308 1204 12314 1216
rect 13280 1213 13308 1244
rect 13354 1232 13360 1284
rect 13412 1272 13418 1284
rect 14277 1275 14335 1281
rect 14277 1272 14289 1275
rect 13412 1244 14289 1272
rect 13412 1232 13418 1244
rect 14277 1241 14289 1244
rect 14323 1272 14335 1275
rect 14918 1272 14924 1284
rect 14323 1244 14924 1272
rect 14323 1241 14335 1244
rect 14277 1235 14335 1241
rect 14918 1232 14924 1244
rect 14976 1272 14982 1284
rect 15378 1272 15384 1284
rect 14976 1244 15384 1272
rect 14976 1232 14982 1244
rect 15378 1232 15384 1244
rect 15436 1272 15442 1284
rect 15657 1275 15715 1281
rect 15657 1272 15669 1275
rect 15436 1244 15669 1272
rect 15436 1232 15442 1244
rect 15657 1241 15669 1244
rect 15703 1272 15715 1275
rect 15703 1244 16606 1272
rect 15703 1241 15715 1244
rect 15657 1235 15715 1241
rect 18230 1232 18236 1284
rect 18288 1272 18294 1284
rect 18325 1275 18383 1281
rect 18325 1272 18337 1275
rect 18288 1244 18337 1272
rect 18288 1232 18294 1244
rect 18325 1241 18337 1244
rect 18371 1241 18383 1275
rect 18325 1235 18383 1241
rect 12345 1207 12403 1213
rect 12345 1204 12357 1207
rect 12308 1176 12357 1204
rect 12308 1164 12314 1176
rect 12345 1173 12357 1176
rect 12391 1173 12403 1207
rect 12345 1167 12403 1173
rect 13265 1207 13323 1213
rect 13265 1173 13277 1207
rect 13311 1173 13323 1207
rect 13630 1204 13636 1216
rect 13591 1176 13636 1204
rect 13265 1167 13323 1173
rect 13630 1164 13636 1176
rect 13688 1164 13694 1216
rect 17954 1164 17960 1216
rect 18012 1204 18018 1216
rect 18049 1207 18107 1213
rect 18049 1204 18061 1207
rect 18012 1176 18061 1204
rect 18012 1164 18018 1176
rect 18049 1173 18061 1176
rect 18095 1173 18107 1207
rect 18506 1204 18512 1216
rect 18467 1176 18512 1204
rect 18049 1167 18107 1173
rect 18506 1164 18512 1176
rect 18564 1164 18570 1216
rect 0 1114 18860 1136
rect 0 1062 4660 1114
rect 4712 1062 4724 1114
rect 4776 1062 4788 1114
rect 4840 1062 4852 1114
rect 4904 1062 4916 1114
rect 4968 1062 7760 1114
rect 7812 1062 7824 1114
rect 7876 1062 7888 1114
rect 7940 1062 7952 1114
rect 8004 1062 8016 1114
rect 8068 1062 10860 1114
rect 10912 1062 10924 1114
rect 10976 1062 10988 1114
rect 11040 1062 11052 1114
rect 11104 1062 11116 1114
rect 11168 1062 13960 1114
rect 14012 1062 14024 1114
rect 14076 1062 14088 1114
rect 14140 1062 14152 1114
rect 14204 1062 14216 1114
rect 14268 1062 17060 1114
rect 17112 1062 17124 1114
rect 17176 1062 17188 1114
rect 17240 1062 17252 1114
rect 17304 1062 17316 1114
rect 17368 1062 18860 1114
rect 0 1040 18860 1062
rect 2317 1003 2375 1009
rect 2317 969 2329 1003
rect 2363 1000 2375 1003
rect 2498 1000 2504 1012
rect 2363 972 2504 1000
rect 2363 969 2375 972
rect 2317 963 2375 969
rect 2498 960 2504 972
rect 2556 960 2562 1012
rect 5626 960 5632 1012
rect 5684 1000 5690 1012
rect 5905 1003 5963 1009
rect 5905 1000 5917 1003
rect 5684 972 5917 1000
rect 5684 960 5690 972
rect 5905 969 5917 972
rect 5951 969 5963 1003
rect 7098 1000 7104 1012
rect 7011 972 7104 1000
rect 5905 963 5963 969
rect 7098 960 7104 972
rect 7156 1000 7162 1012
rect 10318 1000 10324 1012
rect 7156 972 8156 1000
rect 10279 972 10324 1000
rect 7156 960 7162 972
rect 4062 932 4068 944
rect 3910 904 4068 932
rect 4062 892 4068 904
rect 4120 892 4126 944
rect 5442 932 5448 944
rect 4632 904 5212 932
rect 5403 904 5448 932
rect 2501 867 2559 873
rect 2501 833 2513 867
rect 2547 864 2559 867
rect 2590 864 2596 876
rect 2547 836 2596 864
rect 2547 833 2559 836
rect 2501 827 2559 833
rect 2590 824 2596 836
rect 2648 824 2654 876
rect 4632 873 4660 904
rect 5184 876 5212 904
rect 5442 892 5448 904
rect 5500 892 5506 944
rect 5644 904 6040 932
rect 8128 918 8156 972
rect 10318 960 10324 972
rect 10376 960 10382 1012
rect 11330 960 11336 1012
rect 11388 1000 11394 1012
rect 11425 1003 11483 1009
rect 11425 1000 11437 1003
rect 11388 972 11437 1000
rect 11388 960 11394 972
rect 11425 969 11437 972
rect 11471 1000 11483 1003
rect 13354 1000 13360 1012
rect 11471 972 13360 1000
rect 11471 969 11483 972
rect 11425 963 11483 969
rect 9171 935 9229 941
rect 4295 867 4353 873
rect 4295 833 4307 867
rect 4341 864 4353 867
rect 4617 867 4675 873
rect 4617 864 4629 867
rect 4341 836 4629 864
rect 4341 833 4353 836
rect 4295 827 4353 833
rect 4617 833 4629 836
rect 4663 833 4675 867
rect 4982 864 4988 876
rect 4943 836 4988 864
rect 4617 827 4675 833
rect 4982 824 4988 836
rect 5040 824 5046 876
rect 5166 864 5172 876
rect 5079 836 5172 864
rect 5166 824 5172 836
rect 5224 864 5230 876
rect 5644 864 5672 904
rect 6012 873 6040 904
rect 9171 901 9183 935
rect 9217 932 9229 935
rect 9769 935 9827 941
rect 9769 932 9781 935
rect 9217 904 9781 932
rect 9217 901 9229 904
rect 9171 895 9229 901
rect 9769 901 9781 904
rect 9815 932 9827 935
rect 10410 932 10416 944
rect 9815 904 10416 932
rect 9815 901 9827 904
rect 9769 895 9827 901
rect 10410 892 10416 904
rect 10468 892 10474 944
rect 11790 932 11796 944
rect 11751 904 11796 932
rect 11790 892 11796 904
rect 11848 892 11854 944
rect 12820 918 12848 972
rect 13354 960 13360 972
rect 13412 960 13418 1012
rect 13630 960 13636 1012
rect 13688 1000 13694 1012
rect 14185 1003 14243 1009
rect 14185 1000 14197 1003
rect 13688 972 14197 1000
rect 13688 960 13694 972
rect 14185 969 14197 972
rect 14231 969 14243 1003
rect 14185 963 14243 969
rect 15286 960 15292 1012
rect 15344 1000 15350 1012
rect 18230 1000 18236 1012
rect 15344 972 16528 1000
rect 18191 972 18236 1000
rect 15344 960 15350 972
rect 14458 932 14464 944
rect 14419 904 14464 932
rect 14458 892 14464 904
rect 14516 892 14522 944
rect 14918 892 14924 944
rect 14976 932 14982 944
rect 14976 904 15042 932
rect 14976 892 14982 904
rect 5224 836 5672 864
rect 5721 867 5779 873
rect 5224 824 5230 836
rect 5721 833 5733 867
rect 5767 864 5779 867
rect 5813 867 5871 873
rect 5813 864 5825 867
rect 5767 836 5825 864
rect 5767 833 5779 836
rect 5721 827 5779 833
rect 5813 833 5825 836
rect 5859 833 5871 867
rect 5813 827 5871 833
rect 5997 867 6055 873
rect 5997 833 6009 867
rect 6043 833 6055 867
rect 6457 867 6515 873
rect 6457 864 6469 867
rect 5997 827 6055 833
rect 6104 836 6469 864
rect 2866 796 2872 808
rect 2827 768 2872 796
rect 2866 756 2872 768
rect 2924 756 2930 808
rect 3878 756 3884 808
rect 3936 796 3942 808
rect 5350 796 5356 808
rect 3936 768 5356 796
rect 3936 756 3942 768
rect 5350 756 5356 768
rect 5408 796 5414 808
rect 5736 796 5764 827
rect 5408 768 5764 796
rect 5408 756 5414 768
rect 5902 756 5908 808
rect 5960 796 5966 808
rect 6104 796 6132 836
rect 6457 833 6469 836
rect 6503 833 6515 867
rect 6457 827 6515 833
rect 7282 824 7288 876
rect 7340 864 7346 876
rect 7377 867 7435 873
rect 7377 864 7389 867
rect 7340 836 7389 864
rect 7340 824 7346 836
rect 7377 833 7389 836
rect 7423 833 7435 867
rect 7377 827 7435 833
rect 9030 824 9036 876
rect 9088 864 9094 876
rect 9677 867 9735 873
rect 9677 864 9689 867
rect 9088 836 9689 864
rect 9088 824 9094 836
rect 9677 833 9689 836
rect 9723 864 9735 867
rect 9723 836 9812 864
rect 9723 833 9735 836
rect 9677 827 9735 833
rect 5960 768 6132 796
rect 6273 799 6331 805
rect 5960 756 5966 768
rect 6273 765 6285 799
rect 6319 765 6331 799
rect 6273 759 6331 765
rect 5442 688 5448 740
rect 5500 728 5506 740
rect 6288 728 6316 759
rect 6362 756 6368 808
rect 6420 796 6426 808
rect 7742 796 7748 808
rect 6420 768 6465 796
rect 7703 768 7748 796
rect 6420 756 6426 768
rect 7742 756 7748 768
rect 7800 756 7806 808
rect 6546 728 6552 740
rect 5500 700 6552 728
rect 5500 688 5506 700
rect 6546 688 6552 700
rect 6604 688 6610 740
rect 4522 660 4528 672
rect 4483 632 4528 660
rect 4522 620 4528 632
rect 4580 620 4586 672
rect 6822 660 6828 672
rect 6783 632 6828 660
rect 6822 620 6828 632
rect 6880 620 6886 672
rect 9674 660 9680 672
rect 9635 632 9680 660
rect 9674 620 9680 632
rect 9732 620 9738 672
rect 9784 660 9812 836
rect 9858 824 9864 876
rect 9916 864 9922 876
rect 9953 867 10011 873
rect 9953 864 9965 867
rect 9916 836 9965 864
rect 9916 824 9922 836
rect 9953 833 9965 836
rect 9999 833 10011 867
rect 9953 827 10011 833
rect 9968 728 9996 827
rect 10502 824 10508 876
rect 10560 864 10566 876
rect 10689 867 10747 873
rect 10689 864 10701 867
rect 10560 836 10701 864
rect 10560 824 10566 836
rect 10689 833 10701 836
rect 10735 833 10747 867
rect 10689 827 10747 833
rect 10781 867 10839 873
rect 10781 833 10793 867
rect 10827 864 10839 867
rect 10962 864 10968 876
rect 10827 836 10968 864
rect 10827 833 10839 836
rect 10781 827 10839 833
rect 10962 824 10968 836
rect 11020 824 11026 876
rect 11606 864 11612 876
rect 11519 836 11612 864
rect 11606 824 11612 836
rect 11664 824 11670 876
rect 11882 864 11888 876
rect 11716 836 11888 864
rect 10870 756 10876 808
rect 10928 796 10934 808
rect 10928 768 10973 796
rect 10928 756 10934 768
rect 11624 728 11652 824
rect 9968 700 11652 728
rect 11716 660 11744 836
rect 11882 824 11888 836
rect 11940 824 11946 876
rect 12066 864 12072 876
rect 12027 836 12072 864
rect 12066 824 12072 836
rect 12124 824 12130 876
rect 16500 873 16528 972
rect 18230 960 18236 972
rect 18288 960 18294 1012
rect 16942 892 16948 944
rect 17000 932 17006 944
rect 17098 935 17156 941
rect 17098 932 17110 935
rect 17000 904 17110 932
rect 17000 892 17006 904
rect 17098 901 17110 904
rect 17144 901 17156 935
rect 17098 895 17156 901
rect 14001 867 14059 873
rect 14001 833 14013 867
rect 14047 833 14059 867
rect 14001 827 14059 833
rect 16485 867 16543 873
rect 16485 833 16497 867
rect 16531 864 16543 867
rect 16853 867 16911 873
rect 16853 864 16865 867
rect 16531 836 16865 864
rect 16531 833 16543 836
rect 16485 827 16543 833
rect 16853 833 16865 836
rect 16899 833 16911 867
rect 18506 864 18512 876
rect 18467 836 18512 864
rect 16853 827 16911 833
rect 12345 799 12403 805
rect 12345 765 12357 799
rect 12391 796 12403 799
rect 12802 796 12808 808
rect 12391 768 12808 796
rect 12391 765 12403 768
rect 12345 759 12403 765
rect 12802 756 12808 768
rect 12860 756 12866 808
rect 13814 796 13820 808
rect 13775 768 13820 796
rect 13814 756 13820 768
rect 13872 796 13878 808
rect 14016 796 14044 827
rect 18506 824 18512 836
rect 18564 824 18570 876
rect 16206 796 16212 808
rect 13872 768 14044 796
rect 16167 768 16212 796
rect 13872 756 13878 768
rect 16206 756 16212 768
rect 16264 756 16270 808
rect 17862 688 17868 740
rect 17920 728 17926 740
rect 18325 731 18383 737
rect 18325 728 18337 731
rect 17920 700 18337 728
rect 17920 688 17926 700
rect 18325 697 18337 700
rect 18371 697 18383 731
rect 18325 691 18383 697
rect 9784 632 11744 660
rect 11885 663 11943 669
rect 11885 629 11897 663
rect 11931 660 11943 663
rect 12158 660 12164 672
rect 11931 632 12164 660
rect 11931 629 11943 632
rect 11885 623 11943 629
rect 12158 620 12164 632
rect 12216 620 12222 672
rect 0 570 18860 592
rect 0 518 3110 570
rect 3162 518 3174 570
rect 3226 518 3238 570
rect 3290 518 3302 570
rect 3354 518 3366 570
rect 3418 518 6210 570
rect 6262 518 6274 570
rect 6326 518 6338 570
rect 6390 518 6402 570
rect 6454 518 6466 570
rect 6518 518 9310 570
rect 9362 518 9374 570
rect 9426 518 9438 570
rect 9490 518 9502 570
rect 9554 518 9566 570
rect 9618 518 12410 570
rect 12462 518 12474 570
rect 12526 518 12538 570
rect 12590 518 12602 570
rect 12654 518 12666 570
rect 12718 518 15510 570
rect 15562 518 15574 570
rect 15626 518 15638 570
rect 15690 518 15702 570
rect 15754 518 15766 570
rect 15818 518 18860 570
rect 0 496 18860 518
rect 2866 416 2872 468
rect 2924 456 2930 468
rect 3145 459 3203 465
rect 3145 456 3157 459
rect 2924 428 3157 456
rect 2924 416 2930 428
rect 3145 425 3157 428
rect 3191 425 3203 459
rect 3145 419 3203 425
rect 3237 459 3295 465
rect 3237 425 3249 459
rect 3283 456 3295 459
rect 3602 456 3608 468
rect 3283 428 3608 456
rect 3283 425 3295 428
rect 3237 419 3295 425
rect 3602 416 3608 428
rect 3660 416 3666 468
rect 5721 459 5779 465
rect 5721 425 5733 459
rect 5767 456 5779 459
rect 5902 456 5908 468
rect 5767 428 5908 456
rect 5767 425 5779 428
rect 5721 419 5779 425
rect 5902 416 5908 428
rect 5960 416 5966 468
rect 7742 416 7748 468
rect 7800 456 7806 468
rect 8481 459 8539 465
rect 8481 456 8493 459
rect 7800 428 8493 456
rect 7800 416 7806 428
rect 8481 425 8493 428
rect 8527 425 8539 459
rect 10502 456 10508 468
rect 10463 428 10508 456
rect 8481 419 8539 425
rect 10502 416 10508 428
rect 10560 416 10566 468
rect 12802 456 12808 468
rect 12763 428 12808 456
rect 12802 416 12808 428
rect 12860 416 12866 468
rect 14642 416 14648 468
rect 14700 456 14706 468
rect 14737 459 14795 465
rect 14737 456 14749 459
rect 14700 428 14749 456
rect 14700 416 14706 428
rect 14737 425 14749 428
rect 14783 425 14795 459
rect 14737 419 14795 425
rect 15105 459 15163 465
rect 15105 425 15117 459
rect 15151 456 15163 459
rect 16206 456 16212 468
rect 15151 428 16212 456
rect 15151 425 15163 428
rect 15105 419 15163 425
rect 16206 416 16212 428
rect 16264 416 16270 468
rect 16574 416 16580 468
rect 16632 456 16638 468
rect 17313 459 17371 465
rect 17313 456 17325 459
rect 16632 428 17325 456
rect 16632 416 16638 428
rect 17313 425 17325 428
rect 17359 425 17371 459
rect 17313 419 17371 425
rect 17681 459 17739 465
rect 17681 425 17693 459
rect 17727 456 17739 459
rect 18046 456 18052 468
rect 17727 428 18052 456
rect 17727 425 17739 428
rect 17681 419 17739 425
rect 18046 416 18052 428
rect 18104 416 18110 468
rect 18141 459 18199 465
rect 18141 425 18153 459
rect 18187 425 18199 459
rect 18141 419 18199 425
rect 6089 391 6147 397
rect 6089 388 6101 391
rect 3896 360 6101 388
rect 3053 323 3111 329
rect 3053 289 3065 323
rect 3099 320 3111 323
rect 3789 323 3847 329
rect 3789 320 3801 323
rect 3099 292 3801 320
rect 3099 289 3111 292
rect 3053 283 3111 289
rect 3789 289 3801 292
rect 3835 289 3847 323
rect 3789 283 3847 289
rect 3329 255 3387 261
rect 3329 221 3341 255
rect 3375 221 3387 255
rect 3329 215 3387 221
rect 3344 184 3372 215
rect 3602 212 3608 264
rect 3660 252 3666 264
rect 3896 261 3924 360
rect 6089 357 6101 360
rect 6135 357 6147 391
rect 18156 388 18184 419
rect 18414 416 18420 468
rect 18472 456 18478 468
rect 18509 459 18567 465
rect 18509 456 18521 459
rect 18472 428 18521 456
rect 18472 416 18478 428
rect 18509 425 18521 428
rect 18555 425 18567 459
rect 18509 419 18567 425
rect 6089 351 6147 357
rect 17236 360 18184 388
rect 5350 320 5356 332
rect 5311 292 5356 320
rect 5350 280 5356 292
rect 5408 280 5414 332
rect 5994 280 6000 332
rect 6052 320 6058 332
rect 6641 323 6699 329
rect 6641 320 6653 323
rect 6052 292 6653 320
rect 6052 280 6058 292
rect 6641 289 6653 292
rect 6687 289 6699 323
rect 8754 320 8760 332
rect 8715 292 8760 320
rect 6641 283 6699 289
rect 8754 280 8760 292
rect 8812 280 8818 332
rect 9125 323 9183 329
rect 9125 289 9137 323
rect 9171 320 9183 323
rect 9674 320 9680 332
rect 9171 292 9680 320
rect 9171 289 9183 292
rect 9125 283 9183 289
rect 9674 280 9680 292
rect 9732 280 9738 332
rect 10134 320 10140 332
rect 10095 292 10140 320
rect 10134 280 10140 292
rect 10192 280 10198 332
rect 12158 320 12164 332
rect 12119 292 12164 320
rect 12158 280 12164 292
rect 12216 280 12222 332
rect 12250 280 12256 332
rect 12308 320 12314 332
rect 12529 323 12587 329
rect 12529 320 12541 323
rect 12308 292 12541 320
rect 12308 280 12314 292
rect 12529 289 12541 292
rect 12575 289 12587 323
rect 12529 283 12587 289
rect 12618 280 12624 332
rect 12676 320 12682 332
rect 12676 292 14964 320
rect 12676 280 12682 292
rect 3697 255 3755 261
rect 3697 252 3709 255
rect 3660 224 3709 252
rect 3660 212 3666 224
rect 3697 221 3709 224
rect 3743 221 3755 255
rect 3697 215 3755 221
rect 3881 255 3939 261
rect 3881 221 3893 255
rect 3927 221 3939 255
rect 3881 215 3939 221
rect 5166 212 5172 264
rect 5224 252 5230 264
rect 5445 255 5503 261
rect 5445 252 5457 255
rect 5224 224 5457 252
rect 5224 212 5230 224
rect 5445 221 5457 224
rect 5491 221 5503 255
rect 5445 215 5503 221
rect 6457 255 6515 261
rect 6457 221 6469 255
rect 6503 252 6515 255
rect 6822 252 6828 264
rect 6503 224 6828 252
rect 6503 221 6515 224
rect 6457 215 6515 221
rect 6822 212 6828 224
rect 6880 212 6886 264
rect 8662 252 8668 264
rect 8623 224 8668 252
rect 8662 212 8668 224
rect 8720 212 8726 264
rect 10229 255 10287 261
rect 10229 221 10241 255
rect 10275 252 10287 255
rect 10410 252 10416 264
rect 10275 224 10416 252
rect 10275 221 10287 224
rect 10229 215 10287 221
rect 10410 212 10416 224
rect 10468 212 10474 264
rect 14642 252 14648 264
rect 14603 224 14648 252
rect 14642 212 14648 224
rect 14700 212 14706 264
rect 14936 261 14964 292
rect 14921 255 14979 261
rect 14921 221 14933 255
rect 14967 221 14979 255
rect 14921 215 14979 221
rect 16666 212 16672 264
rect 16724 252 16730 264
rect 17236 261 17264 360
rect 17221 255 17279 261
rect 17221 252 17233 255
rect 16724 224 17233 252
rect 16724 212 16730 224
rect 17221 221 17233 224
rect 17267 221 17279 255
rect 17221 215 17279 221
rect 18049 255 18107 261
rect 18049 221 18061 255
rect 18095 252 18107 255
rect 18138 252 18144 264
rect 18095 224 18144 252
rect 18095 221 18107 224
rect 18049 215 18107 221
rect 18138 212 18144 224
rect 18196 212 18202 264
rect 3510 184 3516 196
rect 3344 156 3516 184
rect 3510 144 3516 156
rect 3568 184 3574 196
rect 4522 184 4528 196
rect 3568 156 4528 184
rect 3568 144 3574 156
rect 4522 144 4528 156
rect 4580 144 4586 196
rect 6549 187 6607 193
rect 6549 153 6561 187
rect 6595 184 6607 187
rect 6638 184 6644 196
rect 6595 156 6644 184
rect 6595 153 6607 156
rect 6549 147 6607 153
rect 6638 144 6644 156
rect 6696 144 6702 196
rect 0 26 18860 48
rect 0 -26 4660 26
rect 4712 -26 4724 26
rect 4776 -26 4788 26
rect 4840 -26 4852 26
rect 4904 -26 4916 26
rect 4968 -26 7760 26
rect 7812 -26 7824 26
rect 7876 -26 7888 26
rect 7940 -26 7952 26
rect 8004 -26 8016 26
rect 8068 -26 10860 26
rect 10912 -26 10924 26
rect 10976 -26 10988 26
rect 11040 -26 11052 26
rect 11104 -26 11116 26
rect 11168 -26 13960 26
rect 14012 -26 14024 26
rect 14076 -26 14088 26
rect 14140 -26 14152 26
rect 14204 -26 14216 26
rect 14268 -26 17060 26
rect 17112 -26 17124 26
rect 17176 -26 17188 26
rect 17240 -26 17252 26
rect 17304 -26 17316 26
rect 17368 -26 18860 26
rect 0 -48 18860 -26
<< via1 >>
rect 4660 10854 4712 10906
rect 4724 10854 4776 10906
rect 4788 10854 4840 10906
rect 4852 10854 4904 10906
rect 4916 10854 4968 10906
rect 7760 10854 7812 10906
rect 7824 10854 7876 10906
rect 7888 10854 7940 10906
rect 7952 10854 8004 10906
rect 8016 10854 8068 10906
rect 10860 10854 10912 10906
rect 10924 10854 10976 10906
rect 10988 10854 11040 10906
rect 11052 10854 11104 10906
rect 11116 10854 11168 10906
rect 13960 10854 14012 10906
rect 14024 10854 14076 10906
rect 14088 10854 14140 10906
rect 14152 10854 14204 10906
rect 14216 10854 14268 10906
rect 17060 10854 17112 10906
rect 17124 10854 17176 10906
rect 17188 10854 17240 10906
rect 17252 10854 17304 10906
rect 17316 10854 17368 10906
rect 2412 10752 2464 10804
rect 2044 10684 2096 10736
rect 2412 10616 2464 10668
rect 7104 10752 7156 10804
rect 9956 10752 10008 10804
rect 12808 10752 12860 10804
rect 14740 10752 14792 10804
rect 13544 10727 13596 10736
rect 13544 10693 13553 10727
rect 13553 10693 13587 10727
rect 13587 10693 13596 10727
rect 13544 10684 13596 10693
rect 2872 10616 2924 10668
rect 7472 10659 7524 10668
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 2964 10591 3016 10600
rect 572 10412 624 10464
rect 2964 10557 2973 10591
rect 2973 10557 3007 10591
rect 3007 10557 3016 10591
rect 2964 10548 3016 10557
rect 11244 10616 11296 10668
rect 11796 10616 11848 10668
rect 11152 10548 11204 10600
rect 14648 10548 14700 10600
rect 13728 10480 13780 10532
rect 13912 10480 13964 10532
rect 15108 10659 15160 10668
rect 15108 10625 15117 10659
rect 15117 10625 15151 10659
rect 15151 10625 15160 10659
rect 15108 10616 15160 10625
rect 15292 10616 15344 10668
rect 18052 10659 18104 10668
rect 18052 10625 18061 10659
rect 18061 10625 18095 10659
rect 18095 10625 18104 10659
rect 18052 10616 18104 10625
rect 18788 10616 18840 10668
rect 2504 10412 2556 10464
rect 11060 10455 11112 10464
rect 11060 10421 11069 10455
rect 11069 10421 11103 10455
rect 11103 10421 11112 10455
rect 11060 10412 11112 10421
rect 11612 10412 11664 10464
rect 14372 10412 14424 10464
rect 14832 10412 14884 10464
rect 16212 10412 16264 10464
rect 3110 10310 3162 10362
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 3302 10310 3354 10362
rect 3366 10310 3418 10362
rect 6210 10310 6262 10362
rect 6274 10310 6326 10362
rect 6338 10310 6390 10362
rect 6402 10310 6454 10362
rect 6466 10310 6518 10362
rect 9310 10310 9362 10362
rect 9374 10310 9426 10362
rect 9438 10310 9490 10362
rect 9502 10310 9554 10362
rect 9566 10310 9618 10362
rect 12410 10310 12462 10362
rect 12474 10310 12526 10362
rect 12538 10310 12590 10362
rect 12602 10310 12654 10362
rect 12666 10310 12718 10362
rect 15510 10310 15562 10362
rect 15574 10310 15626 10362
rect 15638 10310 15690 10362
rect 15702 10310 15754 10362
rect 15766 10310 15818 10362
rect 1400 10251 1452 10260
rect 1400 10217 1409 10251
rect 1409 10217 1443 10251
rect 1443 10217 1452 10251
rect 1400 10208 1452 10217
rect 4436 10208 4488 10260
rect 5908 10208 5960 10260
rect 6828 10208 6880 10260
rect 1400 10004 1452 10056
rect 2964 10047 3016 10056
rect 2964 10013 2973 10047
rect 2973 10013 3007 10047
rect 3007 10013 3016 10047
rect 2964 10004 3016 10013
rect 3332 10004 3384 10056
rect 3700 10140 3752 10192
rect 7472 10208 7524 10260
rect 12992 10208 13044 10260
rect 13544 10208 13596 10260
rect 18052 10208 18104 10260
rect 14924 10140 14976 10192
rect 3976 10072 4028 10124
rect 6092 10115 6144 10124
rect 6092 10081 6101 10115
rect 6101 10081 6135 10115
rect 6135 10081 6144 10115
rect 6092 10072 6144 10081
rect 11336 10115 11388 10124
rect 11336 10081 11345 10115
rect 11345 10081 11379 10115
rect 11379 10081 11388 10115
rect 11336 10072 11388 10081
rect 15016 10072 15068 10124
rect 8852 10047 8904 10056
rect 8852 10013 8861 10047
rect 8861 10013 8895 10047
rect 8895 10013 8904 10047
rect 8852 10004 8904 10013
rect 11060 10047 11112 10056
rect 11060 10013 11069 10047
rect 11069 10013 11103 10047
rect 11103 10013 11112 10047
rect 11060 10004 11112 10013
rect 12992 10004 13044 10056
rect 13912 10047 13964 10056
rect 13912 10013 13921 10047
rect 13921 10013 13955 10047
rect 13955 10013 13964 10047
rect 13912 10004 13964 10013
rect 16580 10072 16632 10124
rect 18604 10004 18656 10056
rect 3976 9979 4028 9988
rect 3976 9945 3985 9979
rect 3985 9945 4019 9979
rect 4019 9945 4028 9979
rect 3976 9936 4028 9945
rect 4436 9936 4488 9988
rect 3240 9911 3292 9920
rect 3240 9877 3249 9911
rect 3249 9877 3283 9911
rect 3283 9877 3292 9911
rect 3240 9868 3292 9877
rect 3424 9911 3476 9920
rect 3424 9877 3433 9911
rect 3433 9877 3467 9911
rect 3467 9877 3476 9911
rect 3424 9868 3476 9877
rect 3700 9868 3752 9920
rect 4160 9868 4212 9920
rect 5264 9868 5316 9920
rect 6828 9936 6880 9988
rect 6552 9868 6604 9920
rect 7656 9868 7708 9920
rect 11152 9979 11204 9988
rect 11152 9945 11161 9979
rect 11161 9945 11195 9979
rect 11195 9945 11204 9979
rect 11152 9936 11204 9945
rect 11612 9979 11664 9988
rect 11612 9945 11621 9979
rect 11621 9945 11655 9979
rect 11655 9945 11664 9979
rect 11612 9936 11664 9945
rect 10324 9868 10376 9920
rect 10692 9868 10744 9920
rect 14464 9936 14516 9988
rect 16764 9936 16816 9988
rect 13176 9868 13228 9920
rect 15200 9868 15252 9920
rect 18328 9911 18380 9920
rect 18328 9877 18337 9911
rect 18337 9877 18371 9911
rect 18371 9877 18380 9911
rect 18328 9868 18380 9877
rect 4660 9766 4712 9818
rect 4724 9766 4776 9818
rect 4788 9766 4840 9818
rect 4852 9766 4904 9818
rect 4916 9766 4968 9818
rect 7760 9766 7812 9818
rect 7824 9766 7876 9818
rect 7888 9766 7940 9818
rect 7952 9766 8004 9818
rect 8016 9766 8068 9818
rect 10860 9766 10912 9818
rect 10924 9766 10976 9818
rect 10988 9766 11040 9818
rect 11052 9766 11104 9818
rect 11116 9766 11168 9818
rect 13960 9766 14012 9818
rect 14024 9766 14076 9818
rect 14088 9766 14140 9818
rect 14152 9766 14204 9818
rect 14216 9766 14268 9818
rect 17060 9766 17112 9818
rect 17124 9766 17176 9818
rect 17188 9766 17240 9818
rect 17252 9766 17304 9818
rect 17316 9766 17368 9818
rect 2044 9707 2096 9716
rect 2044 9673 2053 9707
rect 2053 9673 2087 9707
rect 2087 9673 2096 9707
rect 2044 9664 2096 9673
rect 572 9639 624 9648
rect 572 9605 581 9639
rect 581 9605 615 9639
rect 615 9605 624 9639
rect 572 9596 624 9605
rect 2596 9664 2648 9716
rect 2780 9664 2832 9716
rect 3424 9664 3476 9716
rect 3700 9664 3752 9716
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 2136 9528 2188 9537
rect 2504 9571 2556 9580
rect 296 9503 348 9512
rect 296 9469 305 9503
rect 305 9469 339 9503
rect 339 9469 348 9503
rect 296 9460 348 9469
rect 2044 9460 2096 9512
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 2504 9528 2556 9537
rect 3516 9596 3568 9648
rect 2964 9571 3016 9580
rect 2964 9537 2973 9571
rect 2973 9537 3007 9571
rect 3007 9537 3016 9571
rect 2964 9528 3016 9537
rect 3700 9571 3752 9580
rect 3700 9537 3709 9571
rect 3709 9537 3743 9571
rect 3743 9537 3752 9571
rect 3700 9528 3752 9537
rect 3332 9460 3384 9512
rect 4068 9664 4120 9716
rect 7656 9664 7708 9716
rect 8576 9707 8628 9716
rect 8576 9673 8585 9707
rect 8585 9673 8619 9707
rect 8619 9673 8628 9707
rect 8576 9664 8628 9673
rect 11796 9707 11848 9716
rect 11796 9673 11805 9707
rect 11805 9673 11839 9707
rect 11839 9673 11848 9707
rect 11796 9664 11848 9673
rect 12992 9664 13044 9716
rect 14924 9664 14976 9716
rect 5172 9596 5224 9648
rect 5908 9596 5960 9648
rect 4804 9528 4856 9580
rect 5264 9528 5316 9580
rect 10324 9596 10376 9648
rect 3976 9460 4028 9512
rect 4528 9503 4580 9512
rect 4528 9469 4537 9503
rect 4537 9469 4571 9503
rect 4571 9469 4580 9503
rect 4528 9460 4580 9469
rect 5632 9503 5684 9512
rect 756 9324 808 9376
rect 3056 9392 3108 9444
rect 2596 9324 2648 9376
rect 3516 9367 3568 9376
rect 3516 9333 3525 9367
rect 3525 9333 3559 9367
rect 3559 9333 3568 9367
rect 3516 9324 3568 9333
rect 3608 9324 3660 9376
rect 5264 9367 5316 9376
rect 5264 9333 5273 9367
rect 5273 9333 5307 9367
rect 5307 9333 5316 9367
rect 5264 9324 5316 9333
rect 5632 9469 5641 9503
rect 5641 9469 5675 9503
rect 5675 9469 5684 9503
rect 5632 9460 5684 9469
rect 7196 9392 7248 9444
rect 9680 9528 9732 9580
rect 11336 9596 11388 9648
rect 11612 9596 11664 9648
rect 14372 9596 14424 9648
rect 16212 9596 16264 9648
rect 16580 9596 16632 9648
rect 10692 9571 10744 9580
rect 10692 9537 10726 9571
rect 10726 9537 10744 9571
rect 10692 9528 10744 9537
rect 7748 9503 7800 9512
rect 7748 9469 7757 9503
rect 7757 9469 7791 9503
rect 7791 9469 7800 9503
rect 7748 9460 7800 9469
rect 8116 9460 8168 9512
rect 6092 9324 6144 9376
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 7288 9324 7340 9333
rect 8944 9460 8996 9512
rect 8576 9392 8628 9444
rect 10692 9324 10744 9376
rect 13728 9528 13780 9580
rect 15292 9528 15344 9580
rect 16764 9528 16816 9580
rect 14832 9503 14884 9512
rect 14832 9469 14841 9503
rect 14841 9469 14875 9503
rect 14875 9469 14884 9503
rect 14832 9460 14884 9469
rect 15200 9503 15252 9512
rect 15200 9469 15209 9503
rect 15209 9469 15243 9503
rect 15243 9469 15252 9503
rect 15200 9460 15252 9469
rect 14372 9392 14424 9444
rect 12808 9324 12860 9376
rect 13176 9324 13228 9376
rect 13728 9324 13780 9376
rect 14464 9324 14516 9376
rect 17500 9324 17552 9376
rect 3110 9222 3162 9274
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 3302 9222 3354 9274
rect 3366 9222 3418 9274
rect 6210 9222 6262 9274
rect 6274 9222 6326 9274
rect 6338 9222 6390 9274
rect 6402 9222 6454 9274
rect 6466 9222 6518 9274
rect 9310 9222 9362 9274
rect 9374 9222 9426 9274
rect 9438 9222 9490 9274
rect 9502 9222 9554 9274
rect 9566 9222 9618 9274
rect 12410 9222 12462 9274
rect 12474 9222 12526 9274
rect 12538 9222 12590 9274
rect 12602 9222 12654 9274
rect 12666 9222 12718 9274
rect 15510 9222 15562 9274
rect 15574 9222 15626 9274
rect 15638 9222 15690 9274
rect 15702 9222 15754 9274
rect 15766 9222 15818 9274
rect 2412 9120 2464 9172
rect 2780 8984 2832 9036
rect 296 8916 348 8968
rect 756 8916 808 8968
rect 2044 8916 2096 8968
rect 2688 8959 2740 8968
rect 2688 8925 2697 8959
rect 2697 8925 2731 8959
rect 2731 8925 2740 8959
rect 2688 8916 2740 8925
rect 3700 9120 3752 9172
rect 4804 9120 4856 9172
rect 2964 8984 3016 9036
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 296 8780 348 8832
rect 664 8780 716 8832
rect 2688 8780 2740 8832
rect 4160 8984 4212 9036
rect 4804 9027 4856 9036
rect 4804 8993 4813 9027
rect 4813 8993 4847 9027
rect 4847 8993 4856 9027
rect 4804 8984 4856 8993
rect 3608 8916 3660 8968
rect 5632 9120 5684 9172
rect 5816 9052 5868 9104
rect 7748 9120 7800 9172
rect 8852 9120 8904 9172
rect 11244 9120 11296 9172
rect 12900 9120 12952 9172
rect 18328 9120 18380 9172
rect 8760 9052 8812 9104
rect 8944 9052 8996 9104
rect 6460 9027 6512 9036
rect 6460 8993 6469 9027
rect 6469 8993 6503 9027
rect 6503 8993 6512 9027
rect 6460 8984 6512 8993
rect 7288 8984 7340 9036
rect 3792 8848 3844 8900
rect 5356 8916 5408 8968
rect 7012 8959 7064 8968
rect 7012 8925 7021 8959
rect 7021 8925 7055 8959
rect 7055 8925 7064 8959
rect 7012 8916 7064 8925
rect 7196 8916 7248 8968
rect 9680 8984 9732 9036
rect 9956 8984 10008 9036
rect 10416 8984 10468 9036
rect 4988 8848 5040 8900
rect 8852 8916 8904 8968
rect 9312 8959 9364 8968
rect 9312 8925 9321 8959
rect 9321 8925 9355 8959
rect 9355 8925 9364 8959
rect 9772 8959 9824 8968
rect 9312 8916 9364 8925
rect 9772 8925 9781 8959
rect 9781 8925 9815 8959
rect 9815 8925 9824 8959
rect 9772 8916 9824 8925
rect 10324 8959 10376 8968
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 11612 8959 11664 8968
rect 11612 8925 11621 8959
rect 11621 8925 11655 8959
rect 11655 8925 11664 8959
rect 11612 8916 11664 8925
rect 3884 8780 3936 8832
rect 4528 8780 4580 8832
rect 5080 8780 5132 8832
rect 7380 8780 7432 8832
rect 10508 8848 10560 8900
rect 8852 8823 8904 8832
rect 8852 8789 8861 8823
rect 8861 8789 8895 8823
rect 8895 8789 8904 8823
rect 8852 8780 8904 8789
rect 11244 8780 11296 8832
rect 12256 8823 12308 8832
rect 12256 8789 12265 8823
rect 12265 8789 12299 8823
rect 12299 8789 12308 8823
rect 12256 8780 12308 8789
rect 12532 8780 12584 8832
rect 14740 8984 14792 9036
rect 15016 9027 15068 9036
rect 15016 8993 15025 9027
rect 15025 8993 15059 9027
rect 15059 8993 15068 9027
rect 15016 8984 15068 8993
rect 15108 8916 15160 8968
rect 13728 8848 13780 8900
rect 14648 8848 14700 8900
rect 14832 8848 14884 8900
rect 14464 8780 14516 8832
rect 14556 8780 14608 8832
rect 15016 8848 15068 8900
rect 16120 8891 16172 8900
rect 15292 8780 15344 8832
rect 16120 8857 16129 8891
rect 16129 8857 16163 8891
rect 16163 8857 16172 8891
rect 16120 8848 16172 8857
rect 16764 8848 16816 8900
rect 4660 8678 4712 8730
rect 4724 8678 4776 8730
rect 4788 8678 4840 8730
rect 4852 8678 4904 8730
rect 4916 8678 4968 8730
rect 7760 8678 7812 8730
rect 7824 8678 7876 8730
rect 7888 8678 7940 8730
rect 7952 8678 8004 8730
rect 8016 8678 8068 8730
rect 10860 8678 10912 8730
rect 10924 8678 10976 8730
rect 10988 8678 11040 8730
rect 11052 8678 11104 8730
rect 11116 8678 11168 8730
rect 13960 8678 14012 8730
rect 14024 8678 14076 8730
rect 14088 8678 14140 8730
rect 14152 8678 14204 8730
rect 14216 8678 14268 8730
rect 17060 8678 17112 8730
rect 17124 8678 17176 8730
rect 17188 8678 17240 8730
rect 17252 8678 17304 8730
rect 17316 8678 17368 8730
rect 2136 8576 2188 8628
rect 2688 8576 2740 8628
rect 4988 8576 5040 8628
rect 6552 8576 6604 8628
rect 296 8483 348 8492
rect 296 8449 305 8483
rect 305 8449 339 8483
rect 339 8449 348 8483
rect 296 8440 348 8449
rect 664 8483 716 8492
rect 664 8449 673 8483
rect 673 8449 707 8483
rect 707 8449 716 8483
rect 664 8440 716 8449
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 3884 8483 3936 8492
rect 3884 8449 3893 8483
rect 3893 8449 3927 8483
rect 3927 8449 3936 8483
rect 3884 8440 3936 8449
rect 5172 8483 5224 8492
rect 5172 8449 5181 8483
rect 5181 8449 5215 8483
rect 5215 8449 5224 8483
rect 5172 8440 5224 8449
rect 3976 8415 4028 8424
rect 3976 8381 3985 8415
rect 3985 8381 4019 8415
rect 4019 8381 4028 8415
rect 3976 8372 4028 8381
rect 5724 8508 5776 8560
rect 7380 8551 7432 8560
rect 7380 8517 7389 8551
rect 7389 8517 7423 8551
rect 7423 8517 7432 8551
rect 7380 8508 7432 8517
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 6460 8440 6512 8492
rect 7012 8440 7064 8492
rect 7656 8508 7708 8560
rect 9312 8576 9364 8628
rect 11244 8576 11296 8628
rect 12256 8576 12308 8628
rect 13728 8576 13780 8628
rect 9588 8508 9640 8560
rect 10416 8551 10468 8560
rect 10416 8517 10425 8551
rect 10425 8517 10459 8551
rect 10459 8517 10468 8551
rect 10416 8508 10468 8517
rect 11612 8508 11664 8560
rect 12900 8508 12952 8560
rect 16120 8576 16172 8628
rect 4712 8304 4764 8356
rect 5816 8372 5868 8424
rect 7196 8372 7248 8424
rect 7748 8372 7800 8424
rect 8852 8440 8904 8492
rect 9956 8483 10008 8492
rect 9956 8449 9965 8483
rect 9965 8449 9999 8483
rect 9999 8449 10008 8483
rect 9956 8440 10008 8449
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 12532 8483 12584 8492
rect 8944 8304 8996 8356
rect 10048 8304 10100 8356
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 14372 8440 14424 8492
rect 14556 8440 14608 8492
rect 16764 8508 16816 8560
rect 15292 8440 15344 8492
rect 18604 8440 18656 8492
rect 10692 8304 10744 8356
rect 13820 8372 13872 8424
rect 15108 8372 15160 8424
rect 14648 8347 14700 8356
rect 14648 8313 14657 8347
rect 14657 8313 14691 8347
rect 14691 8313 14700 8347
rect 14648 8304 14700 8313
rect 2596 8236 2648 8288
rect 2964 8279 3016 8288
rect 2964 8245 2973 8279
rect 2973 8245 3007 8279
rect 3007 8245 3016 8279
rect 2964 8236 3016 8245
rect 7656 8236 7708 8288
rect 9956 8236 10008 8288
rect 10784 8236 10836 8288
rect 16580 8236 16632 8288
rect 3110 8134 3162 8186
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 3302 8134 3354 8186
rect 3366 8134 3418 8186
rect 6210 8134 6262 8186
rect 6274 8134 6326 8186
rect 6338 8134 6390 8186
rect 6402 8134 6454 8186
rect 6466 8134 6518 8186
rect 9310 8134 9362 8186
rect 9374 8134 9426 8186
rect 9438 8134 9490 8186
rect 9502 8134 9554 8186
rect 9566 8134 9618 8186
rect 12410 8134 12462 8186
rect 12474 8134 12526 8186
rect 12538 8134 12590 8186
rect 12602 8134 12654 8186
rect 12666 8134 12718 8186
rect 15510 8134 15562 8186
rect 15574 8134 15626 8186
rect 15638 8134 15690 8186
rect 15702 8134 15754 8186
rect 15766 8134 15818 8186
rect 4252 8032 4304 8084
rect 12808 8032 12860 8084
rect 14924 8032 14976 8084
rect 2780 7964 2832 8016
rect 2412 7871 2464 7880
rect 572 7692 624 7744
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 2964 7896 3016 7948
rect 4068 7896 4120 7948
rect 5356 7964 5408 8016
rect 7196 7964 7248 8016
rect 4160 7828 4212 7880
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 2228 7692 2280 7744
rect 3056 7692 3108 7744
rect 3976 7692 4028 7744
rect 5080 7871 5132 7880
rect 5080 7837 5089 7871
rect 5089 7837 5123 7871
rect 5123 7837 5132 7871
rect 6920 7896 6972 7948
rect 8116 7896 8168 7948
rect 8392 7896 8444 7948
rect 5080 7828 5132 7837
rect 5080 7692 5132 7744
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 6092 7828 6144 7880
rect 7656 7871 7708 7880
rect 5356 7803 5408 7812
rect 5356 7769 5365 7803
rect 5365 7769 5399 7803
rect 5399 7769 5408 7803
rect 7656 7837 7665 7871
rect 7665 7837 7699 7871
rect 7699 7837 7708 7871
rect 7656 7828 7708 7837
rect 9956 7964 10008 8016
rect 9864 7871 9916 7880
rect 6828 7803 6880 7812
rect 5356 7760 5408 7769
rect 6828 7769 6837 7803
rect 6837 7769 6871 7803
rect 6871 7769 6880 7803
rect 6828 7760 6880 7769
rect 9128 7760 9180 7812
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 5632 7735 5684 7744
rect 5632 7701 5641 7735
rect 5641 7701 5675 7735
rect 5675 7701 5684 7735
rect 5632 7692 5684 7701
rect 6184 7735 6236 7744
rect 6184 7701 6193 7735
rect 6193 7701 6227 7735
rect 6227 7701 6236 7735
rect 6184 7692 6236 7701
rect 7656 7692 7708 7744
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10784 7964 10836 8016
rect 13820 7964 13872 8016
rect 13728 7896 13780 7948
rect 14464 7939 14516 7948
rect 14464 7905 14473 7939
rect 14473 7905 14507 7939
rect 14507 7905 14516 7939
rect 14464 7896 14516 7905
rect 15108 7896 15160 7948
rect 10508 7828 10560 7837
rect 12624 7828 12676 7880
rect 14740 7871 14792 7880
rect 11336 7803 11388 7812
rect 11336 7769 11345 7803
rect 11345 7769 11379 7803
rect 11379 7769 11388 7803
rect 11336 7760 11388 7769
rect 14740 7837 14749 7871
rect 14749 7837 14783 7871
rect 14783 7837 14792 7871
rect 14740 7828 14792 7837
rect 16580 7896 16632 7948
rect 17500 7939 17552 7948
rect 17500 7905 17509 7939
rect 17509 7905 17543 7939
rect 17543 7905 17552 7939
rect 17500 7896 17552 7905
rect 18052 7896 18104 7948
rect 15844 7828 15896 7880
rect 14372 7760 14424 7812
rect 10048 7692 10100 7744
rect 10416 7735 10468 7744
rect 10416 7701 10425 7735
rect 10425 7701 10459 7735
rect 10459 7701 10468 7735
rect 10416 7692 10468 7701
rect 10784 7692 10836 7744
rect 12808 7692 12860 7744
rect 14924 7692 14976 7744
rect 15292 7692 15344 7744
rect 16764 7692 16816 7744
rect 4660 7590 4712 7642
rect 4724 7590 4776 7642
rect 4788 7590 4840 7642
rect 4852 7590 4904 7642
rect 4916 7590 4968 7642
rect 7760 7590 7812 7642
rect 7824 7590 7876 7642
rect 7888 7590 7940 7642
rect 7952 7590 8004 7642
rect 8016 7590 8068 7642
rect 10860 7590 10912 7642
rect 10924 7590 10976 7642
rect 10988 7590 11040 7642
rect 11052 7590 11104 7642
rect 11116 7590 11168 7642
rect 13960 7590 14012 7642
rect 14024 7590 14076 7642
rect 14088 7590 14140 7642
rect 14152 7590 14204 7642
rect 14216 7590 14268 7642
rect 17060 7590 17112 7642
rect 17124 7590 17176 7642
rect 17188 7590 17240 7642
rect 17252 7590 17304 7642
rect 17316 7590 17368 7642
rect 2228 7531 2280 7540
rect 2228 7497 2237 7531
rect 2237 7497 2271 7531
rect 2271 7497 2280 7531
rect 2228 7488 2280 7497
rect 2412 7488 2464 7540
rect 3056 7531 3108 7540
rect 3056 7497 3065 7531
rect 3065 7497 3099 7531
rect 3099 7497 3108 7531
rect 3056 7488 3108 7497
rect 3976 7488 4028 7540
rect 572 7463 624 7472
rect 572 7429 581 7463
rect 581 7429 615 7463
rect 615 7429 624 7463
rect 572 7420 624 7429
rect 2596 7420 2648 7472
rect 2320 7395 2372 7404
rect 2320 7361 2329 7395
rect 2329 7361 2363 7395
rect 2363 7361 2372 7395
rect 2320 7352 2372 7361
rect 6184 7488 6236 7540
rect 12624 7531 12676 7540
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 13176 7488 13228 7540
rect 5908 7420 5960 7472
rect 5632 7352 5684 7404
rect 8760 7395 8812 7404
rect 8760 7361 8769 7395
rect 8769 7361 8803 7395
rect 8803 7361 8812 7395
rect 8760 7352 8812 7361
rect 3792 7284 3844 7336
rect 5080 7284 5132 7336
rect 8852 7284 8904 7336
rect 9680 7284 9732 7336
rect 11428 7420 11480 7472
rect 13563 7463 13615 7472
rect 13563 7429 13587 7463
rect 13587 7429 13615 7463
rect 13563 7420 13615 7429
rect 14556 7420 14608 7472
rect 16764 7420 16816 7472
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 11888 7352 11940 7404
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 12900 7352 12952 7361
rect 13176 7395 13228 7404
rect 13176 7361 13185 7395
rect 13185 7361 13219 7395
rect 13219 7361 13228 7395
rect 13176 7352 13228 7361
rect 13360 7395 13412 7404
rect 13360 7361 13369 7395
rect 13369 7361 13403 7395
rect 13403 7361 13412 7395
rect 13360 7352 13412 7361
rect 13452 7395 13504 7404
rect 13452 7361 13461 7395
rect 13461 7361 13495 7395
rect 13495 7361 13504 7395
rect 13452 7352 13504 7361
rect 14004 7395 14056 7404
rect 14004 7361 14013 7395
rect 14013 7361 14047 7395
rect 14047 7361 14056 7395
rect 14004 7352 14056 7361
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 16856 7352 16908 7404
rect 9956 7216 10008 7268
rect 756 7148 808 7200
rect 2596 7191 2648 7200
rect 2596 7157 2605 7191
rect 2605 7157 2639 7191
rect 2639 7157 2648 7191
rect 2596 7148 2648 7157
rect 5356 7148 5408 7200
rect 5908 7148 5960 7200
rect 8576 7191 8628 7200
rect 8576 7157 8585 7191
rect 8585 7157 8619 7191
rect 8619 7157 8628 7191
rect 8576 7148 8628 7157
rect 12808 7284 12860 7336
rect 14464 7327 14516 7336
rect 14464 7293 14473 7327
rect 14473 7293 14507 7327
rect 14507 7293 14516 7327
rect 14464 7284 14516 7293
rect 14740 7284 14792 7336
rect 13268 7259 13320 7268
rect 13268 7225 13277 7259
rect 13277 7225 13311 7259
rect 13311 7225 13320 7259
rect 13268 7216 13320 7225
rect 13636 7216 13688 7268
rect 10784 7148 10836 7200
rect 11152 7148 11204 7200
rect 11336 7148 11388 7200
rect 13728 7148 13780 7200
rect 14280 7148 14332 7200
rect 15292 7148 15344 7200
rect 16580 7148 16632 7200
rect 3110 7046 3162 7098
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 3302 7046 3354 7098
rect 3366 7046 3418 7098
rect 6210 7046 6262 7098
rect 6274 7046 6326 7098
rect 6338 7046 6390 7098
rect 6402 7046 6454 7098
rect 6466 7046 6518 7098
rect 9310 7046 9362 7098
rect 9374 7046 9426 7098
rect 9438 7046 9490 7098
rect 9502 7046 9554 7098
rect 9566 7046 9618 7098
rect 12410 7046 12462 7098
rect 12474 7046 12526 7098
rect 12538 7046 12590 7098
rect 12602 7046 12654 7098
rect 12666 7046 12718 7098
rect 15510 7046 15562 7098
rect 15574 7046 15626 7098
rect 15638 7046 15690 7098
rect 15702 7046 15754 7098
rect 15766 7046 15818 7098
rect 2780 6944 2832 6996
rect 2964 6944 3016 6996
rect 10324 6944 10376 6996
rect 14372 6987 14424 6996
rect 14372 6953 14381 6987
rect 14381 6953 14415 6987
rect 14415 6953 14424 6987
rect 14372 6944 14424 6953
rect 16672 6944 16724 6996
rect 4160 6808 4212 6860
rect 2320 6715 2372 6724
rect 2320 6681 2329 6715
rect 2329 6681 2363 6715
rect 2363 6681 2372 6715
rect 2320 6672 2372 6681
rect 2412 6672 2464 6724
rect 1952 6647 2004 6656
rect 1952 6613 1961 6647
rect 1961 6613 1995 6647
rect 1995 6613 2004 6647
rect 1952 6604 2004 6613
rect 2044 6604 2096 6656
rect 2964 6783 3016 6792
rect 2964 6749 2973 6783
rect 2973 6749 3007 6783
rect 3007 6749 3016 6783
rect 2964 6740 3016 6749
rect 3792 6740 3844 6792
rect 5448 6808 5500 6860
rect 11152 6876 11204 6928
rect 9128 6851 9180 6860
rect 6736 6672 6788 6724
rect 8208 6740 8260 6792
rect 9128 6817 9137 6851
rect 9137 6817 9171 6851
rect 9171 6817 9180 6851
rect 11520 6876 11572 6928
rect 14004 6876 14056 6928
rect 9128 6808 9180 6817
rect 13728 6808 13780 6860
rect 14464 6808 14516 6860
rect 9312 6740 9364 6792
rect 10784 6740 10836 6792
rect 11612 6740 11664 6792
rect 11888 6740 11940 6792
rect 13820 6740 13872 6792
rect 14372 6740 14424 6792
rect 14648 6740 14700 6792
rect 15292 6740 15344 6792
rect 9680 6672 9732 6724
rect 18420 6808 18472 6860
rect 15844 6783 15896 6792
rect 15844 6749 15853 6783
rect 15853 6749 15887 6783
rect 15887 6749 15896 6783
rect 15844 6740 15896 6749
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 16212 6672 16264 6724
rect 16764 6672 16816 6724
rect 17408 6672 17460 6724
rect 3884 6604 3936 6656
rect 4344 6604 4396 6656
rect 8116 6604 8168 6656
rect 8392 6604 8444 6656
rect 13636 6647 13688 6656
rect 13636 6613 13645 6647
rect 13645 6613 13679 6647
rect 13679 6613 13688 6647
rect 13636 6604 13688 6613
rect 14648 6604 14700 6656
rect 15200 6604 15252 6656
rect 15844 6604 15896 6656
rect 4660 6502 4712 6554
rect 4724 6502 4776 6554
rect 4788 6502 4840 6554
rect 4852 6502 4904 6554
rect 4916 6502 4968 6554
rect 7760 6502 7812 6554
rect 7824 6502 7876 6554
rect 7888 6502 7940 6554
rect 7952 6502 8004 6554
rect 8016 6502 8068 6554
rect 10860 6502 10912 6554
rect 10924 6502 10976 6554
rect 10988 6502 11040 6554
rect 11052 6502 11104 6554
rect 11116 6502 11168 6554
rect 13960 6502 14012 6554
rect 14024 6502 14076 6554
rect 14088 6502 14140 6554
rect 14152 6502 14204 6554
rect 14216 6502 14268 6554
rect 17060 6502 17112 6554
rect 17124 6502 17176 6554
rect 17188 6502 17240 6554
rect 17252 6502 17304 6554
rect 17316 6502 17368 6554
rect 756 6400 808 6452
rect 1860 6332 1912 6384
rect 2964 6400 3016 6452
rect 3884 6443 3936 6452
rect 3884 6409 3893 6443
rect 3893 6409 3927 6443
rect 3927 6409 3936 6443
rect 3884 6400 3936 6409
rect 5172 6400 5224 6452
rect 8576 6400 8628 6452
rect 2412 6264 2464 6316
rect 4252 6307 4304 6316
rect 4252 6273 4261 6307
rect 4261 6273 4295 6307
rect 4295 6273 4304 6307
rect 4252 6264 4304 6273
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 5816 6332 5868 6384
rect 6736 6332 6788 6384
rect 8208 6332 8260 6384
rect 11612 6400 11664 6452
rect 9956 6375 10008 6384
rect 4344 6264 4396 6273
rect 5632 6264 5684 6316
rect 8116 6307 8168 6316
rect 8116 6273 8125 6307
rect 8125 6273 8159 6307
rect 8159 6273 8168 6307
rect 8116 6264 8168 6273
rect 8484 6307 8536 6316
rect 8484 6273 8493 6307
rect 8493 6273 8527 6307
rect 8527 6273 8536 6307
rect 8484 6264 8536 6273
rect 9956 6341 9965 6375
rect 9965 6341 9999 6375
rect 9999 6341 10008 6375
rect 9956 6332 10008 6341
rect 1952 6196 2004 6248
rect 2964 6196 3016 6248
rect 940 6060 992 6112
rect 4068 6128 4120 6180
rect 5448 6239 5500 6248
rect 5448 6205 5457 6239
rect 5457 6205 5491 6239
rect 5491 6205 5500 6239
rect 5448 6196 5500 6205
rect 6920 6196 6972 6248
rect 8392 6239 8444 6248
rect 8392 6205 8401 6239
rect 8401 6205 8435 6239
rect 8435 6205 8444 6239
rect 8392 6196 8444 6205
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9680 6307 9732 6316
rect 9312 6264 9364 6273
rect 9680 6273 9689 6307
rect 9689 6273 9723 6307
rect 9723 6273 9732 6307
rect 9680 6264 9732 6273
rect 11428 6264 11480 6316
rect 12716 6400 12768 6452
rect 10692 6196 10744 6248
rect 2044 6103 2096 6112
rect 2044 6069 2053 6103
rect 2053 6069 2087 6103
rect 2087 6069 2096 6103
rect 2044 6060 2096 6069
rect 2688 6060 2740 6112
rect 7564 6060 7616 6112
rect 8944 6103 8996 6112
rect 8944 6069 8953 6103
rect 8953 6069 8987 6103
rect 8987 6069 8996 6103
rect 8944 6060 8996 6069
rect 11520 6060 11572 6112
rect 13636 6264 13688 6316
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 15108 6332 15160 6384
rect 15844 6400 15896 6452
rect 16672 6443 16724 6452
rect 16672 6409 16681 6443
rect 16681 6409 16715 6443
rect 16715 6409 16724 6443
rect 16672 6400 16724 6409
rect 16856 6443 16908 6452
rect 16856 6409 16865 6443
rect 16865 6409 16899 6443
rect 16899 6409 16908 6443
rect 16856 6400 16908 6409
rect 18052 6443 18104 6452
rect 18052 6409 18061 6443
rect 18061 6409 18095 6443
rect 18095 6409 18104 6443
rect 18052 6400 18104 6409
rect 16212 6264 16264 6316
rect 16672 6264 16724 6316
rect 11980 6196 12032 6248
rect 14372 6196 14424 6248
rect 16948 6264 17000 6316
rect 17408 6239 17460 6248
rect 17408 6205 17417 6239
rect 17417 6205 17451 6239
rect 17451 6205 17460 6239
rect 17408 6196 17460 6205
rect 17500 6196 17552 6248
rect 13728 6060 13780 6112
rect 14556 6103 14608 6112
rect 14556 6069 14565 6103
rect 14565 6069 14599 6103
rect 14599 6069 14608 6103
rect 14556 6060 14608 6069
rect 15292 6060 15344 6112
rect 3110 5958 3162 6010
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 3302 5958 3354 6010
rect 3366 5958 3418 6010
rect 6210 5958 6262 6010
rect 6274 5958 6326 6010
rect 6338 5958 6390 6010
rect 6402 5958 6454 6010
rect 6466 5958 6518 6010
rect 9310 5958 9362 6010
rect 9374 5958 9426 6010
rect 9438 5958 9490 6010
rect 9502 5958 9554 6010
rect 9566 5958 9618 6010
rect 12410 5958 12462 6010
rect 12474 5958 12526 6010
rect 12538 5958 12590 6010
rect 12602 5958 12654 6010
rect 12666 5958 12718 6010
rect 15510 5958 15562 6010
rect 15574 5958 15626 6010
rect 15638 5958 15690 6010
rect 15702 5958 15754 6010
rect 15766 5958 15818 6010
rect 2412 5899 2464 5908
rect 2412 5865 2421 5899
rect 2421 5865 2455 5899
rect 2455 5865 2464 5899
rect 2412 5856 2464 5865
rect 4252 5856 4304 5908
rect 5632 5899 5684 5908
rect 5632 5865 5641 5899
rect 5641 5865 5675 5899
rect 5675 5865 5684 5899
rect 5632 5856 5684 5865
rect 8484 5856 8536 5908
rect 2044 5788 2096 5840
rect 756 5695 808 5704
rect 756 5661 765 5695
rect 765 5661 799 5695
rect 799 5661 808 5695
rect 756 5652 808 5661
rect 2320 5695 2372 5704
rect 2320 5661 2329 5695
rect 2329 5661 2363 5695
rect 2363 5661 2372 5695
rect 2320 5652 2372 5661
rect 3056 5652 3108 5704
rect 4068 5788 4120 5840
rect 4068 5652 4120 5704
rect 3884 5584 3936 5636
rect 6828 5652 6880 5704
rect 7472 5652 7524 5704
rect 7564 5695 7616 5704
rect 7564 5661 7573 5695
rect 7573 5661 7607 5695
rect 7607 5661 7616 5695
rect 7564 5652 7616 5661
rect 15384 5856 15436 5908
rect 16948 5856 17000 5908
rect 11244 5788 11296 5840
rect 11980 5831 12032 5840
rect 11980 5797 11989 5831
rect 11989 5797 12023 5831
rect 12023 5797 12032 5831
rect 11980 5788 12032 5797
rect 5172 5627 5224 5636
rect 5172 5593 5181 5627
rect 5181 5593 5215 5627
rect 5215 5593 5224 5627
rect 5172 5584 5224 5593
rect 8668 5627 8720 5636
rect 8668 5593 8677 5627
rect 8677 5593 8711 5627
rect 8711 5593 8720 5627
rect 8668 5584 8720 5593
rect 480 5516 532 5568
rect 2412 5516 2464 5568
rect 2872 5516 2924 5568
rect 3976 5559 4028 5568
rect 3976 5525 3985 5559
rect 3985 5525 4019 5559
rect 4019 5525 4028 5559
rect 3976 5516 4028 5525
rect 5264 5559 5316 5568
rect 5264 5525 5273 5559
rect 5273 5525 5307 5559
rect 5307 5525 5316 5559
rect 5264 5516 5316 5525
rect 9036 5516 9088 5568
rect 10784 5516 10836 5568
rect 12900 5720 12952 5772
rect 13728 5763 13780 5772
rect 13728 5729 13737 5763
rect 13737 5729 13771 5763
rect 13771 5729 13780 5763
rect 13728 5720 13780 5729
rect 13636 5652 13688 5704
rect 14372 5720 14424 5772
rect 15292 5763 15344 5772
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 16580 5720 16632 5772
rect 14464 5652 14516 5704
rect 15384 5652 15436 5704
rect 18512 5695 18564 5704
rect 18512 5661 18521 5695
rect 18521 5661 18555 5695
rect 18555 5661 18564 5695
rect 18512 5652 18564 5661
rect 13636 5516 13688 5568
rect 15016 5559 15068 5568
rect 15016 5525 15025 5559
rect 15025 5525 15059 5559
rect 15059 5525 15068 5559
rect 15016 5516 15068 5525
rect 15660 5516 15712 5568
rect 16672 5516 16724 5568
rect 18328 5559 18380 5568
rect 18328 5525 18337 5559
rect 18337 5525 18371 5559
rect 18371 5525 18380 5559
rect 18328 5516 18380 5525
rect 4660 5414 4712 5466
rect 4724 5414 4776 5466
rect 4788 5414 4840 5466
rect 4852 5414 4904 5466
rect 4916 5414 4968 5466
rect 7760 5414 7812 5466
rect 7824 5414 7876 5466
rect 7888 5414 7940 5466
rect 7952 5414 8004 5466
rect 8016 5414 8068 5466
rect 10860 5414 10912 5466
rect 10924 5414 10976 5466
rect 10988 5414 11040 5466
rect 11052 5414 11104 5466
rect 11116 5414 11168 5466
rect 13960 5414 14012 5466
rect 14024 5414 14076 5466
rect 14088 5414 14140 5466
rect 14152 5414 14204 5466
rect 14216 5414 14268 5466
rect 17060 5414 17112 5466
rect 17124 5414 17176 5466
rect 17188 5414 17240 5466
rect 17252 5414 17304 5466
rect 17316 5414 17368 5466
rect 2320 5312 2372 5364
rect 5264 5312 5316 5364
rect 1860 5244 1912 5296
rect 2596 5244 2648 5296
rect 7656 5244 7708 5296
rect 8944 5244 8996 5296
rect 480 5219 532 5228
rect 480 5185 489 5219
rect 489 5185 523 5219
rect 523 5185 532 5219
rect 480 5176 532 5185
rect 940 5176 992 5228
rect 4068 5219 4120 5228
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 4068 5176 4120 5185
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 9036 5219 9088 5228
rect 3056 5108 3108 5160
rect 3884 5108 3936 5160
rect 9036 5185 9045 5219
rect 9045 5185 9079 5219
rect 9079 5185 9088 5219
rect 9036 5176 9088 5185
rect 10784 5312 10836 5364
rect 8852 5040 8904 5092
rect 2596 5015 2648 5024
rect 2596 4981 2605 5015
rect 2605 4981 2639 5015
rect 2639 4981 2648 5015
rect 2596 4972 2648 4981
rect 9220 4972 9272 5024
rect 13820 5176 13872 5228
rect 11152 5108 11204 5160
rect 13636 5108 13688 5160
rect 9956 4972 10008 5024
rect 11244 4972 11296 5024
rect 11520 4972 11572 5024
rect 13820 5015 13872 5024
rect 13820 4981 13829 5015
rect 13829 4981 13863 5015
rect 13863 4981 13872 5015
rect 13820 4972 13872 4981
rect 14556 4972 14608 5024
rect 15660 5244 15712 5296
rect 17500 5244 17552 5296
rect 14924 5219 14976 5228
rect 14924 5185 14933 5219
rect 14933 5185 14967 5219
rect 14967 5185 14976 5219
rect 14924 5176 14976 5185
rect 16948 5219 17000 5228
rect 16948 5185 16957 5219
rect 16957 5185 16991 5219
rect 16991 5185 17000 5219
rect 16948 5176 17000 5185
rect 18328 5108 18380 5160
rect 16856 4972 16908 5024
rect 3110 4870 3162 4922
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 3302 4870 3354 4922
rect 3366 4870 3418 4922
rect 6210 4870 6262 4922
rect 6274 4870 6326 4922
rect 6338 4870 6390 4922
rect 6402 4870 6454 4922
rect 6466 4870 6518 4922
rect 9310 4870 9362 4922
rect 9374 4870 9426 4922
rect 9438 4870 9490 4922
rect 9502 4870 9554 4922
rect 9566 4870 9618 4922
rect 12410 4870 12462 4922
rect 12474 4870 12526 4922
rect 12538 4870 12590 4922
rect 12602 4870 12654 4922
rect 12666 4870 12718 4922
rect 15510 4870 15562 4922
rect 15574 4870 15626 4922
rect 15638 4870 15690 4922
rect 15702 4870 15754 4922
rect 15766 4870 15818 4922
rect 11152 4811 11204 4820
rect 11152 4777 11161 4811
rect 11161 4777 11195 4811
rect 11195 4777 11204 4811
rect 11152 4768 11204 4777
rect 13912 4768 13964 4820
rect 2964 4632 3016 4684
rect 6920 4632 6972 4684
rect 9956 4632 10008 4684
rect 6460 4607 6512 4616
rect 6460 4573 6469 4607
rect 6469 4573 6503 4607
rect 6503 4573 6512 4607
rect 6460 4564 6512 4573
rect 7656 4564 7708 4616
rect 11520 4607 11572 4616
rect 11520 4573 11529 4607
rect 11529 4573 11563 4607
rect 11563 4573 11572 4607
rect 13820 4632 13872 4684
rect 15476 4675 15528 4684
rect 15476 4641 15485 4675
rect 15485 4641 15519 4675
rect 15519 4641 15528 4675
rect 15476 4632 15528 4641
rect 16856 4632 16908 4684
rect 11520 4564 11572 4573
rect 3516 4496 3568 4548
rect 480 4428 532 4480
rect 2596 4428 2648 4480
rect 5448 4471 5500 4480
rect 5448 4437 5457 4471
rect 5457 4437 5491 4471
rect 5491 4437 5500 4471
rect 5448 4428 5500 4437
rect 8392 4496 8444 4548
rect 8576 4428 8628 4480
rect 8852 4496 8904 4548
rect 9220 4496 9272 4548
rect 11612 4496 11664 4548
rect 9772 4428 9824 4480
rect 17868 4607 17920 4616
rect 17868 4573 17877 4607
rect 17877 4573 17911 4607
rect 17911 4573 17920 4607
rect 17868 4564 17920 4573
rect 11980 4496 12032 4548
rect 12256 4471 12308 4480
rect 12256 4437 12265 4471
rect 12265 4437 12299 4471
rect 12299 4437 12308 4471
rect 12256 4428 12308 4437
rect 13176 4428 13228 4480
rect 15200 4496 15252 4548
rect 14556 4428 14608 4480
rect 4660 4326 4712 4378
rect 4724 4326 4776 4378
rect 4788 4326 4840 4378
rect 4852 4326 4904 4378
rect 4916 4326 4968 4378
rect 7760 4326 7812 4378
rect 7824 4326 7876 4378
rect 7888 4326 7940 4378
rect 7952 4326 8004 4378
rect 8016 4326 8068 4378
rect 10860 4326 10912 4378
rect 10924 4326 10976 4378
rect 10988 4326 11040 4378
rect 11052 4326 11104 4378
rect 11116 4326 11168 4378
rect 13960 4326 14012 4378
rect 14024 4326 14076 4378
rect 14088 4326 14140 4378
rect 14152 4326 14204 4378
rect 14216 4326 14268 4378
rect 17060 4326 17112 4378
rect 17124 4326 17176 4378
rect 17188 4326 17240 4378
rect 17252 4326 17304 4378
rect 17316 4326 17368 4378
rect 2412 4224 2464 4276
rect 3516 4267 3568 4276
rect 3516 4233 3525 4267
rect 3525 4233 3559 4267
rect 3559 4233 3568 4267
rect 3516 4224 3568 4233
rect 4344 4224 4396 4276
rect 6460 4224 6512 4276
rect 2596 4156 2648 4208
rect 480 4131 532 4140
rect 480 4097 489 4131
rect 489 4097 523 4131
rect 523 4097 532 4131
rect 480 4088 532 4097
rect 2412 4020 2464 4072
rect 2872 4156 2924 4208
rect 3056 4131 3108 4140
rect 3056 4097 3065 4131
rect 3065 4097 3099 4131
rect 3099 4097 3108 4131
rect 3056 4088 3108 4097
rect 3792 4131 3844 4140
rect 3792 4097 3801 4131
rect 3801 4097 3835 4131
rect 3835 4097 3844 4131
rect 3792 4088 3844 4097
rect 4344 4131 4396 4140
rect 4344 4097 4353 4131
rect 4353 4097 4387 4131
rect 4387 4097 4396 4131
rect 4988 4131 5040 4140
rect 4344 4088 4396 4097
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 8668 4156 8720 4208
rect 8852 4224 8904 4276
rect 14740 4224 14792 4276
rect 5448 4088 5500 4140
rect 2780 3884 2832 3936
rect 6920 3952 6972 4004
rect 7656 4088 7708 4140
rect 8576 4131 8628 4140
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 7564 4020 7616 4072
rect 3516 3884 3568 3936
rect 4620 3884 4672 3936
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 10048 4088 10100 4140
rect 9772 4020 9824 4072
rect 10784 4088 10836 4140
rect 11244 4156 11296 4208
rect 12164 4156 12216 4208
rect 11428 4088 11480 4140
rect 11612 4131 11664 4140
rect 11612 4097 11621 4131
rect 11621 4097 11655 4131
rect 11655 4097 11664 4131
rect 11612 4088 11664 4097
rect 10968 4063 11020 4072
rect 9956 3952 10008 4004
rect 10968 4029 10977 4063
rect 10977 4029 11011 4063
rect 11011 4029 11020 4063
rect 10968 4020 11020 4029
rect 11796 4088 11848 4140
rect 12256 4131 12308 4140
rect 12256 4097 12265 4131
rect 12265 4097 12299 4131
rect 12299 4097 12308 4131
rect 12256 4088 12308 4097
rect 13176 4156 13228 4208
rect 14556 4199 14608 4208
rect 14556 4165 14565 4199
rect 14565 4165 14599 4199
rect 14599 4165 14608 4199
rect 14556 4156 14608 4165
rect 12808 4063 12860 4072
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 12808 4020 12860 4029
rect 18512 4131 18564 4140
rect 18512 4097 18521 4131
rect 18521 4097 18555 4131
rect 18555 4097 18564 4131
rect 18512 4088 18564 4097
rect 13820 4020 13872 4072
rect 14832 4020 14884 4072
rect 15476 4020 15528 4072
rect 11888 3927 11940 3936
rect 11888 3893 11897 3927
rect 11897 3893 11931 3927
rect 11931 3893 11940 3927
rect 11888 3884 11940 3893
rect 13728 3884 13780 3936
rect 17776 3884 17828 3936
rect 18328 3927 18380 3936
rect 18328 3893 18337 3927
rect 18337 3893 18371 3927
rect 18371 3893 18380 3927
rect 18328 3884 18380 3893
rect 3110 3782 3162 3834
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 3302 3782 3354 3834
rect 3366 3782 3418 3834
rect 6210 3782 6262 3834
rect 6274 3782 6326 3834
rect 6338 3782 6390 3834
rect 6402 3782 6454 3834
rect 6466 3782 6518 3834
rect 9310 3782 9362 3834
rect 9374 3782 9426 3834
rect 9438 3782 9490 3834
rect 9502 3782 9554 3834
rect 9566 3782 9618 3834
rect 12410 3782 12462 3834
rect 12474 3782 12526 3834
rect 12538 3782 12590 3834
rect 12602 3782 12654 3834
rect 12666 3782 12718 3834
rect 15510 3782 15562 3834
rect 15574 3782 15626 3834
rect 15638 3782 15690 3834
rect 15702 3782 15754 3834
rect 15766 3782 15818 3834
rect 2780 3723 2832 3732
rect 2780 3689 2789 3723
rect 2789 3689 2823 3723
rect 2823 3689 2832 3723
rect 2780 3680 2832 3689
rect 9956 3680 10008 3732
rect 10968 3680 11020 3732
rect 12808 3680 12860 3732
rect 14740 3680 14792 3732
rect 2688 3655 2740 3664
rect 2688 3621 2697 3655
rect 2697 3621 2731 3655
rect 2731 3621 2740 3655
rect 2688 3612 2740 3621
rect 5632 3612 5684 3664
rect 3792 3544 3844 3596
rect 2596 3476 2648 3528
rect 3148 3519 3200 3528
rect 3148 3485 3157 3519
rect 3157 3485 3191 3519
rect 3191 3485 3200 3519
rect 3148 3476 3200 3485
rect 4252 3544 4304 3596
rect 4988 3544 5040 3596
rect 7564 3612 7616 3664
rect 7656 3612 7708 3664
rect 6736 3544 6788 3596
rect 11612 3612 11664 3664
rect 14924 3612 14976 3664
rect 2320 3451 2372 3460
rect 2320 3417 2329 3451
rect 2329 3417 2363 3451
rect 2363 3417 2372 3451
rect 2320 3408 2372 3417
rect 572 3340 624 3392
rect 2872 3340 2924 3392
rect 4068 3519 4120 3528
rect 4068 3485 4077 3519
rect 4077 3485 4111 3519
rect 4111 3485 4120 3519
rect 4068 3476 4120 3485
rect 4620 3476 4672 3528
rect 5448 3408 5500 3460
rect 6644 3476 6696 3528
rect 11888 3544 11940 3596
rect 13636 3544 13688 3596
rect 14648 3544 14700 3596
rect 9772 3519 9824 3528
rect 7380 3408 7432 3460
rect 7564 3408 7616 3460
rect 8208 3408 8260 3460
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 9772 3476 9824 3485
rect 13728 3476 13780 3528
rect 13820 3476 13872 3528
rect 15292 3476 15344 3528
rect 15752 3519 15804 3528
rect 15752 3485 15761 3519
rect 15761 3485 15795 3519
rect 15795 3485 15804 3519
rect 15752 3476 15804 3485
rect 15844 3476 15896 3528
rect 18144 3476 18196 3528
rect 4160 3340 4212 3392
rect 5724 3340 5776 3392
rect 6000 3340 6052 3392
rect 6552 3340 6604 3392
rect 6644 3340 6696 3392
rect 10784 3408 10836 3460
rect 11428 3408 11480 3460
rect 11980 3408 12032 3460
rect 13636 3408 13688 3460
rect 8392 3340 8444 3392
rect 9036 3340 9088 3392
rect 11336 3340 11388 3392
rect 13176 3340 13228 3392
rect 14372 3383 14424 3392
rect 14372 3349 14381 3383
rect 14381 3349 14415 3383
rect 14415 3349 14424 3383
rect 14372 3340 14424 3349
rect 15108 3340 15160 3392
rect 4660 3238 4712 3290
rect 4724 3238 4776 3290
rect 4788 3238 4840 3290
rect 4852 3238 4904 3290
rect 4916 3238 4968 3290
rect 7760 3238 7812 3290
rect 7824 3238 7876 3290
rect 7888 3238 7940 3290
rect 7952 3238 8004 3290
rect 8016 3238 8068 3290
rect 10860 3238 10912 3290
rect 10924 3238 10976 3290
rect 10988 3238 11040 3290
rect 11052 3238 11104 3290
rect 11116 3238 11168 3290
rect 13960 3238 14012 3290
rect 14024 3238 14076 3290
rect 14088 3238 14140 3290
rect 14152 3238 14204 3290
rect 14216 3238 14268 3290
rect 17060 3238 17112 3290
rect 17124 3238 17176 3290
rect 17188 3238 17240 3290
rect 17252 3238 17304 3290
rect 17316 3238 17368 3290
rect 2596 3179 2648 3188
rect 572 3111 624 3120
rect 572 3077 581 3111
rect 581 3077 615 3111
rect 615 3077 624 3111
rect 572 3068 624 3077
rect 2596 3145 2605 3179
rect 2605 3145 2639 3179
rect 2639 3145 2648 3179
rect 2596 3136 2648 3145
rect 3148 3179 3200 3188
rect 3148 3145 3157 3179
rect 3157 3145 3191 3179
rect 3191 3145 3200 3179
rect 3148 3136 3200 3145
rect 2320 3068 2372 3120
rect 4068 3136 4120 3188
rect 5448 3179 5500 3188
rect 5448 3145 5457 3179
rect 5457 3145 5491 3179
rect 5491 3145 5500 3179
rect 5448 3136 5500 3145
rect 5724 3136 5776 3188
rect 9036 3136 9088 3188
rect 2688 3043 2740 3052
rect 296 2975 348 2984
rect 296 2941 305 2975
rect 305 2941 339 2975
rect 339 2941 348 2975
rect 296 2932 348 2941
rect 2688 3009 2697 3043
rect 2697 3009 2731 3043
rect 2731 3009 2740 3043
rect 2688 3000 2740 3009
rect 3700 3043 3752 3052
rect 3700 3009 3709 3043
rect 3709 3009 3743 3043
rect 3743 3009 3752 3043
rect 3700 3000 3752 3009
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 4252 3043 4304 3052
rect 4252 3009 4261 3043
rect 4261 3009 4295 3043
rect 4295 3009 4304 3043
rect 6552 3068 6604 3120
rect 7104 3068 7156 3120
rect 9220 3068 9272 3120
rect 9864 3068 9916 3120
rect 11336 3136 11388 3188
rect 4252 3000 4304 3009
rect 3516 2932 3568 2984
rect 7288 3000 7340 3052
rect 7656 3043 7708 3052
rect 7656 3009 7665 3043
rect 7665 3009 7699 3043
rect 7699 3009 7708 3043
rect 7656 3000 7708 3009
rect 7748 3043 7800 3052
rect 7748 3009 7757 3043
rect 7757 3009 7791 3043
rect 7791 3009 7800 3043
rect 8208 3043 8260 3052
rect 7748 3000 7800 3009
rect 8208 3009 8217 3043
rect 8217 3009 8251 3043
rect 8251 3009 8260 3043
rect 8208 3000 8260 3009
rect 6000 2975 6052 2984
rect 6000 2941 6009 2975
rect 6009 2941 6043 2975
rect 6043 2941 6052 2975
rect 6000 2932 6052 2941
rect 7472 2932 7524 2984
rect 7104 2864 7156 2916
rect 9128 2864 9180 2916
rect 2504 2796 2556 2848
rect 3792 2839 3844 2848
rect 3792 2805 3801 2839
rect 3801 2805 3835 2839
rect 3835 2805 3844 2839
rect 3792 2796 3844 2805
rect 4344 2796 4396 2848
rect 7196 2796 7248 2848
rect 8852 2796 8904 2848
rect 9036 2796 9088 2848
rect 12992 3136 13044 3188
rect 14648 3179 14700 3188
rect 14648 3145 14657 3179
rect 14657 3145 14691 3179
rect 14691 3145 14700 3179
rect 14648 3136 14700 3145
rect 15844 3136 15896 3188
rect 15108 3068 15160 3120
rect 12808 3000 12860 3052
rect 13544 3043 13596 3052
rect 13544 3009 13553 3043
rect 13553 3009 13587 3043
rect 13587 3009 13596 3043
rect 13544 3000 13596 3009
rect 10324 2796 10376 2848
rect 14372 3000 14424 3052
rect 14556 3043 14608 3052
rect 14556 3009 14565 3043
rect 14565 3009 14599 3043
rect 14599 3009 14608 3043
rect 14556 3000 14608 3009
rect 14740 3043 14792 3052
rect 14740 3009 14749 3043
rect 14749 3009 14783 3043
rect 14783 3009 14792 3043
rect 14740 3000 14792 3009
rect 15384 3000 15436 3052
rect 18328 3000 18380 3052
rect 14924 2932 14976 2984
rect 15108 2932 15160 2984
rect 15844 2932 15896 2984
rect 17868 2932 17920 2984
rect 3110 2694 3162 2746
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 3302 2694 3354 2746
rect 3366 2694 3418 2746
rect 6210 2694 6262 2746
rect 6274 2694 6326 2746
rect 6338 2694 6390 2746
rect 6402 2694 6454 2746
rect 6466 2694 6518 2746
rect 9310 2694 9362 2746
rect 9374 2694 9426 2746
rect 9438 2694 9490 2746
rect 9502 2694 9554 2746
rect 9566 2694 9618 2746
rect 12410 2694 12462 2746
rect 12474 2694 12526 2746
rect 12538 2694 12590 2746
rect 12602 2694 12654 2746
rect 12666 2694 12718 2746
rect 15510 2694 15562 2746
rect 15574 2694 15626 2746
rect 15638 2694 15690 2746
rect 15702 2694 15754 2746
rect 15766 2694 15818 2746
rect 3516 2592 3568 2644
rect 3792 2524 3844 2576
rect 3700 2499 3752 2508
rect 3700 2465 3709 2499
rect 3709 2465 3743 2499
rect 3743 2465 3752 2499
rect 3700 2456 3752 2465
rect 7472 2592 7524 2644
rect 7656 2592 7708 2644
rect 10324 2592 10376 2644
rect 7748 2524 7800 2576
rect 5448 2456 5500 2508
rect 7012 2456 7064 2508
rect 8852 2499 8904 2508
rect 5540 2388 5592 2440
rect 6552 2388 6604 2440
rect 7104 2431 7156 2440
rect 5632 2320 5684 2372
rect 6828 2363 6880 2372
rect 6828 2329 6837 2363
rect 6837 2329 6871 2363
rect 6871 2329 6880 2363
rect 6828 2320 6880 2329
rect 848 2252 900 2304
rect 3792 2252 3844 2304
rect 5264 2252 5316 2304
rect 7104 2397 7113 2431
rect 7113 2397 7147 2431
rect 7147 2397 7156 2431
rect 7104 2388 7156 2397
rect 7196 2388 7248 2440
rect 8852 2465 8861 2499
rect 8861 2465 8895 2499
rect 8895 2465 8904 2499
rect 8852 2456 8904 2465
rect 9128 2456 9180 2508
rect 8944 2388 8996 2440
rect 7012 2320 7064 2372
rect 7472 2363 7524 2372
rect 7472 2329 7481 2363
rect 7481 2329 7515 2363
rect 7515 2329 7524 2363
rect 7472 2320 7524 2329
rect 9220 2320 9272 2372
rect 10600 2320 10652 2372
rect 10784 2320 10836 2372
rect 14556 2592 14608 2644
rect 15200 2592 15252 2644
rect 11888 2524 11940 2576
rect 12900 2524 12952 2576
rect 12992 2567 13044 2576
rect 12992 2533 13001 2567
rect 13001 2533 13035 2567
rect 13035 2533 13044 2567
rect 12992 2524 13044 2533
rect 11520 2499 11572 2508
rect 11520 2465 11529 2499
rect 11529 2465 11563 2499
rect 11563 2465 11572 2499
rect 11520 2456 11572 2465
rect 12256 2456 12308 2508
rect 12348 2431 12400 2440
rect 12348 2397 12357 2431
rect 12357 2397 12391 2431
rect 12391 2397 12400 2431
rect 12348 2388 12400 2397
rect 13820 2499 13872 2508
rect 13820 2465 13829 2499
rect 13829 2465 13863 2499
rect 13863 2465 13872 2499
rect 13820 2456 13872 2465
rect 16948 2456 17000 2508
rect 17868 2499 17920 2508
rect 17868 2465 17877 2499
rect 17877 2465 17911 2499
rect 17911 2465 17920 2499
rect 17868 2456 17920 2465
rect 12624 2388 12676 2440
rect 11612 2320 11664 2372
rect 7380 2252 7432 2304
rect 7656 2252 7708 2304
rect 8760 2252 8812 2304
rect 11244 2295 11296 2304
rect 11244 2261 11253 2295
rect 11253 2261 11287 2295
rect 11287 2261 11296 2295
rect 11244 2252 11296 2261
rect 11980 2252 12032 2304
rect 12348 2252 12400 2304
rect 13636 2388 13688 2440
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 13176 2320 13228 2372
rect 14556 2320 14608 2372
rect 17592 2363 17644 2372
rect 14648 2252 14700 2304
rect 15384 2295 15436 2304
rect 15384 2261 15393 2295
rect 15393 2261 15427 2295
rect 15427 2261 15436 2295
rect 17592 2329 17601 2363
rect 17601 2329 17635 2363
rect 17635 2329 17644 2363
rect 17592 2320 17644 2329
rect 15384 2252 15436 2261
rect 16120 2252 16172 2304
rect 4660 2150 4712 2202
rect 4724 2150 4776 2202
rect 4788 2150 4840 2202
rect 4852 2150 4904 2202
rect 4916 2150 4968 2202
rect 7760 2150 7812 2202
rect 7824 2150 7876 2202
rect 7888 2150 7940 2202
rect 7952 2150 8004 2202
rect 8016 2150 8068 2202
rect 10860 2150 10912 2202
rect 10924 2150 10976 2202
rect 10988 2150 11040 2202
rect 11052 2150 11104 2202
rect 11116 2150 11168 2202
rect 13960 2150 14012 2202
rect 14024 2150 14076 2202
rect 14088 2150 14140 2202
rect 14152 2150 14204 2202
rect 14216 2150 14268 2202
rect 17060 2150 17112 2202
rect 17124 2150 17176 2202
rect 17188 2150 17240 2202
rect 17252 2150 17304 2202
rect 17316 2150 17368 2202
rect 1216 2048 1268 2100
rect 2964 2048 3016 2100
rect 3792 2091 3844 2100
rect 848 2023 900 2032
rect 848 1989 857 2023
rect 857 1989 891 2023
rect 891 1989 900 2023
rect 848 1980 900 1989
rect 296 1844 348 1896
rect 1216 1844 1268 1896
rect 2780 1980 2832 2032
rect 2964 1912 3016 1964
rect 3792 2057 3801 2091
rect 3801 2057 3835 2091
rect 3835 2057 3844 2091
rect 3792 2048 3844 2057
rect 4344 2048 4396 2100
rect 5264 2091 5316 2100
rect 5264 2057 5273 2091
rect 5273 2057 5307 2091
rect 5307 2057 5316 2091
rect 5264 2048 5316 2057
rect 5632 2048 5684 2100
rect 6644 2048 6696 2100
rect 6828 2048 6880 2100
rect 7288 2048 7340 2100
rect 10600 2091 10652 2100
rect 3516 1980 3568 2032
rect 7104 1980 7156 2032
rect 7656 1980 7708 2032
rect 10600 2057 10609 2091
rect 10609 2057 10643 2091
rect 10643 2057 10652 2091
rect 10600 2048 10652 2057
rect 11244 2048 11296 2100
rect 12624 2091 12676 2100
rect 12624 2057 12633 2091
rect 12633 2057 12667 2091
rect 12667 2057 12676 2091
rect 12624 2048 12676 2057
rect 14556 2048 14608 2100
rect 3884 1955 3936 1964
rect 2596 1776 2648 1828
rect 3884 1921 3893 1955
rect 3893 1921 3927 1955
rect 3927 1921 3936 1955
rect 3884 1912 3936 1921
rect 5908 1912 5960 1964
rect 6920 1912 6972 1964
rect 7288 1955 7340 1964
rect 7288 1921 7297 1955
rect 7297 1921 7331 1955
rect 7331 1921 7340 1955
rect 7288 1912 7340 1921
rect 9036 1912 9088 1964
rect 9312 1912 9364 1964
rect 9588 1912 9640 1964
rect 11980 1980 12032 2032
rect 5724 1844 5776 1896
rect 6000 1844 6052 1896
rect 6552 1844 6604 1896
rect 7012 1844 7064 1896
rect 8300 1844 8352 1896
rect 9956 1887 10008 1896
rect 9956 1853 9965 1887
rect 9965 1853 9999 1887
rect 9999 1853 10008 1887
rect 9956 1844 10008 1853
rect 12808 1912 12860 1964
rect 6092 1776 6144 1828
rect 12256 1844 12308 1896
rect 14464 1955 14516 1964
rect 14464 1921 14473 1955
rect 14473 1921 14507 1955
rect 14507 1921 14516 1955
rect 14464 1912 14516 1921
rect 14648 1955 14700 1964
rect 14648 1921 14657 1955
rect 14657 1921 14691 1955
rect 14691 1921 14700 1955
rect 14648 1912 14700 1921
rect 16948 2048 17000 2100
rect 14924 1955 14976 1964
rect 14924 1921 14933 1955
rect 14933 1921 14967 1955
rect 14967 1921 14976 1955
rect 15292 1955 15344 1964
rect 14924 1912 14976 1921
rect 15292 1921 15301 1955
rect 15301 1921 15335 1955
rect 15335 1921 15344 1955
rect 15292 1912 15344 1921
rect 15200 1887 15252 1896
rect 15200 1853 15209 1887
rect 15209 1853 15243 1887
rect 15243 1853 15252 1887
rect 15200 1844 15252 1853
rect 16488 1912 16540 1964
rect 10784 1776 10836 1828
rect 2504 1751 2556 1760
rect 2504 1717 2513 1751
rect 2513 1717 2547 1751
rect 2547 1717 2556 1751
rect 2504 1708 2556 1717
rect 2872 1751 2924 1760
rect 2872 1717 2881 1751
rect 2881 1717 2915 1751
rect 2915 1717 2924 1751
rect 2872 1708 2924 1717
rect 3516 1708 3568 1760
rect 6828 1751 6880 1760
rect 6828 1717 6837 1751
rect 6837 1717 6871 1751
rect 6871 1717 6880 1751
rect 6828 1708 6880 1717
rect 7104 1751 7156 1760
rect 7104 1717 7113 1751
rect 7113 1717 7147 1751
rect 7147 1717 7156 1751
rect 7104 1708 7156 1717
rect 9128 1751 9180 1760
rect 9128 1717 9137 1751
rect 9137 1717 9171 1751
rect 9171 1717 9180 1751
rect 9128 1708 9180 1717
rect 11152 1708 11204 1760
rect 14648 1776 14700 1828
rect 15108 1819 15160 1828
rect 15108 1785 15117 1819
rect 15117 1785 15151 1819
rect 15151 1785 15160 1819
rect 15108 1776 15160 1785
rect 12992 1708 13044 1760
rect 14188 1751 14240 1760
rect 14188 1717 14197 1751
rect 14197 1717 14231 1751
rect 14231 1717 14240 1751
rect 16672 1751 16724 1760
rect 14188 1708 14240 1717
rect 16672 1717 16681 1751
rect 16681 1717 16715 1751
rect 16715 1717 16724 1751
rect 16672 1708 16724 1717
rect 3110 1606 3162 1658
rect 3174 1606 3226 1658
rect 3238 1606 3290 1658
rect 3302 1606 3354 1658
rect 3366 1606 3418 1658
rect 6210 1606 6262 1658
rect 6274 1606 6326 1658
rect 6338 1606 6390 1658
rect 6402 1606 6454 1658
rect 6466 1606 6518 1658
rect 9310 1606 9362 1658
rect 9374 1606 9426 1658
rect 9438 1606 9490 1658
rect 9502 1606 9554 1658
rect 9566 1606 9618 1658
rect 12410 1606 12462 1658
rect 12474 1606 12526 1658
rect 12538 1606 12590 1658
rect 12602 1606 12654 1658
rect 12666 1606 12718 1658
rect 15510 1606 15562 1658
rect 15574 1606 15626 1658
rect 15638 1606 15690 1658
rect 15702 1606 15754 1658
rect 15766 1606 15818 1658
rect 2964 1504 3016 1556
rect 3700 1504 3752 1556
rect 5908 1547 5960 1556
rect 5908 1513 5917 1547
rect 5917 1513 5951 1547
rect 5951 1513 5960 1547
rect 5908 1504 5960 1513
rect 6092 1547 6144 1556
rect 6092 1513 6101 1547
rect 6101 1513 6135 1547
rect 6135 1513 6144 1547
rect 6092 1504 6144 1513
rect 9956 1504 10008 1556
rect 11980 1504 12032 1556
rect 14188 1504 14240 1556
rect 17592 1547 17644 1556
rect 17592 1513 17601 1547
rect 17601 1513 17635 1547
rect 17635 1513 17644 1547
rect 17592 1504 17644 1513
rect 2780 1436 2832 1488
rect 3884 1436 3936 1488
rect 1216 1368 1268 1420
rect 2872 1368 2924 1420
rect 5632 1411 5684 1420
rect 3700 1300 3752 1352
rect 5632 1377 5641 1411
rect 5641 1377 5675 1411
rect 5675 1377 5684 1411
rect 5632 1368 5684 1377
rect 6000 1368 6052 1420
rect 7380 1368 7432 1420
rect 9128 1411 9180 1420
rect 9128 1377 9137 1411
rect 9137 1377 9171 1411
rect 9171 1377 9180 1411
rect 9128 1368 9180 1377
rect 4988 1300 5040 1352
rect 6828 1300 6880 1352
rect 8300 1300 8352 1352
rect 8668 1343 8720 1352
rect 8668 1309 8677 1343
rect 8677 1309 8711 1343
rect 8711 1309 8720 1343
rect 8668 1300 8720 1309
rect 8760 1343 8812 1352
rect 8760 1309 8769 1343
rect 8769 1309 8803 1343
rect 8803 1309 8812 1343
rect 8760 1300 8812 1309
rect 10048 1300 10100 1352
rect 2504 1164 2556 1216
rect 2872 1232 2924 1284
rect 3332 1232 3384 1284
rect 6644 1232 6696 1284
rect 10140 1232 10192 1284
rect 10416 1343 10468 1352
rect 10416 1309 10425 1343
rect 10425 1309 10459 1343
rect 10459 1309 10468 1343
rect 11152 1343 11204 1352
rect 10416 1300 10468 1309
rect 11152 1309 11161 1343
rect 11161 1309 11195 1343
rect 11195 1309 11204 1343
rect 11152 1300 11204 1309
rect 11520 1368 11572 1420
rect 14464 1436 14516 1488
rect 12992 1368 13044 1420
rect 13728 1343 13780 1352
rect 13728 1309 13737 1343
rect 13737 1309 13771 1343
rect 13771 1309 13780 1343
rect 14924 1368 14976 1420
rect 15200 1411 15252 1420
rect 15200 1377 15209 1411
rect 15209 1377 15243 1411
rect 15243 1377 15252 1411
rect 15200 1368 15252 1377
rect 16120 1411 16172 1420
rect 16120 1377 16129 1411
rect 16129 1377 16163 1411
rect 16163 1377 16172 1411
rect 16120 1368 16172 1377
rect 13728 1300 13780 1309
rect 14740 1300 14792 1352
rect 15844 1343 15896 1352
rect 15844 1309 15853 1343
rect 15853 1309 15887 1343
rect 15887 1309 15896 1343
rect 15844 1300 15896 1309
rect 17776 1343 17828 1352
rect 17776 1309 17785 1343
rect 17785 1309 17819 1343
rect 17819 1309 17828 1343
rect 17776 1300 17828 1309
rect 17868 1343 17920 1352
rect 17868 1309 17877 1343
rect 17877 1309 17911 1343
rect 17911 1309 17920 1343
rect 18052 1343 18104 1352
rect 17868 1300 17920 1309
rect 18052 1309 18061 1343
rect 18061 1309 18095 1343
rect 18095 1309 18104 1343
rect 18052 1300 18104 1309
rect 18420 1300 18472 1352
rect 3608 1164 3660 1216
rect 4068 1207 4120 1216
rect 4068 1173 4077 1207
rect 4077 1173 4111 1207
rect 4111 1173 4120 1207
rect 4068 1164 4120 1173
rect 7104 1164 7156 1216
rect 8760 1164 8812 1216
rect 10324 1164 10376 1216
rect 11796 1164 11848 1216
rect 12256 1164 12308 1216
rect 13360 1232 13412 1284
rect 14924 1232 14976 1284
rect 15384 1232 15436 1284
rect 18236 1232 18288 1284
rect 13636 1207 13688 1216
rect 13636 1173 13645 1207
rect 13645 1173 13679 1207
rect 13679 1173 13688 1207
rect 13636 1164 13688 1173
rect 17960 1164 18012 1216
rect 18512 1207 18564 1216
rect 18512 1173 18521 1207
rect 18521 1173 18555 1207
rect 18555 1173 18564 1207
rect 18512 1164 18564 1173
rect 4660 1062 4712 1114
rect 4724 1062 4776 1114
rect 4788 1062 4840 1114
rect 4852 1062 4904 1114
rect 4916 1062 4968 1114
rect 7760 1062 7812 1114
rect 7824 1062 7876 1114
rect 7888 1062 7940 1114
rect 7952 1062 8004 1114
rect 8016 1062 8068 1114
rect 10860 1062 10912 1114
rect 10924 1062 10976 1114
rect 10988 1062 11040 1114
rect 11052 1062 11104 1114
rect 11116 1062 11168 1114
rect 13960 1062 14012 1114
rect 14024 1062 14076 1114
rect 14088 1062 14140 1114
rect 14152 1062 14204 1114
rect 14216 1062 14268 1114
rect 17060 1062 17112 1114
rect 17124 1062 17176 1114
rect 17188 1062 17240 1114
rect 17252 1062 17304 1114
rect 17316 1062 17368 1114
rect 2504 960 2556 1012
rect 5632 960 5684 1012
rect 7104 1003 7156 1012
rect 7104 969 7113 1003
rect 7113 969 7147 1003
rect 7147 969 7156 1003
rect 10324 1003 10376 1012
rect 7104 960 7156 969
rect 4068 892 4120 944
rect 5448 935 5500 944
rect 2596 824 2648 876
rect 5448 901 5457 935
rect 5457 901 5491 935
rect 5491 901 5500 935
rect 5448 892 5500 901
rect 10324 969 10333 1003
rect 10333 969 10367 1003
rect 10367 969 10376 1003
rect 10324 960 10376 969
rect 11336 960 11388 1012
rect 4988 867 5040 876
rect 4988 833 4997 867
rect 4997 833 5031 867
rect 5031 833 5040 867
rect 4988 824 5040 833
rect 5172 867 5224 876
rect 5172 833 5181 867
rect 5181 833 5215 867
rect 5215 833 5224 867
rect 10416 892 10468 944
rect 11796 935 11848 944
rect 11796 901 11805 935
rect 11805 901 11839 935
rect 11839 901 11848 935
rect 11796 892 11848 901
rect 13360 960 13412 1012
rect 13636 960 13688 1012
rect 15292 960 15344 1012
rect 18236 1003 18288 1012
rect 14464 935 14516 944
rect 14464 901 14473 935
rect 14473 901 14507 935
rect 14507 901 14516 935
rect 14464 892 14516 901
rect 14924 892 14976 944
rect 5172 824 5224 833
rect 2872 799 2924 808
rect 2872 765 2881 799
rect 2881 765 2915 799
rect 2915 765 2924 799
rect 2872 756 2924 765
rect 3884 756 3936 808
rect 5356 756 5408 808
rect 5908 756 5960 808
rect 7288 824 7340 876
rect 9036 824 9088 876
rect 5448 688 5500 740
rect 6368 799 6420 808
rect 6368 765 6377 799
rect 6377 765 6411 799
rect 6411 765 6420 799
rect 7748 799 7800 808
rect 6368 756 6420 765
rect 7748 765 7757 799
rect 7757 765 7791 799
rect 7791 765 7800 799
rect 7748 756 7800 765
rect 6552 688 6604 740
rect 4528 663 4580 672
rect 4528 629 4537 663
rect 4537 629 4571 663
rect 4571 629 4580 663
rect 4528 620 4580 629
rect 6828 663 6880 672
rect 6828 629 6837 663
rect 6837 629 6871 663
rect 6871 629 6880 663
rect 6828 620 6880 629
rect 9680 663 9732 672
rect 9680 629 9689 663
rect 9689 629 9723 663
rect 9723 629 9732 663
rect 9680 620 9732 629
rect 9864 824 9916 876
rect 10508 824 10560 876
rect 10968 824 11020 876
rect 11612 867 11664 876
rect 11612 833 11621 867
rect 11621 833 11655 867
rect 11655 833 11664 867
rect 11612 824 11664 833
rect 11888 867 11940 876
rect 10876 799 10928 808
rect 10876 765 10885 799
rect 10885 765 10919 799
rect 10919 765 10928 799
rect 10876 756 10928 765
rect 11888 833 11897 867
rect 11897 833 11931 867
rect 11931 833 11940 867
rect 11888 824 11940 833
rect 12072 867 12124 876
rect 12072 833 12081 867
rect 12081 833 12115 867
rect 12115 833 12124 867
rect 12072 824 12124 833
rect 18236 969 18245 1003
rect 18245 969 18279 1003
rect 18279 969 18288 1003
rect 18236 960 18288 969
rect 16948 892 17000 944
rect 18512 867 18564 876
rect 12808 756 12860 808
rect 13820 799 13872 808
rect 13820 765 13829 799
rect 13829 765 13863 799
rect 13863 765 13872 799
rect 18512 833 18521 867
rect 18521 833 18555 867
rect 18555 833 18564 867
rect 18512 824 18564 833
rect 16212 799 16264 808
rect 13820 756 13872 765
rect 16212 765 16221 799
rect 16221 765 16255 799
rect 16255 765 16264 799
rect 16212 756 16264 765
rect 17868 688 17920 740
rect 12164 620 12216 672
rect 3110 518 3162 570
rect 3174 518 3226 570
rect 3238 518 3290 570
rect 3302 518 3354 570
rect 3366 518 3418 570
rect 6210 518 6262 570
rect 6274 518 6326 570
rect 6338 518 6390 570
rect 6402 518 6454 570
rect 6466 518 6518 570
rect 9310 518 9362 570
rect 9374 518 9426 570
rect 9438 518 9490 570
rect 9502 518 9554 570
rect 9566 518 9618 570
rect 12410 518 12462 570
rect 12474 518 12526 570
rect 12538 518 12590 570
rect 12602 518 12654 570
rect 12666 518 12718 570
rect 15510 518 15562 570
rect 15574 518 15626 570
rect 15638 518 15690 570
rect 15702 518 15754 570
rect 15766 518 15818 570
rect 2872 416 2924 468
rect 3608 416 3660 468
rect 5908 416 5960 468
rect 7748 416 7800 468
rect 10508 459 10560 468
rect 10508 425 10517 459
rect 10517 425 10551 459
rect 10551 425 10560 459
rect 10508 416 10560 425
rect 12808 459 12860 468
rect 12808 425 12817 459
rect 12817 425 12851 459
rect 12851 425 12860 459
rect 12808 416 12860 425
rect 14648 416 14700 468
rect 16212 416 16264 468
rect 16580 416 16632 468
rect 18052 416 18104 468
rect 3608 212 3660 264
rect 18420 416 18472 468
rect 5356 323 5408 332
rect 5356 289 5365 323
rect 5365 289 5399 323
rect 5399 289 5408 323
rect 5356 280 5408 289
rect 6000 280 6052 332
rect 8760 323 8812 332
rect 8760 289 8769 323
rect 8769 289 8803 323
rect 8803 289 8812 323
rect 8760 280 8812 289
rect 9680 280 9732 332
rect 10140 323 10192 332
rect 10140 289 10149 323
rect 10149 289 10183 323
rect 10183 289 10192 323
rect 10140 280 10192 289
rect 12164 323 12216 332
rect 12164 289 12173 323
rect 12173 289 12207 323
rect 12207 289 12216 323
rect 12164 280 12216 289
rect 12256 280 12308 332
rect 12624 323 12676 332
rect 12624 289 12633 323
rect 12633 289 12667 323
rect 12667 289 12676 323
rect 12624 280 12676 289
rect 5172 212 5224 264
rect 6828 212 6880 264
rect 8668 255 8720 264
rect 8668 221 8677 255
rect 8677 221 8711 255
rect 8711 221 8720 255
rect 8668 212 8720 221
rect 10416 212 10468 264
rect 14648 255 14700 264
rect 14648 221 14657 255
rect 14657 221 14691 255
rect 14691 221 14700 255
rect 14648 212 14700 221
rect 16672 212 16724 264
rect 18144 212 18196 264
rect 3516 144 3568 196
rect 4528 144 4580 196
rect 6644 144 6696 196
rect 4660 -26 4712 26
rect 4724 -26 4776 26
rect 4788 -26 4840 26
rect 4852 -26 4904 26
rect 4916 -26 4968 26
rect 7760 -26 7812 26
rect 7824 -26 7876 26
rect 7888 -26 7940 26
rect 7952 -26 8004 26
rect 8016 -26 8068 26
rect 10860 -26 10912 26
rect 10924 -26 10976 26
rect 10988 -26 11040 26
rect 11052 -26 11104 26
rect 11116 -26 11168 26
rect 13960 -26 14012 26
rect 14024 -26 14076 26
rect 14088 -26 14140 26
rect 14152 -26 14204 26
rect 14216 -26 14268 26
rect 17060 -26 17112 26
rect 17124 -26 17176 26
rect 17188 -26 17240 26
rect 17252 -26 17304 26
rect 17316 -26 17368 26
<< metal2 >>
rect 1398 11200 1454 12000
rect 4250 11200 4306 12000
rect 7102 11200 7158 12000
rect 9954 11200 10010 12000
rect 12806 11200 12862 12000
rect 15396 11206 15608 11234
rect 572 10464 624 10470
rect 572 10406 624 10412
rect 584 9654 612 10406
rect 1412 10266 1440 11200
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2044 10736 2096 10742
rect 2044 10678 2096 10684
rect 1400 10260 1452 10266
rect 1400 10202 1452 10208
rect 1412 10062 1440 10202
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 2056 9722 2084 10678
rect 2424 10674 2452 10746
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 572 9648 624 9654
rect 572 9590 624 9596
rect 2056 9518 2084 9658
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 296 9512 348 9518
rect 296 9454 348 9460
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 308 8974 336 9454
rect 756 9376 808 9382
rect 756 9318 808 9324
rect 768 8974 796 9318
rect 2056 8974 2084 9454
rect 296 8968 348 8974
rect 296 8910 348 8916
rect 756 8968 808 8974
rect 756 8910 808 8916
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 296 8832 348 8838
rect 296 8774 348 8780
rect 664 8832 716 8838
rect 664 8774 716 8780
rect 308 8498 336 8774
rect 676 8498 704 8774
rect 296 8492 348 8498
rect 296 8434 348 8440
rect 664 8492 716 8498
rect 664 8434 716 8440
rect 572 7744 624 7750
rect 572 7686 624 7692
rect 584 7478 612 7686
rect 572 7472 624 7478
rect 572 7414 624 7420
rect 768 7206 796 8910
rect 2148 8634 2176 9522
rect 2424 9489 2452 10610
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2516 9586 2544 10406
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2410 9480 2466 9489
rect 2410 9415 2466 9424
rect 2424 9178 2452 9415
rect 2608 9382 2636 9658
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2608 8294 2636 9318
rect 2792 9042 2820 9658
rect 2884 9058 2912 10610
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 2976 10062 3004 10542
rect 3110 10364 3418 10384
rect 3110 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3276 10364
rect 3332 10362 3356 10364
rect 3412 10362 3418 10364
rect 3172 10310 3174 10362
rect 3354 10310 3356 10362
rect 3110 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3276 10310
rect 3332 10308 3356 10310
rect 3412 10308 3418 10310
rect 3110 10288 3418 10308
rect 3700 10192 3752 10198
rect 3146 10160 3202 10169
rect 3700 10134 3752 10140
rect 3974 10160 4030 10169
rect 3146 10095 3202 10104
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2976 9160 3004 9522
rect 3160 9466 3188 10095
rect 3332 10056 3384 10062
rect 3238 10024 3294 10033
rect 3384 10016 3648 10044
rect 3332 9998 3384 10004
rect 3238 9959 3294 9968
rect 3252 9926 3280 9959
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3436 9722 3464 9862
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3332 9512 3384 9518
rect 3068 9450 3188 9466
rect 3056 9444 3188 9450
rect 3108 9438 3188 9444
rect 3330 9480 3332 9489
rect 3384 9480 3386 9489
rect 3330 9415 3386 9424
rect 3056 9386 3108 9392
rect 3528 9382 3556 9590
rect 3620 9382 3648 10016
rect 3712 9926 3740 10134
rect 3974 10095 3976 10104
rect 4028 10095 4030 10104
rect 3976 10066 4028 10072
rect 3974 10024 4030 10033
rect 3974 9959 3976 9968
rect 4028 9959 4030 9968
rect 3976 9930 4028 9936
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 3700 9716 3752 9722
rect 4068 9716 4120 9722
rect 3752 9676 4068 9704
rect 3700 9658 3752 9664
rect 4068 9658 4120 9664
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3110 9276 3418 9296
rect 3110 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3276 9276
rect 3332 9274 3356 9276
rect 3412 9274 3418 9276
rect 3172 9222 3174 9274
rect 3354 9222 3356 9274
rect 3110 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3276 9222
rect 3332 9220 3356 9222
rect 3412 9220 3418 9222
rect 3110 9200 3418 9220
rect 2976 9132 3096 9160
rect 2884 9042 3004 9058
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2884 9036 3016 9042
rect 2884 9030 2964 9036
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2700 8838 2728 8910
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2700 8634 2728 8774
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2884 8498 2912 9030
rect 2964 8978 3016 8984
rect 3068 8974 3096 9132
rect 3620 8974 3648 9318
rect 3712 9178 3740 9522
rect 3976 9512 4028 9518
rect 3804 9472 3976 9500
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3804 8906 3832 9472
rect 3976 9454 4028 9460
rect 4172 9042 4200 9862
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 2240 7546 2268 7686
rect 2424 7546 2452 7822
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2608 7478 2636 8230
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 2596 7472 2648 7478
rect 2596 7414 2648 7420
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 756 7200 808 7206
rect 756 7142 808 7148
rect 768 6458 796 7142
rect 2332 6730 2360 7346
rect 2608 7206 2636 7414
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2320 6724 2372 6730
rect 2320 6666 2372 6672
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 756 6452 808 6458
rect 756 6394 808 6400
rect 768 5710 796 6394
rect 1860 6384 1912 6390
rect 1860 6326 1912 6332
rect 940 6112 992 6118
rect 940 6054 992 6060
rect 756 5704 808 5710
rect 756 5646 808 5652
rect 480 5568 532 5574
rect 480 5510 532 5516
rect 492 5234 520 5510
rect 952 5234 980 6054
rect 1872 5302 1900 6326
rect 1964 6254 1992 6598
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 2056 6118 2084 6598
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 2056 5846 2084 6054
rect 2044 5840 2096 5846
rect 2044 5782 2096 5788
rect 2332 5794 2360 6666
rect 2424 6322 2452 6666
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2424 5914 2452 6258
rect 2608 6100 2636 7142
rect 2792 7002 2820 7958
rect 2976 7954 3004 8230
rect 3110 8188 3418 8208
rect 3110 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3276 8188
rect 3332 8186 3356 8188
rect 3412 8186 3418 8188
rect 3172 8134 3174 8186
rect 3354 8134 3356 8186
rect 3110 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3276 8134
rect 3332 8132 3356 8134
rect 3412 8132 3418 8134
rect 3110 8112 3418 8132
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 3068 7546 3096 7686
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3804 7342 3832 8842
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3896 8498 3924 8774
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 3988 7750 4016 8366
rect 4264 8090 4292 11200
rect 4660 10908 4968 10928
rect 4660 10906 4666 10908
rect 4722 10906 4746 10908
rect 4802 10906 4826 10908
rect 4882 10906 4906 10908
rect 4962 10906 4968 10908
rect 4722 10854 4724 10906
rect 4904 10854 4906 10906
rect 4660 10852 4666 10854
rect 4722 10852 4746 10854
rect 4802 10852 4826 10854
rect 4882 10852 4906 10854
rect 4962 10852 4968 10854
rect 4660 10832 4968 10852
rect 7116 10810 7144 11200
rect 7760 10908 8068 10928
rect 7760 10906 7766 10908
rect 7822 10906 7846 10908
rect 7902 10906 7926 10908
rect 7982 10906 8006 10908
rect 8062 10906 8068 10908
rect 7822 10854 7824 10906
rect 8004 10854 8006 10906
rect 7760 10852 7766 10854
rect 7822 10852 7846 10854
rect 7902 10852 7926 10854
rect 7982 10852 8006 10854
rect 8062 10852 8068 10854
rect 7760 10832 8068 10852
rect 9968 10810 9996 11200
rect 10860 10908 11168 10928
rect 10860 10906 10866 10908
rect 10922 10906 10946 10908
rect 11002 10906 11026 10908
rect 11082 10906 11106 10908
rect 11162 10906 11168 10908
rect 10922 10854 10924 10906
rect 11104 10854 11106 10906
rect 10860 10852 10866 10854
rect 10922 10852 10946 10854
rect 11002 10852 11026 10854
rect 11082 10852 11106 10854
rect 11162 10852 11168 10854
rect 10860 10832 11168 10852
rect 12820 10810 12848 11200
rect 13960 10908 14268 10928
rect 13960 10906 13966 10908
rect 14022 10906 14046 10908
rect 14102 10906 14126 10908
rect 14182 10906 14206 10908
rect 14262 10906 14268 10908
rect 14022 10854 14024 10906
rect 14204 10854 14206 10906
rect 13960 10852 13966 10854
rect 14022 10852 14046 10854
rect 14102 10852 14126 10854
rect 14182 10852 14206 10854
rect 14262 10852 14268 10854
rect 13960 10832 14268 10852
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 6210 10364 6518 10384
rect 6210 10362 6216 10364
rect 6272 10362 6296 10364
rect 6352 10362 6376 10364
rect 6432 10362 6456 10364
rect 6512 10362 6518 10364
rect 6272 10310 6274 10362
rect 6454 10310 6456 10362
rect 6210 10308 6216 10310
rect 6272 10308 6296 10310
rect 6352 10308 6376 10310
rect 6432 10308 6456 10310
rect 6512 10308 6518 10310
rect 6210 10288 6518 10308
rect 7484 10266 7512 10610
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 9310 10364 9618 10384
rect 9310 10362 9316 10364
rect 9372 10362 9396 10364
rect 9452 10362 9476 10364
rect 9532 10362 9556 10364
rect 9612 10362 9618 10364
rect 9372 10310 9374 10362
rect 9554 10310 9556 10362
rect 9310 10308 9316 10310
rect 9372 10308 9396 10310
rect 9452 10308 9476 10310
rect 9532 10308 9556 10310
rect 9612 10308 9618 10310
rect 9310 10288 9618 10308
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 4448 9994 4476 10202
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 4660 9820 4968 9840
rect 4660 9818 4666 9820
rect 4722 9818 4746 9820
rect 4802 9818 4826 9820
rect 4882 9818 4906 9820
rect 4962 9818 4968 9820
rect 4722 9766 4724 9818
rect 4904 9766 4906 9818
rect 4660 9764 4666 9766
rect 4722 9764 4746 9766
rect 4802 9764 4826 9766
rect 4882 9764 4906 9766
rect 4962 9764 4968 9766
rect 4660 9744 4968 9764
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4540 8838 4568 9454
rect 4816 9178 4844 9522
rect 5184 9364 5212 9590
rect 5276 9586 5304 9862
rect 5920 9654 5948 10202
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5264 9376 5316 9382
rect 5184 9336 5264 9364
rect 5264 9318 5316 9324
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4816 9042 4844 9114
rect 4804 9036 4856 9042
rect 4804 8978 4856 8984
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4660 8732 4968 8752
rect 4660 8730 4666 8732
rect 4722 8730 4746 8732
rect 4802 8730 4826 8732
rect 4882 8730 4906 8732
rect 4962 8730 4968 8732
rect 4722 8678 4724 8730
rect 4904 8678 4906 8730
rect 4660 8676 4666 8678
rect 4722 8676 4746 8678
rect 4802 8676 4826 8678
rect 4882 8676 4906 8678
rect 4962 8676 4968 8678
rect 4660 8656 4968 8676
rect 5000 8634 5028 8842
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3988 7546 4016 7686
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3110 7100 3418 7120
rect 3110 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3276 7100
rect 3332 7098 3356 7100
rect 3412 7098 3418 7100
rect 3172 7046 3174 7098
rect 3354 7046 3356 7098
rect 3110 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3276 7046
rect 3332 7044 3356 7046
rect 3412 7044 3418 7046
rect 3110 7024 3418 7044
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 2976 6798 3004 6938
rect 3804 6798 3832 7278
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 2976 6458 3004 6734
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 6458 3924 6598
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 2976 6254 3004 6394
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 4080 6186 4108 7890
rect 4724 7886 4752 8298
rect 5092 7886 5120 8774
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 4172 6866 4200 7822
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4660 7644 4968 7664
rect 4660 7642 4666 7644
rect 4722 7642 4746 7644
rect 4802 7642 4826 7644
rect 4882 7642 4906 7644
rect 4962 7642 4968 7644
rect 4722 7590 4724 7642
rect 4904 7590 4906 7642
rect 4660 7588 4666 7590
rect 4722 7588 4746 7590
rect 4802 7588 4826 7590
rect 4882 7588 4906 7590
rect 4962 7588 4968 7590
rect 4660 7568 4968 7588
rect 5092 7342 5120 7686
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4356 6322 4384 6598
rect 4660 6556 4968 6576
rect 4660 6554 4666 6556
rect 4722 6554 4746 6556
rect 4802 6554 4826 6556
rect 4882 6554 4906 6556
rect 4962 6554 4968 6556
rect 4722 6502 4724 6554
rect 4904 6502 4906 6554
rect 4660 6500 4666 6502
rect 4722 6500 4746 6502
rect 4802 6500 4826 6502
rect 4882 6500 4906 6502
rect 4962 6500 4968 6502
rect 4660 6480 4968 6500
rect 5184 6458 5212 8434
rect 5276 7188 5304 9318
rect 5644 9178 5672 9454
rect 6104 9382 6132 10066
rect 6840 9994 6868 10202
rect 11072 10062 11100 10406
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5368 8498 5396 8910
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 5368 7818 5396 7958
rect 5736 7886 5764 8502
rect 5828 8430 5856 9046
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5644 7410 5672 7686
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5356 7200 5408 7206
rect 5276 7160 5356 7188
rect 5356 7142 5408 7148
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 2688 6112 2740 6118
rect 2608 6072 2688 6100
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2332 5766 2452 5794
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2332 5370 2360 5646
rect 2424 5574 2452 5766
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2608 5302 2636 6072
rect 2688 6054 2740 6060
rect 3110 6012 3418 6032
rect 3110 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3276 6012
rect 3332 6010 3356 6012
rect 3412 6010 3418 6012
rect 3172 5958 3174 6010
rect 3354 5958 3356 6010
rect 3110 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3276 5958
rect 3332 5956 3356 5958
rect 3412 5956 3418 5958
rect 3110 5936 3418 5956
rect 4080 5846 4108 6122
rect 4264 5914 4292 6258
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4068 5840 4120 5846
rect 3988 5788 4068 5794
rect 3988 5782 4120 5788
rect 3988 5766 4108 5782
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2872 5568 2924 5574
rect 3068 5556 3096 5646
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 2924 5528 3096 5556
rect 2872 5510 2924 5516
rect 1860 5296 1912 5302
rect 1860 5238 1912 5244
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 480 5228 532 5234
rect 480 5170 532 5176
rect 940 5228 992 5234
rect 940 5170 992 5176
rect 2608 5030 2636 5238
rect 3068 5166 3096 5528
rect 3896 5166 3924 5578
rect 3988 5574 4016 5766
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 4080 5234 4108 5646
rect 5184 5642 5212 6394
rect 5460 6254 5488 6802
rect 5828 6390 5856 8366
rect 6104 7886 6132 9318
rect 6210 9276 6518 9296
rect 6210 9274 6216 9276
rect 6272 9274 6296 9276
rect 6352 9274 6376 9276
rect 6432 9274 6456 9276
rect 6512 9274 6518 9276
rect 6272 9222 6274 9274
rect 6454 9222 6456 9274
rect 6210 9220 6216 9222
rect 6272 9220 6296 9222
rect 6352 9220 6376 9222
rect 6432 9220 6456 9222
rect 6512 9220 6518 9222
rect 6210 9200 6518 9220
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6472 8498 6500 8978
rect 6564 8634 6592 9862
rect 7668 9722 7696 9862
rect 7760 9820 8068 9840
rect 7760 9818 7766 9820
rect 7822 9818 7846 9820
rect 7902 9818 7926 9820
rect 7982 9818 8006 9820
rect 8062 9818 8068 9820
rect 7822 9766 7824 9818
rect 8004 9766 8006 9818
rect 7760 9764 7766 9766
rect 7822 9764 7846 9766
rect 7902 9764 7926 9766
rect 7982 9764 8006 9766
rect 8062 9764 8068 9766
rect 7760 9744 8068 9764
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7208 8974 7236 9386
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 9042 7328 9318
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 7024 8498 7052 8910
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8566 7420 8774
rect 7668 8566 7696 9658
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 7760 9178 7788 9454
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7760 8732 8068 8752
rect 7760 8730 7766 8732
rect 7822 8730 7846 8732
rect 7902 8730 7926 8732
rect 7982 8730 8006 8732
rect 8062 8730 8068 8732
rect 7822 8678 7824 8730
rect 8004 8678 8006 8730
rect 7760 8676 7766 8678
rect 7822 8676 7846 8678
rect 7902 8676 7926 8678
rect 7982 8676 8006 8678
rect 8062 8676 8068 8678
rect 7760 8656 8068 8676
rect 7380 8560 7432 8566
rect 7380 8502 7432 8508
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 6210 8188 6518 8208
rect 6210 8186 6216 8188
rect 6272 8186 6296 8188
rect 6352 8186 6376 8188
rect 6432 8186 6456 8188
rect 6512 8186 6518 8188
rect 6272 8134 6274 8186
rect 6454 8134 6456 8186
rect 6210 8132 6216 8134
rect 6272 8132 6296 8134
rect 6352 8132 6376 8134
rect 6432 8132 6456 8134
rect 6512 8132 6518 8134
rect 6210 8112 6518 8132
rect 7208 8022 7236 8366
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6196 7546 6224 7686
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 5908 7472 5960 7478
rect 5908 7414 5960 7420
rect 5920 7206 5948 7414
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 6210 7100 6518 7120
rect 6210 7098 6216 7100
rect 6272 7098 6296 7100
rect 6352 7098 6376 7100
rect 6432 7098 6456 7100
rect 6512 7098 6518 7100
rect 6272 7046 6274 7098
rect 6454 7046 6456 7098
rect 6210 7044 6216 7046
rect 6272 7044 6296 7046
rect 6352 7044 6376 7046
rect 6432 7044 6456 7046
rect 6512 7044 6518 7046
rect 6210 7024 6518 7044
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6748 6390 6776 6666
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5644 5914 5672 6258
rect 6210 6012 6518 6032
rect 6210 6010 6216 6012
rect 6272 6010 6296 6012
rect 6352 6010 6376 6012
rect 6432 6010 6456 6012
rect 6512 6010 6518 6012
rect 6272 5958 6274 6010
rect 6454 5958 6456 6010
rect 6210 5956 6216 5958
rect 6272 5956 6296 5958
rect 6352 5956 6376 5958
rect 6432 5956 6456 5958
rect 6512 5956 6518 5958
rect 6210 5936 6518 5956
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 6840 5710 6868 7754
rect 6932 6254 6960 7890
rect 7668 7886 7696 8230
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7656 7744 7708 7750
rect 7760 7732 7788 8366
rect 8128 7954 8156 9454
rect 8588 9450 8616 9658
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8864 9178 8892 9998
rect 11164 9994 11192 10542
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10336 9654 10364 9862
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8956 9110 8984 9454
rect 9310 9276 9618 9296
rect 9310 9274 9316 9276
rect 9372 9274 9396 9276
rect 9452 9274 9476 9276
rect 9532 9274 9556 9276
rect 9612 9274 9618 9276
rect 9372 9222 9374 9274
rect 9554 9222 9556 9274
rect 9310 9220 9316 9222
rect 9372 9220 9396 9222
rect 9452 9220 9476 9222
rect 9532 9220 9556 9222
rect 9612 9220 9618 9222
rect 9310 9200 9618 9220
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 8772 8956 8800 9046
rect 8852 8968 8904 8974
rect 8772 8928 8852 8956
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 7708 7704 7788 7732
rect 7656 7686 7708 7692
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7576 5710 7604 6054
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 5172 5636 5224 5642
rect 5172 5578 5224 5584
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 4660 5468 4968 5488
rect 4660 5466 4666 5468
rect 4722 5466 4746 5468
rect 4802 5466 4826 5468
rect 4882 5466 4906 5468
rect 4962 5466 4968 5468
rect 4722 5414 4724 5466
rect 4904 5414 4906 5466
rect 4660 5412 4666 5414
rect 4722 5412 4746 5414
rect 4802 5412 4826 5414
rect 4882 5412 4906 5414
rect 4962 5412 4968 5414
rect 4660 5392 4968 5412
rect 5276 5370 5304 5510
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 7484 5234 7512 5646
rect 7668 5302 7696 7686
rect 7760 7644 8068 7664
rect 7760 7642 7766 7644
rect 7822 7642 7846 7644
rect 7902 7642 7926 7644
rect 7982 7642 8006 7644
rect 8062 7642 8068 7644
rect 7822 7590 7824 7642
rect 8004 7590 8006 7642
rect 7760 7588 7766 7590
rect 7822 7588 7846 7590
rect 7902 7588 7926 7590
rect 7982 7588 8006 7590
rect 8062 7588 8068 7590
rect 7760 7568 8068 7588
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 7760 6556 8068 6576
rect 7760 6554 7766 6556
rect 7822 6554 7846 6556
rect 7902 6554 7926 6556
rect 7982 6554 8006 6556
rect 8062 6554 8068 6556
rect 7822 6502 7824 6554
rect 8004 6502 8006 6554
rect 7760 6500 7766 6502
rect 7822 6500 7846 6502
rect 7902 6500 7926 6502
rect 7982 6500 8006 6502
rect 8062 6500 8068 6502
rect 7760 6480 8068 6500
rect 8128 6322 8156 6598
rect 8220 6390 8248 6734
rect 8404 6662 8432 7890
rect 8772 7410 8800 8928
rect 8852 8910 8904 8916
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8864 8498 8892 8774
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8956 8362 8984 9046
rect 9692 9042 9720 9522
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9324 8634 9352 8910
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9588 8560 9640 8566
rect 9784 8514 9812 8910
rect 9640 8508 9812 8514
rect 9588 8502 9812 8508
rect 9600 8486 9812 8502
rect 9968 8498 9996 8978
rect 10336 8974 10364 9590
rect 10704 9586 10732 9862
rect 10860 9820 11168 9840
rect 10860 9818 10866 9820
rect 10922 9818 10946 9820
rect 11002 9818 11026 9820
rect 11082 9818 11106 9820
rect 11162 9818 11168 9820
rect 10922 9766 10924 9818
rect 11104 9766 11106 9818
rect 10860 9764 10866 9766
rect 10922 9764 10946 9766
rect 11002 9764 11026 9766
rect 11082 9764 11106 9766
rect 11162 9764 11168 9766
rect 10860 9744 11168 9764
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10324 8968 10376 8974
rect 10244 8928 10324 8956
rect 10244 8498 10272 8928
rect 10324 8910 10376 8916
rect 10428 8566 10456 8978
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 9784 8242 9812 8486
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 9956 8288 10008 8294
rect 9784 8236 9956 8242
rect 9784 8230 10008 8236
rect 9784 8214 9996 8230
rect 9310 8188 9618 8208
rect 9310 8186 9316 8188
rect 9372 8186 9396 8188
rect 9452 8186 9476 8188
rect 9532 8186 9556 8188
rect 9612 8186 9618 8188
rect 9372 8134 9374 8186
rect 9554 8134 9556 8186
rect 9310 8132 9316 8134
rect 9372 8132 9396 8134
rect 9452 8132 9476 8134
rect 9532 8132 9556 8134
rect 9612 8132 9618 8134
rect 9310 8112 9618 8132
rect 9876 7886 9904 8214
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8404 6254 8432 6598
rect 8588 6458 8616 7142
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8496 5914 8524 6258
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 7760 5468 8068 5488
rect 7760 5466 7766 5468
rect 7822 5466 7846 5468
rect 7902 5466 7926 5468
rect 7982 5466 8006 5468
rect 8062 5466 8068 5468
rect 7822 5414 7824 5466
rect 8004 5414 8006 5466
rect 7760 5412 7766 5414
rect 7822 5412 7846 5414
rect 7902 5412 7926 5414
rect 7982 5412 8006 5414
rect 8062 5412 8068 5414
rect 7760 5392 8068 5412
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2608 4486 2636 4966
rect 3110 4924 3418 4944
rect 3110 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3276 4924
rect 3332 4922 3356 4924
rect 3412 4922 3418 4924
rect 3172 4870 3174 4922
rect 3354 4870 3356 4922
rect 3110 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3276 4870
rect 3332 4868 3356 4870
rect 3412 4868 3418 4870
rect 3110 4848 3418 4868
rect 6210 4924 6518 4944
rect 6210 4922 6216 4924
rect 6272 4922 6296 4924
rect 6352 4922 6376 4924
rect 6432 4922 6456 4924
rect 6512 4922 6518 4924
rect 6272 4870 6274 4922
rect 6454 4870 6456 4922
rect 6210 4868 6216 4870
rect 6272 4868 6296 4870
rect 6352 4868 6376 4870
rect 6432 4868 6456 4870
rect 6512 4868 6518 4870
rect 6210 4848 6518 4868
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 480 4480 532 4486
rect 480 4422 532 4428
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 492 4146 520 4422
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 480 4140 532 4146
rect 480 4082 532 4088
rect 2424 4078 2452 4218
rect 2608 4214 2636 4422
rect 2596 4208 2648 4214
rect 2596 4150 2648 4156
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2792 3738 2820 3878
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2688 3664 2740 3670
rect 2688 3606 2740 3612
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 2320 3460 2372 3466
rect 2320 3402 2372 3408
rect 572 3392 624 3398
rect 572 3334 624 3340
rect 584 3126 612 3334
rect 2332 3126 2360 3402
rect 2608 3194 2636 3470
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 572 3120 624 3126
rect 572 3062 624 3068
rect 2320 3120 2372 3126
rect 2320 3062 2372 3068
rect 2700 3058 2728 3606
rect 2884 3398 2912 4150
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 296 2984 348 2990
rect 296 2926 348 2932
rect 308 1902 336 2926
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 848 2304 900 2310
rect 848 2246 900 2252
rect 860 2038 888 2246
rect 1216 2100 1268 2106
rect 1216 2042 1268 2048
rect 848 2032 900 2038
rect 848 1974 900 1980
rect 1228 1902 1256 2042
rect 296 1896 348 1902
rect 296 1838 348 1844
rect 1216 1896 1268 1902
rect 1216 1838 1268 1844
rect 1228 1426 1256 1838
rect 2516 1766 2544 2790
rect 2976 2106 3004 4626
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 3516 4548 3568 4554
rect 3516 4490 3568 4496
rect 3528 4282 3556 4490
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 4660 4380 4968 4400
rect 4660 4378 4666 4380
rect 4722 4378 4746 4380
rect 4802 4378 4826 4380
rect 4882 4378 4906 4380
rect 4962 4378 4968 4380
rect 4722 4326 4724 4378
rect 4904 4326 4906 4378
rect 4660 4324 4666 4326
rect 4722 4324 4746 4326
rect 4802 4324 4826 4326
rect 4882 4324 4906 4326
rect 4962 4324 4968 4326
rect 4660 4304 4968 4324
rect 3516 4276 3568 4282
rect 3516 4218 3568 4224
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 3054 4176 3110 4185
rect 3054 4111 3056 4120
rect 3108 4111 3110 4120
rect 3514 4176 3570 4185
rect 4356 4146 4384 4218
rect 4986 4176 5042 4185
rect 3514 4111 3570 4120
rect 3792 4140 3844 4146
rect 3056 4082 3108 4088
rect 3528 3942 3556 4111
rect 3792 4082 3844 4088
rect 4344 4140 4396 4146
rect 5460 4146 5488 4422
rect 6472 4282 6500 4558
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 4986 4111 4988 4120
rect 4344 4082 4396 4088
rect 5040 4111 5042 4120
rect 5448 4140 5500 4146
rect 4988 4082 5040 4088
rect 5448 4082 5500 4088
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3110 3836 3418 3856
rect 3110 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3276 3836
rect 3332 3834 3356 3836
rect 3412 3834 3418 3836
rect 3172 3782 3174 3834
rect 3354 3782 3356 3834
rect 3110 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3276 3782
rect 3332 3780 3356 3782
rect 3412 3780 3418 3782
rect 3110 3760 3418 3780
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 3160 3194 3188 3470
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3528 2990 3556 3878
rect 3804 3602 3832 4082
rect 6932 4010 6960 4626
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7668 4146 7696 4558
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 7760 4380 8068 4400
rect 7760 4378 7766 4380
rect 7822 4378 7846 4380
rect 7902 4378 7926 4380
rect 7982 4378 8006 4380
rect 8062 4378 8068 4380
rect 7822 4326 7824 4378
rect 8004 4326 8006 4378
rect 7760 4324 7766 4326
rect 7822 4324 7846 4326
rect 7902 4324 7926 4326
rect 7982 4324 8006 4326
rect 8062 4324 8068 4326
rect 7760 4304 8068 4324
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 3792 3596 3844 3602
rect 3792 3538 3844 3544
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4080 3194 4108 3470
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4172 3058 4200 3334
rect 4264 3058 4292 3538
rect 4632 3534 4660 3878
rect 5000 3602 5028 3878
rect 6210 3836 6518 3856
rect 6210 3834 6216 3836
rect 6272 3834 6296 3836
rect 6352 3834 6376 3836
rect 6432 3834 6456 3836
rect 6512 3834 6518 3836
rect 6272 3782 6274 3834
rect 6454 3782 6456 3834
rect 6210 3780 6216 3782
rect 6272 3780 6296 3782
rect 6352 3780 6376 3782
rect 6432 3780 6456 3782
rect 6512 3780 6518 3782
rect 6210 3760 6518 3780
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 4660 3292 4968 3312
rect 4660 3290 4666 3292
rect 4722 3290 4746 3292
rect 4802 3290 4826 3292
rect 4882 3290 4906 3292
rect 4962 3290 4968 3292
rect 4722 3238 4724 3290
rect 4904 3238 4906 3290
rect 4660 3236 4666 3238
rect 4722 3236 4746 3238
rect 4802 3236 4826 3238
rect 4882 3236 4906 3238
rect 4962 3236 4968 3238
rect 4660 3216 4968 3236
rect 5460 3194 5488 3402
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3110 2748 3418 2768
rect 3110 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3276 2748
rect 3332 2746 3356 2748
rect 3412 2746 3418 2748
rect 3172 2694 3174 2746
rect 3354 2694 3356 2746
rect 3110 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3276 2694
rect 3332 2692 3356 2694
rect 3412 2692 3418 2694
rect 3110 2672 3418 2692
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 2964 2100 3016 2106
rect 2964 2042 3016 2048
rect 3528 2038 3556 2586
rect 3712 2514 3740 2994
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 3804 2582 3832 2790
rect 3792 2576 3844 2582
rect 3792 2518 3844 2524
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 3804 2106 3832 2246
rect 4356 2106 4384 2790
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 4660 2204 4968 2224
rect 4660 2202 4666 2204
rect 4722 2202 4746 2204
rect 4802 2202 4826 2204
rect 4882 2202 4906 2204
rect 4962 2202 4968 2204
rect 4722 2150 4724 2202
rect 4904 2150 4906 2202
rect 4660 2148 4666 2150
rect 4722 2148 4746 2150
rect 4802 2148 4826 2150
rect 4882 2148 4906 2150
rect 4962 2148 4968 2150
rect 4660 2128 4968 2148
rect 5276 2106 5304 2246
rect 3792 2100 3844 2106
rect 3792 2042 3844 2048
rect 4344 2100 4396 2106
rect 4344 2042 4396 2048
rect 5264 2100 5316 2106
rect 5264 2042 5316 2048
rect 2780 2032 2832 2038
rect 2780 1974 2832 1980
rect 3516 2032 3568 2038
rect 3516 1974 3568 1980
rect 2596 1828 2648 1834
rect 2596 1770 2648 1776
rect 2504 1760 2556 1766
rect 2504 1702 2556 1708
rect 1216 1420 1268 1426
rect 1216 1362 1268 1368
rect 2516 1222 2544 1702
rect 2504 1216 2556 1222
rect 2504 1158 2556 1164
rect 2516 1018 2544 1158
rect 2504 1012 2556 1018
rect 2504 954 2556 960
rect 2608 882 2636 1770
rect 2792 1494 2820 1974
rect 2964 1964 3016 1970
rect 2964 1906 3016 1912
rect 2872 1760 2924 1766
rect 2872 1702 2924 1708
rect 2780 1488 2832 1494
rect 2780 1430 2832 1436
rect 2792 1306 2820 1430
rect 2884 1426 2912 1702
rect 2976 1562 3004 1906
rect 3528 1766 3556 1974
rect 3884 1964 3936 1970
rect 3884 1906 3936 1912
rect 3516 1760 3568 1766
rect 3516 1702 3568 1708
rect 3110 1660 3418 1680
rect 3110 1658 3116 1660
rect 3172 1658 3196 1660
rect 3252 1658 3276 1660
rect 3332 1658 3356 1660
rect 3412 1658 3418 1660
rect 3172 1606 3174 1658
rect 3354 1606 3356 1658
rect 3110 1604 3116 1606
rect 3172 1604 3196 1606
rect 3252 1604 3276 1606
rect 3332 1604 3356 1606
rect 3412 1604 3418 1606
rect 3110 1584 3418 1604
rect 2964 1556 3016 1562
rect 2964 1498 3016 1504
rect 2872 1420 2924 1426
rect 2872 1362 2924 1368
rect 2792 1290 2912 1306
rect 2792 1284 2924 1290
rect 2792 1278 2872 1284
rect 2872 1226 2924 1232
rect 3332 1284 3384 1290
rect 3332 1226 3384 1232
rect 2596 876 2648 882
rect 2596 818 2648 824
rect 2872 808 2924 814
rect 2872 750 2924 756
rect 2884 474 2912 750
rect 3344 728 3372 1226
rect 3528 864 3556 1702
rect 3700 1556 3752 1562
rect 3700 1498 3752 1504
rect 3712 1358 3740 1498
rect 3896 1494 3924 1906
rect 3884 1488 3936 1494
rect 3884 1430 3936 1436
rect 3700 1352 3752 1358
rect 3606 1320 3662 1329
rect 3700 1294 3752 1300
rect 3606 1255 3662 1264
rect 3620 1222 3648 1255
rect 3608 1216 3660 1222
rect 3608 1158 3660 1164
rect 3528 836 3648 864
rect 3344 700 3556 728
rect 3110 572 3418 592
rect 3110 570 3116 572
rect 3172 570 3196 572
rect 3252 570 3276 572
rect 3332 570 3356 572
rect 3412 570 3418 572
rect 3172 518 3174 570
rect 3354 518 3356 570
rect 3110 516 3116 518
rect 3172 516 3196 518
rect 3252 516 3276 518
rect 3332 516 3356 518
rect 3412 516 3418 518
rect 3110 496 3418 516
rect 2872 468 2924 474
rect 2872 410 2924 416
rect 3528 202 3556 700
rect 3620 474 3648 836
rect 3896 814 3924 1430
rect 4988 1352 5040 1358
rect 4988 1294 5040 1300
rect 4068 1216 4120 1222
rect 4068 1158 4120 1164
rect 4080 950 4108 1158
rect 4660 1116 4968 1136
rect 4660 1114 4666 1116
rect 4722 1114 4746 1116
rect 4802 1114 4826 1116
rect 4882 1114 4906 1116
rect 4962 1114 4968 1116
rect 4722 1062 4724 1114
rect 4904 1062 4906 1114
rect 4660 1060 4666 1062
rect 4722 1060 4746 1062
rect 4802 1060 4826 1062
rect 4882 1060 4906 1062
rect 4962 1060 4968 1062
rect 4660 1040 4968 1060
rect 4068 944 4120 950
rect 4068 886 4120 892
rect 5000 882 5028 1294
rect 5460 950 5488 2450
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5552 1329 5580 2382
rect 5644 2378 5672 3606
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6656 3398 6684 3470
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 5736 3194 5764 3334
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5632 2372 5684 2378
rect 5632 2314 5684 2320
rect 5644 2106 5672 2314
rect 5632 2100 5684 2106
rect 5632 2042 5684 2048
rect 5736 1902 5764 3130
rect 6012 2990 6040 3334
rect 6564 3126 6592 3334
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 6210 2748 6518 2768
rect 6210 2746 6216 2748
rect 6272 2746 6296 2748
rect 6352 2746 6376 2748
rect 6432 2746 6456 2748
rect 6512 2746 6518 2748
rect 6272 2694 6274 2746
rect 6454 2694 6456 2746
rect 6210 2692 6216 2694
rect 6272 2692 6296 2694
rect 6352 2692 6376 2694
rect 6432 2692 6456 2694
rect 6512 2692 6518 2694
rect 6210 2672 6518 2692
rect 6564 2446 6592 3062
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 6656 2106 6684 3334
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 5908 1964 5960 1970
rect 5908 1906 5960 1912
rect 5724 1896 5776 1902
rect 5724 1838 5776 1844
rect 5920 1562 5948 1906
rect 6000 1896 6052 1902
rect 6000 1838 6052 1844
rect 6552 1896 6604 1902
rect 6552 1838 6604 1844
rect 5908 1556 5960 1562
rect 5908 1498 5960 1504
rect 6012 1426 6040 1838
rect 6092 1828 6144 1834
rect 6092 1770 6144 1776
rect 6104 1562 6132 1770
rect 6210 1660 6518 1680
rect 6210 1658 6216 1660
rect 6272 1658 6296 1660
rect 6352 1658 6376 1660
rect 6432 1658 6456 1660
rect 6512 1658 6518 1660
rect 6272 1606 6274 1658
rect 6454 1606 6456 1658
rect 6210 1604 6216 1606
rect 6272 1604 6296 1606
rect 6352 1604 6376 1606
rect 6432 1604 6456 1606
rect 6512 1604 6518 1606
rect 6210 1584 6518 1604
rect 6092 1556 6144 1562
rect 6092 1498 6144 1504
rect 5632 1420 5684 1426
rect 5632 1362 5684 1368
rect 6000 1420 6052 1426
rect 6000 1362 6052 1368
rect 5538 1320 5594 1329
rect 5538 1255 5594 1264
rect 5644 1018 5672 1362
rect 5632 1012 5684 1018
rect 5632 954 5684 960
rect 5448 944 5500 950
rect 5448 886 5500 892
rect 4988 876 5040 882
rect 4988 818 5040 824
rect 5172 876 5224 882
rect 5172 818 5224 824
rect 3884 808 3936 814
rect 3884 750 3936 756
rect 4528 672 4580 678
rect 4528 614 4580 620
rect 3608 468 3660 474
rect 3608 410 3660 416
rect 3620 270 3648 410
rect 3608 264 3660 270
rect 3608 206 3660 212
rect 4540 202 4568 614
rect 5184 270 5212 818
rect 5356 808 5408 814
rect 5356 750 5408 756
rect 5368 338 5396 750
rect 5460 746 5488 886
rect 5908 808 5960 814
rect 5908 750 5960 756
rect 5448 740 5500 746
rect 5448 682 5500 688
rect 5920 474 5948 750
rect 5908 468 5960 474
rect 5908 410 5960 416
rect 6012 338 6040 1362
rect 6368 808 6420 814
rect 6366 776 6368 785
rect 6420 776 6422 785
rect 6564 746 6592 1838
rect 6656 1290 6684 2042
rect 6644 1284 6696 1290
rect 6644 1226 6696 1232
rect 6642 776 6698 785
rect 6366 711 6422 720
rect 6552 740 6604 746
rect 6748 762 6776 3538
rect 6932 2530 6960 3946
rect 7576 3670 7604 4014
rect 7668 3670 7696 4082
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7576 3466 7604 3606
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 7104 3120 7156 3126
rect 7104 3062 7156 3068
rect 7116 2922 7144 3062
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 6932 2514 7052 2530
rect 6932 2508 7064 2514
rect 6932 2502 7012 2508
rect 6828 2372 6880 2378
rect 6828 2314 6880 2320
rect 6840 2106 6868 2314
rect 6828 2100 6880 2106
rect 6828 2042 6880 2048
rect 6932 1970 6960 2502
rect 7012 2450 7064 2456
rect 7116 2446 7144 2858
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7208 2446 7236 2790
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7012 2372 7064 2378
rect 7012 2314 7064 2320
rect 6920 1964 6972 1970
rect 6920 1906 6972 1912
rect 7024 1902 7052 2314
rect 7300 2122 7328 2994
rect 7392 2310 7420 3402
rect 7760 3292 8068 3312
rect 7760 3290 7766 3292
rect 7822 3290 7846 3292
rect 7902 3290 7926 3292
rect 7982 3290 8006 3292
rect 8062 3290 8068 3292
rect 7822 3238 7824 3290
rect 8004 3238 8006 3290
rect 7760 3236 7766 3238
rect 7822 3236 7846 3238
rect 7902 3236 7926 3238
rect 7982 3236 8006 3238
rect 8062 3236 8068 3238
rect 7760 3216 8068 3236
rect 8220 3058 8248 3402
rect 8404 3398 8432 4490
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8588 4146 8616 4422
rect 8680 4214 8708 5578
rect 8864 5098 8892 7278
rect 9140 6866 9168 7754
rect 9968 7562 9996 7958
rect 10060 7886 10088 8298
rect 10520 7886 10548 8842
rect 10704 8362 10732 9318
rect 11256 9178 11284 10610
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11348 9654 11376 10066
rect 11624 9994 11652 10406
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11808 9722 11836 10610
rect 12410 10364 12718 10384
rect 12410 10362 12416 10364
rect 12472 10362 12496 10364
rect 12552 10362 12576 10364
rect 12632 10362 12656 10364
rect 12712 10362 12718 10364
rect 12472 10310 12474 10362
rect 12654 10310 12656 10362
rect 12410 10308 12416 10310
rect 12472 10308 12496 10310
rect 12552 10308 12576 10310
rect 12632 10308 12656 10310
rect 12712 10308 12718 10310
rect 12410 10288 12718 10308
rect 13556 10266 13584 10678
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13004 10062 13032 10202
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 13004 9722 13032 9998
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 12992 9716 13044 9722
rect 12992 9658 13044 9664
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11612 9648 11664 9654
rect 11612 9590 11664 9596
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 10860 8732 11168 8752
rect 10860 8730 10866 8732
rect 10922 8730 10946 8732
rect 11002 8730 11026 8732
rect 11082 8730 11106 8732
rect 11162 8730 11168 8732
rect 10922 8678 10924 8730
rect 11104 8678 11106 8730
rect 10860 8676 10866 8678
rect 10922 8676 10946 8678
rect 11002 8676 11026 8678
rect 11082 8676 11106 8678
rect 11162 8676 11168 8678
rect 10860 8656 11168 8676
rect 11256 8634 11284 8774
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10060 7750 10088 7822
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10336 7562 10364 7822
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 9968 7534 10364 7562
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9310 7100 9618 7120
rect 9310 7098 9316 7100
rect 9372 7098 9396 7100
rect 9452 7098 9476 7100
rect 9532 7098 9556 7100
rect 9612 7098 9618 7100
rect 9372 7046 9374 7098
rect 9554 7046 9556 7098
rect 9310 7044 9316 7046
rect 9372 7044 9396 7046
rect 9452 7044 9476 7046
rect 9532 7044 9556 7046
rect 9612 7044 9618 7046
rect 9310 7024 9618 7044
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9324 6322 9352 6734
rect 9692 6730 9720 7278
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9692 6322 9720 6666
rect 9968 6390 9996 7210
rect 10336 7002 10364 7534
rect 10428 7410 10456 7686
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 10704 6254 10732 8298
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10796 8022 10824 8230
rect 10784 8016 10836 8022
rect 10784 7958 10836 7964
rect 11348 7936 11376 9590
rect 11624 8974 11652 9590
rect 13188 9382 13216 9862
rect 13740 9586 13768 10474
rect 13924 10062 13952 10474
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14384 10282 14412 10406
rect 14384 10254 14504 10282
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 14476 9994 14504 10254
rect 14464 9988 14516 9994
rect 14464 9930 14516 9936
rect 13960 9820 14268 9840
rect 13960 9818 13966 9820
rect 14022 9818 14046 9820
rect 14102 9818 14126 9820
rect 14182 9818 14206 9820
rect 14262 9818 14268 9820
rect 14022 9766 14024 9818
rect 14204 9766 14206 9818
rect 13960 9764 13966 9766
rect 14022 9764 14046 9766
rect 14102 9764 14126 9766
rect 14182 9764 14206 9766
rect 14262 9764 14268 9766
rect 13960 9744 14268 9764
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 14384 9450 14412 9590
rect 14372 9444 14424 9450
rect 14372 9386 14424 9392
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 12410 9276 12718 9296
rect 12410 9274 12416 9276
rect 12472 9274 12496 9276
rect 12552 9274 12576 9276
rect 12632 9274 12656 9276
rect 12712 9274 12718 9276
rect 12472 9222 12474 9274
rect 12654 9222 12656 9274
rect 12410 9220 12416 9222
rect 12472 9220 12496 9222
rect 12552 9220 12576 9222
rect 12632 9220 12656 9222
rect 12712 9220 12718 9222
rect 12410 9200 12718 9220
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11624 8566 11652 8910
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12268 8634 12296 8774
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11256 7908 11376 7936
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10796 7206 10824 7686
rect 10860 7644 11168 7664
rect 10860 7642 10866 7644
rect 10922 7642 10946 7644
rect 11002 7642 11026 7644
rect 11082 7642 11106 7644
rect 11162 7642 11168 7644
rect 10922 7590 10924 7642
rect 11104 7590 11106 7642
rect 10860 7588 10866 7590
rect 10922 7588 10946 7590
rect 11002 7588 11026 7590
rect 11082 7588 11106 7590
rect 11162 7588 11168 7590
rect 10860 7568 11168 7588
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11164 6934 11192 7142
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8956 5302 8984 6054
rect 9310 6012 9618 6032
rect 9310 6010 9316 6012
rect 9372 6010 9396 6012
rect 9452 6010 9476 6012
rect 9532 6010 9556 6012
rect 9612 6010 9618 6012
rect 9372 5958 9374 6010
rect 9554 5958 9556 6010
rect 9310 5956 9316 5958
rect 9372 5956 9396 5958
rect 9452 5956 9476 5958
rect 9532 5956 9556 5958
rect 9612 5956 9618 5958
rect 9310 5936 9618 5956
rect 10796 5574 10824 6734
rect 10860 6556 11168 6576
rect 10860 6554 10866 6556
rect 10922 6554 10946 6556
rect 11002 6554 11026 6556
rect 11082 6554 11106 6556
rect 11162 6554 11168 6556
rect 10922 6502 10924 6554
rect 11104 6502 11106 6554
rect 10860 6500 10866 6502
rect 10922 6500 10946 6502
rect 11002 6500 11026 6502
rect 11082 6500 11106 6502
rect 11162 6500 11168 6502
rect 10860 6480 11168 6500
rect 11256 5846 11284 7908
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11348 7206 11376 7754
rect 11428 7472 11480 7478
rect 11428 7414 11480 7420
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11440 6322 11468 7414
rect 11624 7018 11652 8502
rect 12544 8498 12572 8774
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12410 8188 12718 8208
rect 12410 8186 12416 8188
rect 12472 8186 12496 8188
rect 12552 8186 12576 8188
rect 12632 8186 12656 8188
rect 12712 8186 12718 8188
rect 12472 8134 12474 8186
rect 12654 8134 12656 8186
rect 12410 8132 12416 8134
rect 12472 8132 12496 8134
rect 12552 8132 12576 8134
rect 12632 8132 12656 8134
rect 12712 8132 12718 8134
rect 12410 8112 12718 8132
rect 12820 8090 12848 9318
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12912 8566 12940 9114
rect 13740 8906 13768 9318
rect 13728 8900 13780 8906
rect 13728 8842 13780 8848
rect 13740 8634 13768 8842
rect 13960 8732 14268 8752
rect 13960 8730 13966 8732
rect 14022 8730 14046 8732
rect 14102 8730 14126 8732
rect 14182 8730 14206 8732
rect 14262 8730 14268 8732
rect 14022 8678 14024 8730
rect 14204 8678 14206 8730
rect 13960 8676 13966 8678
rect 14022 8676 14046 8678
rect 14102 8676 14126 8678
rect 14182 8676 14206 8678
rect 14262 8676 14268 8678
rect 13960 8656 14268 8676
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 14384 8498 14412 9386
rect 14476 9382 14504 9930
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14660 8906 14688 10542
rect 14752 9042 14780 10746
rect 15108 10668 15160 10674
rect 14936 10628 15108 10656
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14844 9518 14872 10406
rect 14936 10198 14964 10628
rect 15108 10610 15160 10616
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 14924 10192 14976 10198
rect 14924 10134 14976 10140
rect 14936 9722 14964 10134
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 14924 9716 14976 9722
rect 14924 9658 14976 9664
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14648 8900 14700 8906
rect 14648 8842 14700 8848
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 13832 8022 13860 8366
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 14476 7954 14504 8774
rect 14568 8498 14596 8774
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12636 7546 12664 7822
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11532 6990 11652 7018
rect 11532 6934 11560 6990
rect 11520 6928 11572 6934
rect 11520 6870 11572 6876
rect 11428 6316 11480 6322
rect 11428 6258 11480 6264
rect 11532 6118 11560 6870
rect 11900 6798 11928 7346
rect 12820 7342 12848 7686
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13188 7410 13216 7482
rect 13563 7472 13615 7478
rect 13450 7440 13506 7449
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13360 7404 13412 7410
rect 13615 7432 13676 7460
rect 13563 7414 13615 7420
rect 13450 7375 13452 7384
rect 13360 7346 13412 7352
rect 13504 7375 13506 7384
rect 13648 7392 13676 7432
rect 13740 7392 13768 7890
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 13960 7644 14268 7664
rect 13960 7642 13966 7644
rect 14022 7642 14046 7644
rect 14102 7642 14126 7644
rect 14182 7642 14206 7644
rect 14262 7642 14268 7644
rect 14022 7590 14024 7642
rect 14204 7590 14206 7642
rect 13960 7588 13966 7590
rect 14022 7588 14046 7590
rect 14102 7588 14126 7590
rect 14182 7588 14206 7590
rect 14262 7588 14268 7590
rect 13960 7568 14268 7588
rect 13648 7364 13768 7392
rect 13452 7346 13504 7352
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12410 7100 12718 7120
rect 12410 7098 12416 7100
rect 12472 7098 12496 7100
rect 12552 7098 12576 7100
rect 12632 7098 12656 7100
rect 12712 7098 12718 7100
rect 12472 7046 12474 7098
rect 12654 7046 12656 7098
rect 12410 7044 12416 7046
rect 12472 7044 12496 7046
rect 12552 7044 12576 7046
rect 12632 7044 12656 7046
rect 12712 7044 12718 7046
rect 12410 7024 12718 7044
rect 11612 6792 11664 6798
rect 11610 6760 11612 6769
rect 11888 6792 11940 6798
rect 11664 6760 11666 6769
rect 11888 6734 11940 6740
rect 11610 6695 11666 6704
rect 11624 6458 11652 6695
rect 12820 6474 12848 7278
rect 12728 6458 12848 6474
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 12716 6452 12848 6458
rect 12768 6446 12848 6452
rect 12716 6394 12768 6400
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11992 5846 12020 6190
rect 12410 6012 12718 6032
rect 12410 6010 12416 6012
rect 12472 6010 12496 6012
rect 12552 6010 12576 6012
rect 12632 6010 12656 6012
rect 12712 6010 12718 6012
rect 12472 5958 12474 6010
rect 12654 5958 12656 6010
rect 12410 5956 12416 5958
rect 12472 5956 12496 5958
rect 12552 5956 12576 5958
rect 12632 5956 12656 5958
rect 12712 5956 12718 5958
rect 12410 5936 12718 5956
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 8944 5296 8996 5302
rect 8944 5238 8996 5244
rect 9048 5234 9076 5510
rect 10796 5370 10824 5510
rect 10860 5468 11168 5488
rect 10860 5466 10866 5468
rect 10922 5466 10946 5468
rect 11002 5466 11026 5468
rect 11082 5466 11106 5468
rect 11162 5466 11168 5468
rect 10922 5414 10924 5466
rect 11104 5414 11106 5466
rect 10860 5412 10866 5414
rect 10922 5412 10946 5414
rect 11002 5412 11026 5414
rect 11082 5412 11106 5414
rect 11162 5412 11168 5414
rect 10860 5392 11168 5412
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 8852 5092 8904 5098
rect 8852 5034 8904 5040
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9232 4554 9260 4966
rect 9310 4924 9618 4944
rect 9310 4922 9316 4924
rect 9372 4922 9396 4924
rect 9452 4922 9476 4924
rect 9532 4922 9556 4924
rect 9612 4922 9618 4924
rect 9372 4870 9374 4922
rect 9554 4870 9556 4922
rect 9310 4868 9316 4870
rect 9372 4868 9396 4870
rect 9452 4868 9476 4870
rect 9532 4868 9556 4870
rect 9612 4868 9618 4870
rect 9310 4848 9618 4868
rect 9968 4690 9996 4966
rect 11164 4826 11192 5102
rect 11256 5030 11284 5782
rect 12912 5778 12940 7346
rect 13266 7304 13322 7313
rect 13372 7290 13400 7346
rect 13372 7274 13676 7290
rect 13372 7268 13688 7274
rect 13372 7262 13636 7268
rect 13266 7239 13268 7248
rect 13320 7239 13322 7248
rect 13268 7210 13320 7216
rect 13636 7210 13688 7216
rect 13740 7206 13768 7364
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 14016 6934 14044 7346
rect 14292 7206 14320 7346
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14384 7002 14412 7754
rect 14556 7472 14608 7478
rect 14554 7440 14556 7449
rect 14608 7440 14610 7449
rect 14554 7375 14610 7384
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14004 6928 14056 6934
rect 14004 6870 14056 6876
rect 14476 6866 14504 7278
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13648 6322 13676 6598
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13740 6118 13768 6802
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 13728 6112 13780 6118
rect 13648 6060 13728 6066
rect 13648 6054 13780 6060
rect 13648 6038 13768 6054
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 13648 5710 13676 6038
rect 13726 5808 13782 5817
rect 13726 5743 13728 5752
rect 13780 5743 13782 5752
rect 13728 5714 13780 5720
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13648 5166 13676 5510
rect 13832 5234 13860 6734
rect 13960 6556 14268 6576
rect 13960 6554 13966 6556
rect 14022 6554 14046 6556
rect 14102 6554 14126 6556
rect 14182 6554 14206 6556
rect 14262 6554 14268 6556
rect 14022 6502 14024 6554
rect 14204 6502 14206 6554
rect 13960 6500 13966 6502
rect 14022 6500 14046 6502
rect 14102 6500 14126 6502
rect 14182 6500 14206 6502
rect 14262 6500 14268 6502
rect 13960 6480 14268 6500
rect 14384 6254 14412 6734
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14384 5778 14412 6190
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14476 5710 14504 6802
rect 14568 6644 14596 7375
rect 14660 6798 14688 8298
rect 14752 7886 14780 8978
rect 14832 8900 14884 8906
rect 14832 8842 14884 8848
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14740 7336 14792 7342
rect 14738 7304 14740 7313
rect 14792 7304 14794 7313
rect 14738 7239 14794 7248
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14648 6656 14700 6662
rect 14568 6616 14648 6644
rect 14648 6598 14700 6604
rect 14660 6322 14688 6598
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 13960 5468 14268 5488
rect 13960 5466 13966 5468
rect 14022 5466 14046 5468
rect 14102 5466 14126 5468
rect 14182 5466 14206 5468
rect 14262 5466 14268 5468
rect 14022 5414 14024 5466
rect 14204 5414 14206 5466
rect 13960 5412 13966 5414
rect 14022 5412 14046 5414
rect 14102 5412 14126 5414
rect 14182 5412 14206 5414
rect 14262 5412 14268 5414
rect 13960 5392 14268 5412
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 13832 5114 13860 5170
rect 13832 5086 13952 5114
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 9956 4684 10008 4690
rect 9876 4644 9956 4672
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 8864 4282 8892 4490
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8668 4208 8720 4214
rect 8668 4150 8720 4156
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 9784 4078 9812 4422
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9310 3836 9618 3856
rect 9310 3834 9316 3836
rect 9372 3834 9396 3836
rect 9452 3834 9476 3836
rect 9532 3834 9556 3836
rect 9612 3834 9618 3836
rect 9372 3782 9374 3834
rect 9554 3782 9556 3834
rect 9310 3780 9316 3782
rect 9372 3780 9396 3782
rect 9452 3780 9476 3782
rect 9532 3780 9556 3782
rect 9612 3780 9618 3782
rect 9310 3760 9618 3780
rect 9784 3534 9812 4014
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 9048 3194 9076 3334
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7484 2650 7512 2926
rect 7668 2650 7696 2994
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 7484 2378 7512 2586
rect 7760 2582 7788 2994
rect 9048 2854 9076 3130
rect 9876 3126 9904 4644
rect 9956 4626 10008 4632
rect 10860 4380 11168 4400
rect 10860 4378 10866 4380
rect 10922 4378 10946 4380
rect 11002 4378 11026 4380
rect 11082 4378 11106 4380
rect 11162 4378 11168 4380
rect 10922 4326 10924 4378
rect 11104 4326 11106 4378
rect 10860 4324 10866 4326
rect 10922 4324 10946 4326
rect 11002 4324 11026 4326
rect 11082 4324 11106 4326
rect 11162 4324 11168 4326
rect 10860 4304 11168 4324
rect 11256 4214 11284 4966
rect 11532 4622 11560 4966
rect 12410 4924 12718 4944
rect 12410 4922 12416 4924
rect 12472 4922 12496 4924
rect 12552 4922 12576 4924
rect 12632 4922 12656 4924
rect 12712 4922 12718 4924
rect 12472 4870 12474 4922
rect 12654 4870 12656 4922
rect 12410 4868 12416 4870
rect 12472 4868 12496 4870
rect 12552 4868 12576 4870
rect 12632 4868 12656 4870
rect 12712 4868 12718 4870
rect 12410 4848 12718 4868
rect 13832 4690 13860 4966
rect 13924 4826 13952 5086
rect 14568 5030 14596 6054
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 11244 4208 11296 4214
rect 11244 4150 11296 4156
rect 11624 4162 11652 4490
rect 11624 4146 11836 4162
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11612 4140 11848 4146
rect 11664 4134 11796 4140
rect 11612 4082 11664 4088
rect 11796 4082 11848 4088
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9968 3738 9996 3946
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 9128 2916 9180 2922
rect 9128 2858 9180 2864
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 8864 2514 8892 2790
rect 8852 2508 8904 2514
rect 8852 2450 8904 2456
rect 8944 2440 8996 2446
rect 7654 2408 7710 2417
rect 7472 2372 7524 2378
rect 9048 2417 9076 2790
rect 9140 2514 9168 2858
rect 9232 2530 9260 3062
rect 9310 2748 9618 2768
rect 9310 2746 9316 2748
rect 9372 2746 9396 2748
rect 9452 2746 9476 2748
rect 9532 2746 9556 2748
rect 9612 2746 9618 2748
rect 9372 2694 9374 2746
rect 9554 2694 9556 2746
rect 9310 2692 9316 2694
rect 9372 2692 9396 2694
rect 9452 2692 9476 2694
rect 9532 2692 9556 2694
rect 9612 2692 9618 2694
rect 9310 2672 9618 2692
rect 9128 2508 9180 2514
rect 9232 2502 9352 2530
rect 9128 2450 9180 2456
rect 8944 2382 8996 2388
rect 9034 2408 9090 2417
rect 7654 2343 7710 2352
rect 7472 2314 7524 2320
rect 7668 2310 7696 2343
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 7300 2106 7420 2122
rect 7288 2100 7420 2106
rect 7340 2094 7420 2100
rect 7288 2042 7340 2048
rect 7104 2032 7156 2038
rect 7104 1974 7156 1980
rect 7012 1896 7064 1902
rect 7012 1838 7064 1844
rect 7116 1766 7144 1974
rect 7288 1964 7340 1970
rect 7288 1906 7340 1912
rect 6828 1760 6880 1766
rect 6828 1702 6880 1708
rect 7104 1760 7156 1766
rect 7104 1702 7156 1708
rect 6840 1358 6868 1702
rect 6828 1352 6880 1358
rect 6828 1294 6880 1300
rect 7116 1222 7144 1702
rect 7104 1216 7156 1222
rect 7104 1158 7156 1164
rect 7116 1018 7144 1158
rect 7104 1012 7156 1018
rect 7104 954 7156 960
rect 7300 882 7328 1906
rect 7392 1426 7420 2094
rect 7668 2038 7696 2246
rect 7760 2204 8068 2224
rect 7760 2202 7766 2204
rect 7822 2202 7846 2204
rect 7902 2202 7926 2204
rect 7982 2202 8006 2204
rect 8062 2202 8068 2204
rect 7822 2150 7824 2202
rect 8004 2150 8006 2202
rect 7760 2148 7766 2150
rect 7822 2148 7846 2150
rect 7902 2148 7926 2150
rect 7982 2148 8006 2150
rect 8062 2148 8068 2150
rect 7760 2128 8068 2148
rect 7656 2032 7708 2038
rect 7656 1974 7708 1980
rect 8300 1896 8352 1902
rect 8300 1838 8352 1844
rect 7380 1420 7432 1426
rect 7380 1362 7432 1368
rect 8312 1358 8340 1838
rect 8772 1358 8800 2246
rect 8956 1952 8984 2382
rect 9034 2343 9090 2352
rect 9218 2408 9274 2417
rect 9218 2343 9220 2352
rect 9272 2343 9274 2352
rect 9220 2314 9272 2320
rect 9324 1970 9352 2502
rect 9036 1964 9088 1970
rect 8956 1924 9036 1952
rect 9036 1906 9088 1912
rect 9312 1964 9364 1970
rect 9312 1906 9364 1912
rect 9588 1964 9640 1970
rect 9588 1906 9640 1912
rect 8300 1352 8352 1358
rect 8300 1294 8352 1300
rect 8668 1352 8720 1358
rect 8668 1294 8720 1300
rect 8760 1352 8812 1358
rect 8760 1294 8812 1300
rect 7760 1116 8068 1136
rect 7760 1114 7766 1116
rect 7822 1114 7846 1116
rect 7902 1114 7926 1116
rect 7982 1114 8006 1116
rect 8062 1114 8068 1116
rect 7822 1062 7824 1114
rect 8004 1062 8006 1114
rect 7760 1060 7766 1062
rect 7822 1060 7846 1062
rect 7902 1060 7926 1062
rect 7982 1060 8006 1062
rect 8062 1060 8068 1062
rect 7760 1040 8068 1060
rect 7288 876 7340 882
rect 7288 818 7340 824
rect 6698 734 6776 762
rect 7748 808 7800 814
rect 7748 750 7800 756
rect 6642 711 6698 720
rect 6552 682 6604 688
rect 6210 572 6518 592
rect 6210 570 6216 572
rect 6272 570 6296 572
rect 6352 570 6376 572
rect 6432 570 6456 572
rect 6512 570 6518 572
rect 6272 518 6274 570
rect 6454 518 6456 570
rect 6210 516 6216 518
rect 6272 516 6296 518
rect 6352 516 6376 518
rect 6432 516 6456 518
rect 6512 516 6518 518
rect 6210 496 6518 516
rect 5356 332 5408 338
rect 5356 274 5408 280
rect 6000 332 6052 338
rect 6000 274 6052 280
rect 5172 264 5224 270
rect 5172 206 5224 212
rect 6656 202 6684 711
rect 6828 672 6880 678
rect 6828 614 6880 620
rect 6840 270 6868 614
rect 7760 474 7788 750
rect 7748 468 7800 474
rect 7748 410 7800 416
rect 8680 270 8708 1294
rect 8760 1216 8812 1222
rect 8760 1158 8812 1164
rect 8772 338 8800 1158
rect 9048 882 9076 1906
rect 9600 1816 9628 1906
rect 9956 1896 10008 1902
rect 9956 1838 10008 1844
rect 9600 1788 9720 1816
rect 9128 1760 9180 1766
rect 9128 1702 9180 1708
rect 9140 1426 9168 1702
rect 9310 1660 9618 1680
rect 9310 1658 9316 1660
rect 9372 1658 9396 1660
rect 9452 1658 9476 1660
rect 9532 1658 9556 1660
rect 9612 1658 9618 1660
rect 9372 1606 9374 1658
rect 9554 1606 9556 1658
rect 9310 1604 9316 1606
rect 9372 1604 9396 1606
rect 9452 1604 9476 1606
rect 9532 1604 9556 1606
rect 9612 1604 9618 1606
rect 9310 1584 9618 1604
rect 9128 1420 9180 1426
rect 9128 1362 9180 1368
rect 9036 876 9088 882
rect 9692 864 9720 1788
rect 9968 1562 9996 1838
rect 9956 1556 10008 1562
rect 9956 1498 10008 1504
rect 10060 1358 10088 4082
rect 10796 3466 10824 4082
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10980 3738 11008 4014
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11440 3466 11468 4082
rect 11624 3670 11652 4082
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11900 3602 11928 3878
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11992 3466 12020 4490
rect 14568 4486 14596 4966
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 12164 4208 12216 4214
rect 12164 4150 12216 4156
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 10336 2650 10364 2790
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10796 2378 10824 3402
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 10860 3292 11168 3312
rect 10860 3290 10866 3292
rect 10922 3290 10946 3292
rect 11002 3290 11026 3292
rect 11082 3290 11106 3292
rect 11162 3290 11168 3292
rect 10922 3238 10924 3290
rect 11104 3238 11106 3290
rect 10860 3236 10866 3238
rect 10922 3236 10946 3238
rect 11002 3236 11026 3238
rect 11082 3236 11106 3238
rect 11162 3236 11168 3238
rect 10860 3216 11168 3236
rect 11348 3194 11376 3334
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 10600 2372 10652 2378
rect 10600 2314 10652 2320
rect 10784 2372 10836 2378
rect 10784 2314 10836 2320
rect 10612 2106 10640 2314
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 10860 2204 11168 2224
rect 10860 2202 10866 2204
rect 10922 2202 10946 2204
rect 11002 2202 11026 2204
rect 11082 2202 11106 2204
rect 11162 2202 11168 2204
rect 10922 2150 10924 2202
rect 11104 2150 11106 2202
rect 10860 2148 10866 2150
rect 10922 2148 10946 2150
rect 11002 2148 11026 2150
rect 11082 2148 11106 2150
rect 11162 2148 11168 2150
rect 10860 2128 11168 2148
rect 11256 2106 11284 2246
rect 10600 2100 10652 2106
rect 10600 2042 10652 2048
rect 11244 2100 11296 2106
rect 11244 2042 11296 2048
rect 10784 1828 10836 1834
rect 10784 1770 10836 1776
rect 10048 1352 10100 1358
rect 10048 1294 10100 1300
rect 10416 1352 10468 1358
rect 10416 1294 10468 1300
rect 10140 1284 10192 1290
rect 10140 1226 10192 1232
rect 9864 876 9916 882
rect 9692 836 9864 864
rect 9036 818 9088 824
rect 9864 818 9916 824
rect 9680 672 9732 678
rect 9680 614 9732 620
rect 9310 572 9618 592
rect 9310 570 9316 572
rect 9372 570 9396 572
rect 9452 570 9476 572
rect 9532 570 9556 572
rect 9612 570 9618 572
rect 9372 518 9374 570
rect 9554 518 9556 570
rect 9310 516 9316 518
rect 9372 516 9396 518
rect 9452 516 9476 518
rect 9532 516 9556 518
rect 9612 516 9618 518
rect 9310 496 9618 516
rect 9692 338 9720 614
rect 10152 338 10180 1226
rect 10324 1216 10376 1222
rect 10324 1158 10376 1164
rect 10336 1018 10364 1158
rect 10324 1012 10376 1018
rect 10324 954 10376 960
rect 10428 950 10456 1294
rect 10416 944 10468 950
rect 10416 886 10468 892
rect 8760 332 8812 338
rect 8760 274 8812 280
rect 9680 332 9732 338
rect 9680 274 9732 280
rect 10140 332 10192 338
rect 10140 274 10192 280
rect 10428 270 10456 886
rect 10508 876 10560 882
rect 10508 818 10560 824
rect 10520 474 10548 818
rect 10796 796 10824 1770
rect 11152 1760 11204 1766
rect 11152 1702 11204 1708
rect 11164 1358 11192 1702
rect 11152 1352 11204 1358
rect 11152 1294 11204 1300
rect 10860 1116 11168 1136
rect 10860 1114 10866 1116
rect 10922 1114 10946 1116
rect 11002 1114 11026 1116
rect 11082 1114 11106 1116
rect 11162 1114 11168 1116
rect 10922 1062 10924 1114
rect 11104 1062 11106 1114
rect 10860 1060 10866 1062
rect 10922 1060 10946 1062
rect 11002 1060 11026 1062
rect 11082 1060 11106 1062
rect 11162 1060 11168 1062
rect 10860 1040 11168 1060
rect 11348 1018 11376 3130
rect 11888 2576 11940 2582
rect 11888 2518 11940 2524
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 11532 1426 11560 2450
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 11520 1420 11572 1426
rect 11520 1362 11572 1368
rect 11336 1012 11388 1018
rect 11336 954 11388 960
rect 11624 882 11652 2314
rect 11796 1216 11848 1222
rect 11796 1158 11848 1164
rect 11808 950 11836 1158
rect 11796 944 11848 950
rect 11794 912 11796 921
rect 11848 912 11850 921
rect 10968 876 11020 882
rect 10968 818 11020 824
rect 11612 876 11664 882
rect 11900 882 11928 2518
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11992 2038 12020 2246
rect 11980 2032 12032 2038
rect 11980 1974 12032 1980
rect 11992 1562 12020 1974
rect 11980 1556 12032 1562
rect 11980 1498 12032 1504
rect 11794 847 11850 856
rect 11888 876 11940 882
rect 11612 818 11664 824
rect 11888 818 11940 824
rect 12072 876 12124 882
rect 12176 864 12204 4150
rect 12268 4146 12296 4422
rect 13188 4214 13216 4422
rect 13960 4380 14268 4400
rect 13960 4378 13966 4380
rect 14022 4378 14046 4380
rect 14102 4378 14126 4380
rect 14182 4378 14206 4380
rect 14262 4378 14268 4380
rect 14022 4326 14024 4378
rect 14204 4326 14206 4378
rect 13960 4324 13966 4326
rect 14022 4324 14046 4326
rect 14102 4324 14126 4326
rect 14182 4324 14206 4326
rect 14262 4324 14268 4326
rect 13960 4304 14268 4324
rect 14568 4214 14596 4422
rect 14740 4276 14792 4282
rect 14740 4218 14792 4224
rect 13176 4208 13228 4214
rect 13176 4150 13228 4156
rect 14556 4208 14608 4214
rect 14556 4150 14608 4156
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12410 3836 12718 3856
rect 12410 3834 12416 3836
rect 12472 3834 12496 3836
rect 12552 3834 12576 3836
rect 12632 3834 12656 3836
rect 12712 3834 12718 3836
rect 12472 3782 12474 3834
rect 12654 3782 12656 3834
rect 12410 3780 12416 3782
rect 12472 3780 12496 3782
rect 12552 3780 12576 3782
rect 12632 3780 12656 3782
rect 12712 3780 12718 3782
rect 12410 3760 12718 3780
rect 12820 3738 12848 4014
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 13188 3398 13216 4150
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13648 3466 13676 3538
rect 13740 3534 13768 3878
rect 13832 3534 13860 4014
rect 14752 3738 14780 4218
rect 14844 4078 14872 8842
rect 14936 8090 14964 9658
rect 15028 9042 15056 10066
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15212 9518 15240 9862
rect 15304 9586 15332 10610
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15016 8900 15068 8906
rect 15016 8842 15068 8848
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14936 5234 14964 7686
rect 15028 6769 15056 8842
rect 15120 8430 15148 8910
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15304 8498 15332 8774
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15120 7954 15148 8366
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15014 6760 15070 6769
rect 15014 6695 15070 6704
rect 15028 5574 15056 6695
rect 15120 6390 15148 7890
rect 15304 7750 15332 8434
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15304 6798 15332 7142
rect 15292 6792 15344 6798
rect 15212 6740 15292 6746
rect 15212 6734 15344 6740
rect 15212 6718 15332 6734
rect 15212 6662 15240 6718
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15304 5778 15332 6054
rect 15396 5914 15424 11206
rect 15580 11098 15608 11206
rect 15658 11200 15714 12000
rect 18510 11200 18566 12000
rect 18786 11248 18842 11257
rect 15672 11098 15700 11200
rect 15580 11070 15700 11098
rect 17060 10908 17368 10928
rect 17060 10906 17066 10908
rect 17122 10906 17146 10908
rect 17202 10906 17226 10908
rect 17282 10906 17306 10908
rect 17362 10906 17368 10908
rect 17122 10854 17124 10906
rect 17304 10854 17306 10906
rect 17060 10852 17066 10854
rect 17122 10852 17146 10854
rect 17202 10852 17226 10854
rect 17282 10852 17306 10854
rect 17362 10852 17368 10854
rect 17060 10832 17368 10852
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 15510 10364 15818 10384
rect 15510 10362 15516 10364
rect 15572 10362 15596 10364
rect 15652 10362 15676 10364
rect 15732 10362 15756 10364
rect 15812 10362 15818 10364
rect 15572 10310 15574 10362
rect 15754 10310 15756 10362
rect 15510 10308 15516 10310
rect 15572 10308 15596 10310
rect 15652 10308 15676 10310
rect 15732 10308 15756 10310
rect 15812 10308 15818 10310
rect 15510 10288 15818 10308
rect 16224 9654 16252 10406
rect 18064 10266 18092 10610
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16592 9654 16620 10066
rect 16764 9988 16816 9994
rect 16764 9930 16816 9936
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16776 9586 16804 9930
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 17060 9820 17368 9840
rect 17060 9818 17066 9820
rect 17122 9818 17146 9820
rect 17202 9818 17226 9820
rect 17282 9818 17306 9820
rect 17362 9818 17368 9820
rect 17122 9766 17124 9818
rect 17304 9766 17306 9818
rect 17060 9764 17066 9766
rect 17122 9764 17146 9766
rect 17202 9764 17226 9766
rect 17282 9764 17306 9766
rect 17362 9764 17368 9766
rect 17060 9744 17368 9764
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 15510 9276 15818 9296
rect 15510 9274 15516 9276
rect 15572 9274 15596 9276
rect 15652 9274 15676 9276
rect 15732 9274 15756 9276
rect 15812 9274 15818 9276
rect 15572 9222 15574 9274
rect 15754 9222 15756 9274
rect 15510 9220 15516 9222
rect 15572 9220 15596 9222
rect 15652 9220 15676 9222
rect 15732 9220 15756 9222
rect 15812 9220 15818 9222
rect 15510 9200 15818 9220
rect 16776 8906 16804 9522
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 16120 8900 16172 8906
rect 16120 8842 16172 8848
rect 16764 8900 16816 8906
rect 16764 8842 16816 8848
rect 16132 8634 16160 8842
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16776 8566 16804 8842
rect 17060 8732 17368 8752
rect 17060 8730 17066 8732
rect 17122 8730 17146 8732
rect 17202 8730 17226 8732
rect 17282 8730 17306 8732
rect 17362 8730 17368 8732
rect 17122 8678 17124 8730
rect 17304 8678 17306 8730
rect 17060 8676 17066 8678
rect 17122 8676 17146 8678
rect 17202 8676 17226 8678
rect 17282 8676 17306 8678
rect 17362 8676 17368 8678
rect 17060 8656 17368 8676
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 16580 8288 16632 8294
rect 16580 8230 16632 8236
rect 15510 8188 15818 8208
rect 15510 8186 15516 8188
rect 15572 8186 15596 8188
rect 15652 8186 15676 8188
rect 15732 8186 15756 8188
rect 15812 8186 15818 8188
rect 15572 8134 15574 8186
rect 15754 8134 15756 8186
rect 15510 8132 15516 8134
rect 15572 8132 15596 8134
rect 15652 8132 15676 8134
rect 15732 8132 15756 8134
rect 15812 8132 15818 8134
rect 15510 8112 15818 8132
rect 16592 7954 16620 8230
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15510 7100 15818 7120
rect 15510 7098 15516 7100
rect 15572 7098 15596 7100
rect 15652 7098 15676 7100
rect 15732 7098 15756 7100
rect 15812 7098 15818 7100
rect 15572 7046 15574 7098
rect 15754 7046 15756 7098
rect 15510 7044 15516 7046
rect 15572 7044 15596 7046
rect 15652 7044 15676 7046
rect 15732 7044 15756 7046
rect 15812 7044 15818 7046
rect 15510 7024 15818 7044
rect 15856 6798 15884 7822
rect 16776 7750 16804 8502
rect 17512 7954 17540 9318
rect 18340 9178 18368 9862
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 18524 8514 18552 11200
rect 18786 11183 18842 11192
rect 18800 10674 18828 11183
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18616 9761 18644 9998
rect 18602 9752 18658 9761
rect 18602 9687 18658 9696
rect 18432 8486 18552 8514
rect 18604 8492 18656 8498
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16776 7478 16804 7686
rect 17060 7644 17368 7664
rect 17060 7642 17066 7644
rect 17122 7642 17146 7644
rect 17202 7642 17226 7644
rect 17282 7642 17306 7644
rect 17362 7642 17368 7644
rect 17122 7590 17124 7642
rect 17304 7590 17306 7642
rect 17060 7588 17066 7590
rect 17122 7588 17146 7590
rect 17202 7588 17226 7590
rect 17282 7588 17306 7590
rect 17362 7588 17368 7590
rect 17060 7568 17368 7588
rect 16764 7472 16816 7478
rect 16764 7414 16816 7420
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 16212 6724 16264 6730
rect 16212 6666 16264 6672
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 15856 6458 15884 6598
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 16224 6322 16252 6666
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 15510 6012 15818 6032
rect 15510 6010 15516 6012
rect 15572 6010 15596 6012
rect 15652 6010 15676 6012
rect 15732 6010 15756 6012
rect 15812 6010 15818 6012
rect 15572 5958 15574 6010
rect 15754 5958 15756 6010
rect 15510 5956 15516 5958
rect 15572 5956 15596 5958
rect 15652 5956 15676 5958
rect 15732 5956 15756 5958
rect 15812 5956 15818 5958
rect 15510 5936 15818 5956
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 16592 5778 16620 7142
rect 16672 6996 16724 7002
rect 16672 6938 16724 6944
rect 16684 6458 16712 6938
rect 16776 6730 16804 7414
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16776 6338 16804 6666
rect 16868 6458 16896 7346
rect 17408 6724 17460 6730
rect 17408 6666 17460 6672
rect 17060 6556 17368 6576
rect 17060 6554 17066 6556
rect 17122 6554 17146 6556
rect 17202 6554 17226 6556
rect 17282 6554 17306 6556
rect 17362 6554 17368 6556
rect 17122 6502 17124 6554
rect 17304 6502 17306 6554
rect 17060 6500 17066 6502
rect 17122 6500 17146 6502
rect 17202 6500 17226 6502
rect 17282 6500 17306 6502
rect 17362 6500 17368 6502
rect 17060 6480 17368 6500
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16684 6322 16804 6338
rect 16672 6316 16804 6322
rect 16724 6310 16804 6316
rect 16948 6316 17000 6322
rect 16672 6258 16724 6264
rect 16948 6258 17000 6264
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14648 3596 14700 3602
rect 14648 3538 14700 3544
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 12410 2748 12718 2768
rect 12410 2746 12416 2748
rect 12472 2746 12496 2748
rect 12552 2746 12576 2748
rect 12632 2746 12656 2748
rect 12712 2746 12718 2748
rect 12472 2694 12474 2746
rect 12654 2694 12656 2746
rect 12410 2692 12416 2694
rect 12472 2692 12496 2694
rect 12552 2692 12576 2694
rect 12632 2692 12656 2694
rect 12712 2692 12718 2694
rect 12410 2672 12718 2692
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 12268 1902 12296 2450
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12360 2310 12388 2382
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 12636 2106 12664 2382
rect 12624 2100 12676 2106
rect 12624 2042 12676 2048
rect 12820 1970 12848 2994
rect 13004 2582 13032 3130
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 12900 2576 12952 2582
rect 12900 2518 12952 2524
rect 12992 2576 13044 2582
rect 12992 2518 13044 2524
rect 12912 2394 12940 2518
rect 13556 2428 13584 2994
rect 13648 2774 13676 3402
rect 13648 2746 13768 2774
rect 13636 2440 13688 2446
rect 13556 2400 13636 2428
rect 12912 2378 13216 2394
rect 13636 2382 13688 2388
rect 12912 2372 13228 2378
rect 12912 2366 13176 2372
rect 13176 2314 13228 2320
rect 12808 1964 12860 1970
rect 12808 1906 12860 1912
rect 12256 1896 12308 1902
rect 12256 1838 12308 1844
rect 12992 1760 13044 1766
rect 12992 1702 13044 1708
rect 12410 1660 12718 1680
rect 12410 1658 12416 1660
rect 12472 1658 12496 1660
rect 12552 1658 12576 1660
rect 12632 1658 12656 1660
rect 12712 1658 12718 1660
rect 12472 1606 12474 1658
rect 12654 1606 12656 1658
rect 12410 1604 12416 1606
rect 12472 1604 12496 1606
rect 12552 1604 12576 1606
rect 12632 1604 12656 1606
rect 12712 1604 12718 1606
rect 12410 1584 12718 1604
rect 13004 1426 13032 1702
rect 12992 1420 13044 1426
rect 12992 1362 13044 1368
rect 13740 1358 13768 2746
rect 13832 2514 13860 3470
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 13960 3292 14268 3312
rect 13960 3290 13966 3292
rect 14022 3290 14046 3292
rect 14102 3290 14126 3292
rect 14182 3290 14206 3292
rect 14262 3290 14268 3292
rect 14022 3238 14024 3290
rect 14204 3238 14206 3290
rect 13960 3236 13966 3238
rect 14022 3236 14046 3238
rect 14102 3236 14126 3238
rect 14182 3236 14206 3238
rect 14262 3236 14268 3238
rect 13960 3216 14268 3236
rect 14384 3058 14412 3334
rect 14660 3194 14688 3538
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 14752 3058 14780 3674
rect 14936 3670 14964 5170
rect 15396 4706 15424 5646
rect 16684 5574 16712 6258
rect 16960 5914 16988 6258
rect 17420 6254 17448 6666
rect 18064 6458 18092 7890
rect 18432 6866 18460 8486
rect 18604 8434 18656 8440
rect 18616 8265 18644 8434
rect 18602 8256 18658 8265
rect 18602 8191 18658 8200
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18512 6792 18564 6798
rect 18510 6760 18512 6769
rect 18564 6760 18566 6769
rect 18510 6695 18566 6704
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17500 6248 17552 6254
rect 17500 6190 17552 6196
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 15672 5302 15700 5510
rect 15660 5296 15712 5302
rect 15660 5238 15712 5244
rect 16960 5234 16988 5850
rect 17420 5817 17448 6190
rect 17406 5808 17462 5817
rect 17406 5743 17462 5752
rect 17060 5468 17368 5488
rect 17060 5466 17066 5468
rect 17122 5466 17146 5468
rect 17202 5466 17226 5468
rect 17282 5466 17306 5468
rect 17362 5466 17368 5468
rect 17122 5414 17124 5466
rect 17304 5414 17306 5466
rect 17060 5412 17066 5414
rect 17122 5412 17146 5414
rect 17202 5412 17226 5414
rect 17282 5412 17306 5414
rect 17362 5412 17368 5414
rect 17060 5392 17368 5412
rect 17512 5302 17540 6190
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18328 5568 18380 5574
rect 18328 5510 18380 5516
rect 17500 5296 17552 5302
rect 17500 5238 17552 5244
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 18340 5166 18368 5510
rect 18524 5273 18552 5646
rect 18510 5264 18566 5273
rect 18510 5199 18566 5208
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 15510 4924 15818 4944
rect 15510 4922 15516 4924
rect 15572 4922 15596 4924
rect 15652 4922 15676 4924
rect 15732 4922 15756 4924
rect 15812 4922 15818 4924
rect 15572 4870 15574 4922
rect 15754 4870 15756 4922
rect 15510 4868 15516 4870
rect 15572 4868 15596 4870
rect 15652 4868 15676 4870
rect 15732 4868 15756 4870
rect 15812 4868 15818 4870
rect 15510 4848 15818 4868
rect 15396 4690 15516 4706
rect 16868 4690 16896 4966
rect 15396 4684 15528 4690
rect 15396 4678 15476 4684
rect 15476 4626 15528 4632
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 15200 4548 15252 4554
rect 15200 4490 15252 4496
rect 14924 3664 14976 3670
rect 14924 3606 14976 3612
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14568 2650 14596 2994
rect 14936 2990 14964 3606
rect 15108 3392 15160 3398
rect 15108 3334 15160 3340
rect 15120 3126 15148 3334
rect 15108 3120 15160 3126
rect 15108 3062 15160 3068
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 15108 2984 15160 2990
rect 15108 2926 15160 2932
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 14568 2378 14596 2586
rect 14556 2372 14608 2378
rect 14556 2314 14608 2320
rect 13960 2204 14268 2224
rect 13960 2202 13966 2204
rect 14022 2202 14046 2204
rect 14102 2202 14126 2204
rect 14182 2202 14206 2204
rect 14262 2202 14268 2204
rect 14022 2150 14024 2202
rect 14204 2150 14206 2202
rect 13960 2148 13966 2150
rect 14022 2148 14046 2150
rect 14102 2148 14126 2150
rect 14182 2148 14206 2150
rect 14262 2148 14268 2150
rect 13960 2128 14268 2148
rect 14568 2106 14596 2314
rect 14648 2304 14700 2310
rect 14648 2246 14700 2252
rect 14556 2100 14608 2106
rect 14556 2042 14608 2048
rect 14464 1964 14516 1970
rect 14568 1952 14596 2042
rect 14660 1970 14688 2246
rect 14516 1924 14596 1952
rect 14648 1964 14700 1970
rect 14464 1906 14516 1912
rect 14924 1964 14976 1970
rect 14700 1924 14780 1952
rect 14648 1906 14700 1912
rect 14648 1828 14700 1834
rect 14648 1770 14700 1776
rect 14188 1760 14240 1766
rect 14188 1702 14240 1708
rect 14200 1562 14228 1702
rect 14188 1556 14240 1562
rect 14188 1498 14240 1504
rect 14464 1488 14516 1494
rect 14464 1430 14516 1436
rect 13728 1352 13780 1358
rect 13728 1294 13780 1300
rect 13360 1284 13412 1290
rect 13360 1226 13412 1232
rect 12256 1216 12308 1222
rect 12256 1158 12308 1164
rect 12124 836 12204 864
rect 12072 818 12124 824
rect 10876 808 10928 814
rect 10796 768 10876 796
rect 10980 785 11008 818
rect 10876 750 10928 756
rect 10966 776 11022 785
rect 10966 711 11022 720
rect 12164 672 12216 678
rect 12164 614 12216 620
rect 10508 468 10560 474
rect 10508 410 10560 416
rect 12176 338 12204 614
rect 12268 338 12296 1158
rect 13372 1018 13400 1226
rect 13636 1216 13688 1222
rect 13636 1158 13688 1164
rect 13648 1018 13676 1158
rect 13960 1116 14268 1136
rect 13960 1114 13966 1116
rect 14022 1114 14046 1116
rect 14102 1114 14126 1116
rect 14182 1114 14206 1116
rect 14262 1114 14268 1116
rect 14022 1062 14024 1114
rect 14204 1062 14206 1114
rect 13960 1060 13966 1062
rect 14022 1060 14046 1062
rect 14102 1060 14126 1062
rect 14182 1060 14206 1062
rect 14262 1060 14268 1062
rect 13960 1040 14268 1060
rect 13360 1012 13412 1018
rect 13360 954 13412 960
rect 13636 1012 13688 1018
rect 13636 954 13688 960
rect 14476 950 14504 1430
rect 14464 944 14516 950
rect 13818 912 13874 921
rect 14464 886 14516 892
rect 13818 847 13874 856
rect 13832 814 13860 847
rect 12808 808 12860 814
rect 12808 750 12860 756
rect 13820 808 13872 814
rect 13820 750 13872 756
rect 12410 572 12718 592
rect 12410 570 12416 572
rect 12472 570 12496 572
rect 12552 570 12576 572
rect 12632 570 12656 572
rect 12712 570 12718 572
rect 12472 518 12474 570
rect 12654 518 12656 570
rect 12410 516 12416 518
rect 12472 516 12496 518
rect 12552 516 12576 518
rect 12632 516 12656 518
rect 12712 516 12718 518
rect 12410 496 12718 516
rect 12820 474 12848 750
rect 14660 474 14688 1770
rect 14752 1358 14780 1924
rect 14924 1906 14976 1912
rect 14936 1426 14964 1906
rect 15120 1834 15148 2926
rect 15212 2650 15240 4490
rect 17060 4380 17368 4400
rect 17060 4378 17066 4380
rect 17122 4378 17146 4380
rect 17202 4378 17226 4380
rect 17282 4378 17306 4380
rect 17362 4378 17368 4380
rect 17122 4326 17124 4378
rect 17304 4326 17306 4378
rect 17060 4324 17066 4326
rect 17122 4324 17146 4326
rect 17202 4324 17226 4326
rect 17282 4324 17306 4326
rect 17362 4324 17368 4326
rect 17060 4304 17368 4324
rect 15476 4072 15528 4078
rect 15304 4032 15476 4060
rect 15304 3534 15332 4032
rect 15476 4014 15528 4020
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 15510 3836 15818 3856
rect 15510 3834 15516 3836
rect 15572 3834 15596 3836
rect 15652 3834 15676 3836
rect 15732 3834 15756 3836
rect 15812 3834 15818 3836
rect 15572 3782 15574 3834
rect 15754 3782 15756 3834
rect 15510 3780 15516 3782
rect 15572 3780 15596 3782
rect 15652 3780 15676 3782
rect 15732 3780 15756 3782
rect 15812 3780 15818 3782
rect 15510 3760 15818 3780
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15304 1970 15332 3470
rect 15764 3074 15792 3470
rect 15856 3194 15884 3470
rect 17060 3292 17368 3312
rect 17060 3290 17066 3292
rect 17122 3290 17146 3292
rect 17202 3290 17226 3292
rect 17282 3290 17306 3292
rect 17362 3290 17368 3292
rect 17122 3238 17124 3290
rect 17304 3238 17306 3290
rect 17060 3236 17066 3238
rect 17122 3236 17146 3238
rect 17202 3236 17226 3238
rect 17282 3236 17306 3238
rect 17362 3236 17368 3238
rect 17060 3216 17368 3236
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 15384 3052 15436 3058
rect 15764 3046 15884 3074
rect 15384 2994 15436 3000
rect 15396 2310 15424 2994
rect 15856 2990 15884 3046
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15510 2748 15818 2768
rect 15510 2746 15516 2748
rect 15572 2746 15596 2748
rect 15652 2746 15676 2748
rect 15732 2746 15756 2748
rect 15812 2746 15818 2748
rect 15572 2694 15574 2746
rect 15754 2694 15756 2746
rect 15510 2692 15516 2694
rect 15572 2692 15596 2694
rect 15652 2692 15676 2694
rect 15732 2692 15756 2694
rect 15812 2692 15818 2694
rect 15510 2672 15818 2692
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 15292 1964 15344 1970
rect 15292 1906 15344 1912
rect 15200 1896 15252 1902
rect 15200 1838 15252 1844
rect 15108 1828 15160 1834
rect 15108 1770 15160 1776
rect 15212 1426 15240 1838
rect 14924 1420 14976 1426
rect 14924 1362 14976 1368
rect 15200 1420 15252 1426
rect 15200 1362 15252 1368
rect 14740 1352 14792 1358
rect 14740 1294 14792 1300
rect 14924 1284 14976 1290
rect 14924 1226 14976 1232
rect 14936 950 14964 1226
rect 15304 1018 15332 1906
rect 15396 1290 15424 2246
rect 15510 1660 15818 1680
rect 15510 1658 15516 1660
rect 15572 1658 15596 1660
rect 15652 1658 15676 1660
rect 15732 1658 15756 1660
rect 15812 1658 15818 1660
rect 15572 1606 15574 1658
rect 15754 1606 15756 1658
rect 15510 1604 15516 1606
rect 15572 1604 15596 1606
rect 15652 1604 15676 1606
rect 15732 1604 15756 1606
rect 15812 1604 15818 1606
rect 15510 1584 15818 1604
rect 15856 1358 15884 2926
rect 16948 2508 17000 2514
rect 16948 2450 17000 2456
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16132 1426 16160 2246
rect 16960 2106 16988 2450
rect 17592 2372 17644 2378
rect 17592 2314 17644 2320
rect 17060 2204 17368 2224
rect 17060 2202 17066 2204
rect 17122 2202 17146 2204
rect 17202 2202 17226 2204
rect 17282 2202 17306 2204
rect 17362 2202 17368 2204
rect 17122 2150 17124 2202
rect 17304 2150 17306 2202
rect 17060 2148 17066 2150
rect 17122 2148 17146 2150
rect 17202 2148 17226 2150
rect 17282 2148 17306 2150
rect 17362 2148 17368 2150
rect 17060 2128 17368 2148
rect 16948 2100 17000 2106
rect 16948 2042 17000 2048
rect 16488 1964 16540 1970
rect 16540 1924 16620 1952
rect 16488 1906 16540 1912
rect 16120 1420 16172 1426
rect 16120 1362 16172 1368
rect 15844 1352 15896 1358
rect 15844 1294 15896 1300
rect 15384 1284 15436 1290
rect 15384 1226 15436 1232
rect 15292 1012 15344 1018
rect 15292 954 15344 960
rect 14924 944 14976 950
rect 14924 886 14976 892
rect 16212 808 16264 814
rect 16212 750 16264 756
rect 15510 572 15818 592
rect 15510 570 15516 572
rect 15572 570 15596 572
rect 15652 570 15676 572
rect 15732 570 15756 572
rect 15812 570 15818 572
rect 15572 518 15574 570
rect 15754 518 15756 570
rect 15510 516 15516 518
rect 15572 516 15596 518
rect 15652 516 15676 518
rect 15732 516 15756 518
rect 15812 516 15818 518
rect 15510 496 15818 516
rect 16224 474 16252 750
rect 16592 474 16620 1924
rect 16672 1760 16724 1766
rect 16672 1702 16724 1708
rect 12808 468 12860 474
rect 12808 410 12860 416
rect 14648 468 14700 474
rect 14648 410 14700 416
rect 16212 468 16264 474
rect 16212 410 16264 416
rect 16580 468 16632 474
rect 16580 410 16632 416
rect 14646 368 14702 377
rect 12164 332 12216 338
rect 12164 274 12216 280
rect 12256 332 12308 338
rect 12256 274 12308 280
rect 12624 332 12676 338
rect 14646 303 14702 312
rect 12624 274 12676 280
rect 6828 264 6880 270
rect 8668 264 8720 270
rect 6828 206 6880 212
rect 8666 232 8668 241
rect 10416 264 10468 270
rect 8720 232 8722 241
rect 3516 196 3568 202
rect 3516 138 3568 144
rect 4528 196 4580 202
rect 4528 138 4580 144
rect 6644 196 6696 202
rect 12636 241 12664 274
rect 14660 270 14688 303
rect 16684 270 16712 1702
rect 16960 950 16988 2042
rect 17604 1562 17632 2314
rect 17592 1556 17644 1562
rect 17592 1498 17644 1504
rect 17788 1358 17816 3878
rect 17880 2990 17908 4558
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 17868 2984 17920 2990
rect 17868 2926 17920 2932
rect 17880 2514 17908 2926
rect 17868 2508 17920 2514
rect 17868 2450 17920 2456
rect 17776 1352 17828 1358
rect 17776 1294 17828 1300
rect 17868 1352 17920 1358
rect 17868 1294 17920 1300
rect 18052 1352 18104 1358
rect 18052 1294 18104 1300
rect 17060 1116 17368 1136
rect 17060 1114 17066 1116
rect 17122 1114 17146 1116
rect 17202 1114 17226 1116
rect 17282 1114 17306 1116
rect 17362 1114 17368 1116
rect 17122 1062 17124 1114
rect 17304 1062 17306 1114
rect 17060 1060 17066 1062
rect 17122 1060 17146 1062
rect 17202 1060 17226 1062
rect 17282 1060 17306 1062
rect 17362 1060 17368 1062
rect 17060 1040 17368 1060
rect 16948 944 17000 950
rect 16948 886 17000 892
rect 17880 746 17908 1294
rect 17960 1216 18012 1222
rect 17960 1158 18012 1164
rect 17868 740 17920 746
rect 17868 682 17920 688
rect 17972 377 18000 1158
rect 18064 474 18092 1294
rect 18156 785 18184 3470
rect 18340 3058 18368 3878
rect 18524 3777 18552 4082
rect 18510 3768 18566 3777
rect 18510 3703 18566 3712
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18524 2281 18552 2382
rect 18510 2272 18566 2281
rect 18510 2207 18566 2216
rect 18420 1352 18472 1358
rect 18420 1294 18472 1300
rect 18236 1284 18288 1290
rect 18236 1226 18288 1232
rect 18248 1018 18276 1226
rect 18236 1012 18288 1018
rect 18236 954 18288 960
rect 18142 776 18198 785
rect 18142 711 18198 720
rect 18052 468 18104 474
rect 18052 410 18104 416
rect 17958 368 18014 377
rect 17958 303 18014 312
rect 18156 270 18184 711
rect 18432 474 18460 1294
rect 18512 1216 18564 1222
rect 18512 1158 18564 1164
rect 18524 882 18552 1158
rect 18512 876 18564 882
rect 18512 818 18564 824
rect 18524 785 18552 818
rect 18510 776 18566 785
rect 18510 711 18566 720
rect 18420 468 18472 474
rect 18420 410 18472 416
rect 14648 264 14700 270
rect 10416 206 10468 212
rect 12622 232 12678 241
rect 8666 167 8722 176
rect 14648 206 14700 212
rect 16672 264 16724 270
rect 16672 206 16724 212
rect 18144 264 18196 270
rect 18144 206 18196 212
rect 12622 167 12678 176
rect 6644 138 6696 144
rect 4660 28 4968 48
rect 4660 26 4666 28
rect 4722 26 4746 28
rect 4802 26 4826 28
rect 4882 26 4906 28
rect 4962 26 4968 28
rect 4722 -26 4724 26
rect 4904 -26 4906 26
rect 4660 -28 4666 -26
rect 4722 -28 4746 -26
rect 4802 -28 4826 -26
rect 4882 -28 4906 -26
rect 4962 -28 4968 -26
rect 4660 -48 4968 -28
rect 7760 28 8068 48
rect 7760 26 7766 28
rect 7822 26 7846 28
rect 7902 26 7926 28
rect 7982 26 8006 28
rect 8062 26 8068 28
rect 7822 -26 7824 26
rect 8004 -26 8006 26
rect 7760 -28 7766 -26
rect 7822 -28 7846 -26
rect 7902 -28 7926 -26
rect 7982 -28 8006 -26
rect 8062 -28 8068 -26
rect 7760 -48 8068 -28
rect 10860 28 11168 48
rect 10860 26 10866 28
rect 10922 26 10946 28
rect 11002 26 11026 28
rect 11082 26 11106 28
rect 11162 26 11168 28
rect 10922 -26 10924 26
rect 11104 -26 11106 26
rect 10860 -28 10866 -26
rect 10922 -28 10946 -26
rect 11002 -28 11026 -26
rect 11082 -28 11106 -26
rect 11162 -28 11168 -26
rect 10860 -48 11168 -28
rect 13960 28 14268 48
rect 13960 26 13966 28
rect 14022 26 14046 28
rect 14102 26 14126 28
rect 14182 26 14206 28
rect 14262 26 14268 28
rect 14022 -26 14024 26
rect 14204 -26 14206 26
rect 13960 -28 13966 -26
rect 14022 -28 14046 -26
rect 14102 -28 14126 -26
rect 14182 -28 14206 -26
rect 14262 -28 14268 -26
rect 13960 -48 14268 -28
rect 17060 28 17368 48
rect 17060 26 17066 28
rect 17122 26 17146 28
rect 17202 26 17226 28
rect 17282 26 17306 28
rect 17362 26 17368 28
rect 17122 -26 17124 26
rect 17304 -26 17306 26
rect 17060 -28 17066 -26
rect 17122 -28 17146 -26
rect 17202 -28 17226 -26
rect 17282 -28 17306 -26
rect 17362 -28 17368 -26
rect 17060 -48 17368 -28
<< via2 >>
rect 2410 9424 2466 9480
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 3276 10362 3332 10364
rect 3356 10362 3412 10364
rect 3116 10310 3162 10362
rect 3162 10310 3172 10362
rect 3196 10310 3226 10362
rect 3226 10310 3238 10362
rect 3238 10310 3252 10362
rect 3276 10310 3290 10362
rect 3290 10310 3302 10362
rect 3302 10310 3332 10362
rect 3356 10310 3366 10362
rect 3366 10310 3412 10362
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 3276 10308 3332 10310
rect 3356 10308 3412 10310
rect 3146 10104 3202 10160
rect 3238 9968 3294 10024
rect 3330 9460 3332 9480
rect 3332 9460 3384 9480
rect 3384 9460 3386 9480
rect 3330 9424 3386 9460
rect 3974 10124 4030 10160
rect 3974 10104 3976 10124
rect 3976 10104 4028 10124
rect 4028 10104 4030 10124
rect 3974 9988 4030 10024
rect 3974 9968 3976 9988
rect 3976 9968 4028 9988
rect 4028 9968 4030 9988
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 3276 9274 3332 9276
rect 3356 9274 3412 9276
rect 3116 9222 3162 9274
rect 3162 9222 3172 9274
rect 3196 9222 3226 9274
rect 3226 9222 3238 9274
rect 3238 9222 3252 9274
rect 3276 9222 3290 9274
rect 3290 9222 3302 9274
rect 3302 9222 3332 9274
rect 3356 9222 3366 9274
rect 3366 9222 3412 9274
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3276 9220 3332 9222
rect 3356 9220 3412 9222
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 3276 8186 3332 8188
rect 3356 8186 3412 8188
rect 3116 8134 3162 8186
rect 3162 8134 3172 8186
rect 3196 8134 3226 8186
rect 3226 8134 3238 8186
rect 3238 8134 3252 8186
rect 3276 8134 3290 8186
rect 3290 8134 3302 8186
rect 3302 8134 3332 8186
rect 3356 8134 3366 8186
rect 3366 8134 3412 8186
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 3276 8132 3332 8134
rect 3356 8132 3412 8134
rect 4666 10906 4722 10908
rect 4746 10906 4802 10908
rect 4826 10906 4882 10908
rect 4906 10906 4962 10908
rect 4666 10854 4712 10906
rect 4712 10854 4722 10906
rect 4746 10854 4776 10906
rect 4776 10854 4788 10906
rect 4788 10854 4802 10906
rect 4826 10854 4840 10906
rect 4840 10854 4852 10906
rect 4852 10854 4882 10906
rect 4906 10854 4916 10906
rect 4916 10854 4962 10906
rect 4666 10852 4722 10854
rect 4746 10852 4802 10854
rect 4826 10852 4882 10854
rect 4906 10852 4962 10854
rect 7766 10906 7822 10908
rect 7846 10906 7902 10908
rect 7926 10906 7982 10908
rect 8006 10906 8062 10908
rect 7766 10854 7812 10906
rect 7812 10854 7822 10906
rect 7846 10854 7876 10906
rect 7876 10854 7888 10906
rect 7888 10854 7902 10906
rect 7926 10854 7940 10906
rect 7940 10854 7952 10906
rect 7952 10854 7982 10906
rect 8006 10854 8016 10906
rect 8016 10854 8062 10906
rect 7766 10852 7822 10854
rect 7846 10852 7902 10854
rect 7926 10852 7982 10854
rect 8006 10852 8062 10854
rect 10866 10906 10922 10908
rect 10946 10906 11002 10908
rect 11026 10906 11082 10908
rect 11106 10906 11162 10908
rect 10866 10854 10912 10906
rect 10912 10854 10922 10906
rect 10946 10854 10976 10906
rect 10976 10854 10988 10906
rect 10988 10854 11002 10906
rect 11026 10854 11040 10906
rect 11040 10854 11052 10906
rect 11052 10854 11082 10906
rect 11106 10854 11116 10906
rect 11116 10854 11162 10906
rect 10866 10852 10922 10854
rect 10946 10852 11002 10854
rect 11026 10852 11082 10854
rect 11106 10852 11162 10854
rect 13966 10906 14022 10908
rect 14046 10906 14102 10908
rect 14126 10906 14182 10908
rect 14206 10906 14262 10908
rect 13966 10854 14012 10906
rect 14012 10854 14022 10906
rect 14046 10854 14076 10906
rect 14076 10854 14088 10906
rect 14088 10854 14102 10906
rect 14126 10854 14140 10906
rect 14140 10854 14152 10906
rect 14152 10854 14182 10906
rect 14206 10854 14216 10906
rect 14216 10854 14262 10906
rect 13966 10852 14022 10854
rect 14046 10852 14102 10854
rect 14126 10852 14182 10854
rect 14206 10852 14262 10854
rect 6216 10362 6272 10364
rect 6296 10362 6352 10364
rect 6376 10362 6432 10364
rect 6456 10362 6512 10364
rect 6216 10310 6262 10362
rect 6262 10310 6272 10362
rect 6296 10310 6326 10362
rect 6326 10310 6338 10362
rect 6338 10310 6352 10362
rect 6376 10310 6390 10362
rect 6390 10310 6402 10362
rect 6402 10310 6432 10362
rect 6456 10310 6466 10362
rect 6466 10310 6512 10362
rect 6216 10308 6272 10310
rect 6296 10308 6352 10310
rect 6376 10308 6432 10310
rect 6456 10308 6512 10310
rect 9316 10362 9372 10364
rect 9396 10362 9452 10364
rect 9476 10362 9532 10364
rect 9556 10362 9612 10364
rect 9316 10310 9362 10362
rect 9362 10310 9372 10362
rect 9396 10310 9426 10362
rect 9426 10310 9438 10362
rect 9438 10310 9452 10362
rect 9476 10310 9490 10362
rect 9490 10310 9502 10362
rect 9502 10310 9532 10362
rect 9556 10310 9566 10362
rect 9566 10310 9612 10362
rect 9316 10308 9372 10310
rect 9396 10308 9452 10310
rect 9476 10308 9532 10310
rect 9556 10308 9612 10310
rect 4666 9818 4722 9820
rect 4746 9818 4802 9820
rect 4826 9818 4882 9820
rect 4906 9818 4962 9820
rect 4666 9766 4712 9818
rect 4712 9766 4722 9818
rect 4746 9766 4776 9818
rect 4776 9766 4788 9818
rect 4788 9766 4802 9818
rect 4826 9766 4840 9818
rect 4840 9766 4852 9818
rect 4852 9766 4882 9818
rect 4906 9766 4916 9818
rect 4916 9766 4962 9818
rect 4666 9764 4722 9766
rect 4746 9764 4802 9766
rect 4826 9764 4882 9766
rect 4906 9764 4962 9766
rect 4666 8730 4722 8732
rect 4746 8730 4802 8732
rect 4826 8730 4882 8732
rect 4906 8730 4962 8732
rect 4666 8678 4712 8730
rect 4712 8678 4722 8730
rect 4746 8678 4776 8730
rect 4776 8678 4788 8730
rect 4788 8678 4802 8730
rect 4826 8678 4840 8730
rect 4840 8678 4852 8730
rect 4852 8678 4882 8730
rect 4906 8678 4916 8730
rect 4916 8678 4962 8730
rect 4666 8676 4722 8678
rect 4746 8676 4802 8678
rect 4826 8676 4882 8678
rect 4906 8676 4962 8678
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 3276 7098 3332 7100
rect 3356 7098 3412 7100
rect 3116 7046 3162 7098
rect 3162 7046 3172 7098
rect 3196 7046 3226 7098
rect 3226 7046 3238 7098
rect 3238 7046 3252 7098
rect 3276 7046 3290 7098
rect 3290 7046 3302 7098
rect 3302 7046 3332 7098
rect 3356 7046 3366 7098
rect 3366 7046 3412 7098
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3276 7044 3332 7046
rect 3356 7044 3412 7046
rect 4666 7642 4722 7644
rect 4746 7642 4802 7644
rect 4826 7642 4882 7644
rect 4906 7642 4962 7644
rect 4666 7590 4712 7642
rect 4712 7590 4722 7642
rect 4746 7590 4776 7642
rect 4776 7590 4788 7642
rect 4788 7590 4802 7642
rect 4826 7590 4840 7642
rect 4840 7590 4852 7642
rect 4852 7590 4882 7642
rect 4906 7590 4916 7642
rect 4916 7590 4962 7642
rect 4666 7588 4722 7590
rect 4746 7588 4802 7590
rect 4826 7588 4882 7590
rect 4906 7588 4962 7590
rect 4666 6554 4722 6556
rect 4746 6554 4802 6556
rect 4826 6554 4882 6556
rect 4906 6554 4962 6556
rect 4666 6502 4712 6554
rect 4712 6502 4722 6554
rect 4746 6502 4776 6554
rect 4776 6502 4788 6554
rect 4788 6502 4802 6554
rect 4826 6502 4840 6554
rect 4840 6502 4852 6554
rect 4852 6502 4882 6554
rect 4906 6502 4916 6554
rect 4916 6502 4962 6554
rect 4666 6500 4722 6502
rect 4746 6500 4802 6502
rect 4826 6500 4882 6502
rect 4906 6500 4962 6502
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 3276 6010 3332 6012
rect 3356 6010 3412 6012
rect 3116 5958 3162 6010
rect 3162 5958 3172 6010
rect 3196 5958 3226 6010
rect 3226 5958 3238 6010
rect 3238 5958 3252 6010
rect 3276 5958 3290 6010
rect 3290 5958 3302 6010
rect 3302 5958 3332 6010
rect 3356 5958 3366 6010
rect 3366 5958 3412 6010
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 3276 5956 3332 5958
rect 3356 5956 3412 5958
rect 6216 9274 6272 9276
rect 6296 9274 6352 9276
rect 6376 9274 6432 9276
rect 6456 9274 6512 9276
rect 6216 9222 6262 9274
rect 6262 9222 6272 9274
rect 6296 9222 6326 9274
rect 6326 9222 6338 9274
rect 6338 9222 6352 9274
rect 6376 9222 6390 9274
rect 6390 9222 6402 9274
rect 6402 9222 6432 9274
rect 6456 9222 6466 9274
rect 6466 9222 6512 9274
rect 6216 9220 6272 9222
rect 6296 9220 6352 9222
rect 6376 9220 6432 9222
rect 6456 9220 6512 9222
rect 7766 9818 7822 9820
rect 7846 9818 7902 9820
rect 7926 9818 7982 9820
rect 8006 9818 8062 9820
rect 7766 9766 7812 9818
rect 7812 9766 7822 9818
rect 7846 9766 7876 9818
rect 7876 9766 7888 9818
rect 7888 9766 7902 9818
rect 7926 9766 7940 9818
rect 7940 9766 7952 9818
rect 7952 9766 7982 9818
rect 8006 9766 8016 9818
rect 8016 9766 8062 9818
rect 7766 9764 7822 9766
rect 7846 9764 7902 9766
rect 7926 9764 7982 9766
rect 8006 9764 8062 9766
rect 7766 8730 7822 8732
rect 7846 8730 7902 8732
rect 7926 8730 7982 8732
rect 8006 8730 8062 8732
rect 7766 8678 7812 8730
rect 7812 8678 7822 8730
rect 7846 8678 7876 8730
rect 7876 8678 7888 8730
rect 7888 8678 7902 8730
rect 7926 8678 7940 8730
rect 7940 8678 7952 8730
rect 7952 8678 7982 8730
rect 8006 8678 8016 8730
rect 8016 8678 8062 8730
rect 7766 8676 7822 8678
rect 7846 8676 7902 8678
rect 7926 8676 7982 8678
rect 8006 8676 8062 8678
rect 6216 8186 6272 8188
rect 6296 8186 6352 8188
rect 6376 8186 6432 8188
rect 6456 8186 6512 8188
rect 6216 8134 6262 8186
rect 6262 8134 6272 8186
rect 6296 8134 6326 8186
rect 6326 8134 6338 8186
rect 6338 8134 6352 8186
rect 6376 8134 6390 8186
rect 6390 8134 6402 8186
rect 6402 8134 6432 8186
rect 6456 8134 6466 8186
rect 6466 8134 6512 8186
rect 6216 8132 6272 8134
rect 6296 8132 6352 8134
rect 6376 8132 6432 8134
rect 6456 8132 6512 8134
rect 6216 7098 6272 7100
rect 6296 7098 6352 7100
rect 6376 7098 6432 7100
rect 6456 7098 6512 7100
rect 6216 7046 6262 7098
rect 6262 7046 6272 7098
rect 6296 7046 6326 7098
rect 6326 7046 6338 7098
rect 6338 7046 6352 7098
rect 6376 7046 6390 7098
rect 6390 7046 6402 7098
rect 6402 7046 6432 7098
rect 6456 7046 6466 7098
rect 6466 7046 6512 7098
rect 6216 7044 6272 7046
rect 6296 7044 6352 7046
rect 6376 7044 6432 7046
rect 6456 7044 6512 7046
rect 6216 6010 6272 6012
rect 6296 6010 6352 6012
rect 6376 6010 6432 6012
rect 6456 6010 6512 6012
rect 6216 5958 6262 6010
rect 6262 5958 6272 6010
rect 6296 5958 6326 6010
rect 6326 5958 6338 6010
rect 6338 5958 6352 6010
rect 6376 5958 6390 6010
rect 6390 5958 6402 6010
rect 6402 5958 6432 6010
rect 6456 5958 6466 6010
rect 6466 5958 6512 6010
rect 6216 5956 6272 5958
rect 6296 5956 6352 5958
rect 6376 5956 6432 5958
rect 6456 5956 6512 5958
rect 9316 9274 9372 9276
rect 9396 9274 9452 9276
rect 9476 9274 9532 9276
rect 9556 9274 9612 9276
rect 9316 9222 9362 9274
rect 9362 9222 9372 9274
rect 9396 9222 9426 9274
rect 9426 9222 9438 9274
rect 9438 9222 9452 9274
rect 9476 9222 9490 9274
rect 9490 9222 9502 9274
rect 9502 9222 9532 9274
rect 9556 9222 9566 9274
rect 9566 9222 9612 9274
rect 9316 9220 9372 9222
rect 9396 9220 9452 9222
rect 9476 9220 9532 9222
rect 9556 9220 9612 9222
rect 4666 5466 4722 5468
rect 4746 5466 4802 5468
rect 4826 5466 4882 5468
rect 4906 5466 4962 5468
rect 4666 5414 4712 5466
rect 4712 5414 4722 5466
rect 4746 5414 4776 5466
rect 4776 5414 4788 5466
rect 4788 5414 4802 5466
rect 4826 5414 4840 5466
rect 4840 5414 4852 5466
rect 4852 5414 4882 5466
rect 4906 5414 4916 5466
rect 4916 5414 4962 5466
rect 4666 5412 4722 5414
rect 4746 5412 4802 5414
rect 4826 5412 4882 5414
rect 4906 5412 4962 5414
rect 7766 7642 7822 7644
rect 7846 7642 7902 7644
rect 7926 7642 7982 7644
rect 8006 7642 8062 7644
rect 7766 7590 7812 7642
rect 7812 7590 7822 7642
rect 7846 7590 7876 7642
rect 7876 7590 7888 7642
rect 7888 7590 7902 7642
rect 7926 7590 7940 7642
rect 7940 7590 7952 7642
rect 7952 7590 7982 7642
rect 8006 7590 8016 7642
rect 8016 7590 8062 7642
rect 7766 7588 7822 7590
rect 7846 7588 7902 7590
rect 7926 7588 7982 7590
rect 8006 7588 8062 7590
rect 7766 6554 7822 6556
rect 7846 6554 7902 6556
rect 7926 6554 7982 6556
rect 8006 6554 8062 6556
rect 7766 6502 7812 6554
rect 7812 6502 7822 6554
rect 7846 6502 7876 6554
rect 7876 6502 7888 6554
rect 7888 6502 7902 6554
rect 7926 6502 7940 6554
rect 7940 6502 7952 6554
rect 7952 6502 7982 6554
rect 8006 6502 8016 6554
rect 8016 6502 8062 6554
rect 7766 6500 7822 6502
rect 7846 6500 7902 6502
rect 7926 6500 7982 6502
rect 8006 6500 8062 6502
rect 10866 9818 10922 9820
rect 10946 9818 11002 9820
rect 11026 9818 11082 9820
rect 11106 9818 11162 9820
rect 10866 9766 10912 9818
rect 10912 9766 10922 9818
rect 10946 9766 10976 9818
rect 10976 9766 10988 9818
rect 10988 9766 11002 9818
rect 11026 9766 11040 9818
rect 11040 9766 11052 9818
rect 11052 9766 11082 9818
rect 11106 9766 11116 9818
rect 11116 9766 11162 9818
rect 10866 9764 10922 9766
rect 10946 9764 11002 9766
rect 11026 9764 11082 9766
rect 11106 9764 11162 9766
rect 9316 8186 9372 8188
rect 9396 8186 9452 8188
rect 9476 8186 9532 8188
rect 9556 8186 9612 8188
rect 9316 8134 9362 8186
rect 9362 8134 9372 8186
rect 9396 8134 9426 8186
rect 9426 8134 9438 8186
rect 9438 8134 9452 8186
rect 9476 8134 9490 8186
rect 9490 8134 9502 8186
rect 9502 8134 9532 8186
rect 9556 8134 9566 8186
rect 9566 8134 9612 8186
rect 9316 8132 9372 8134
rect 9396 8132 9452 8134
rect 9476 8132 9532 8134
rect 9556 8132 9612 8134
rect 7766 5466 7822 5468
rect 7846 5466 7902 5468
rect 7926 5466 7982 5468
rect 8006 5466 8062 5468
rect 7766 5414 7812 5466
rect 7812 5414 7822 5466
rect 7846 5414 7876 5466
rect 7876 5414 7888 5466
rect 7888 5414 7902 5466
rect 7926 5414 7940 5466
rect 7940 5414 7952 5466
rect 7952 5414 7982 5466
rect 8006 5414 8016 5466
rect 8016 5414 8062 5466
rect 7766 5412 7822 5414
rect 7846 5412 7902 5414
rect 7926 5412 7982 5414
rect 8006 5412 8062 5414
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 3276 4922 3332 4924
rect 3356 4922 3412 4924
rect 3116 4870 3162 4922
rect 3162 4870 3172 4922
rect 3196 4870 3226 4922
rect 3226 4870 3238 4922
rect 3238 4870 3252 4922
rect 3276 4870 3290 4922
rect 3290 4870 3302 4922
rect 3302 4870 3332 4922
rect 3356 4870 3366 4922
rect 3366 4870 3412 4922
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 3276 4868 3332 4870
rect 3356 4868 3412 4870
rect 6216 4922 6272 4924
rect 6296 4922 6352 4924
rect 6376 4922 6432 4924
rect 6456 4922 6512 4924
rect 6216 4870 6262 4922
rect 6262 4870 6272 4922
rect 6296 4870 6326 4922
rect 6326 4870 6338 4922
rect 6338 4870 6352 4922
rect 6376 4870 6390 4922
rect 6390 4870 6402 4922
rect 6402 4870 6432 4922
rect 6456 4870 6466 4922
rect 6466 4870 6512 4922
rect 6216 4868 6272 4870
rect 6296 4868 6352 4870
rect 6376 4868 6432 4870
rect 6456 4868 6512 4870
rect 4666 4378 4722 4380
rect 4746 4378 4802 4380
rect 4826 4378 4882 4380
rect 4906 4378 4962 4380
rect 4666 4326 4712 4378
rect 4712 4326 4722 4378
rect 4746 4326 4776 4378
rect 4776 4326 4788 4378
rect 4788 4326 4802 4378
rect 4826 4326 4840 4378
rect 4840 4326 4852 4378
rect 4852 4326 4882 4378
rect 4906 4326 4916 4378
rect 4916 4326 4962 4378
rect 4666 4324 4722 4326
rect 4746 4324 4802 4326
rect 4826 4324 4882 4326
rect 4906 4324 4962 4326
rect 3054 4140 3110 4176
rect 3054 4120 3056 4140
rect 3056 4120 3108 4140
rect 3108 4120 3110 4140
rect 3514 4120 3570 4176
rect 4986 4140 5042 4176
rect 4986 4120 4988 4140
rect 4988 4120 5040 4140
rect 5040 4120 5042 4140
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 3276 3834 3332 3836
rect 3356 3834 3412 3836
rect 3116 3782 3162 3834
rect 3162 3782 3172 3834
rect 3196 3782 3226 3834
rect 3226 3782 3238 3834
rect 3238 3782 3252 3834
rect 3276 3782 3290 3834
rect 3290 3782 3302 3834
rect 3302 3782 3332 3834
rect 3356 3782 3366 3834
rect 3366 3782 3412 3834
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 3276 3780 3332 3782
rect 3356 3780 3412 3782
rect 7766 4378 7822 4380
rect 7846 4378 7902 4380
rect 7926 4378 7982 4380
rect 8006 4378 8062 4380
rect 7766 4326 7812 4378
rect 7812 4326 7822 4378
rect 7846 4326 7876 4378
rect 7876 4326 7888 4378
rect 7888 4326 7902 4378
rect 7926 4326 7940 4378
rect 7940 4326 7952 4378
rect 7952 4326 7982 4378
rect 8006 4326 8016 4378
rect 8016 4326 8062 4378
rect 7766 4324 7822 4326
rect 7846 4324 7902 4326
rect 7926 4324 7982 4326
rect 8006 4324 8062 4326
rect 6216 3834 6272 3836
rect 6296 3834 6352 3836
rect 6376 3834 6432 3836
rect 6456 3834 6512 3836
rect 6216 3782 6262 3834
rect 6262 3782 6272 3834
rect 6296 3782 6326 3834
rect 6326 3782 6338 3834
rect 6338 3782 6352 3834
rect 6376 3782 6390 3834
rect 6390 3782 6402 3834
rect 6402 3782 6432 3834
rect 6456 3782 6466 3834
rect 6466 3782 6512 3834
rect 6216 3780 6272 3782
rect 6296 3780 6352 3782
rect 6376 3780 6432 3782
rect 6456 3780 6512 3782
rect 4666 3290 4722 3292
rect 4746 3290 4802 3292
rect 4826 3290 4882 3292
rect 4906 3290 4962 3292
rect 4666 3238 4712 3290
rect 4712 3238 4722 3290
rect 4746 3238 4776 3290
rect 4776 3238 4788 3290
rect 4788 3238 4802 3290
rect 4826 3238 4840 3290
rect 4840 3238 4852 3290
rect 4852 3238 4882 3290
rect 4906 3238 4916 3290
rect 4916 3238 4962 3290
rect 4666 3236 4722 3238
rect 4746 3236 4802 3238
rect 4826 3236 4882 3238
rect 4906 3236 4962 3238
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 3276 2746 3332 2748
rect 3356 2746 3412 2748
rect 3116 2694 3162 2746
rect 3162 2694 3172 2746
rect 3196 2694 3226 2746
rect 3226 2694 3238 2746
rect 3238 2694 3252 2746
rect 3276 2694 3290 2746
rect 3290 2694 3302 2746
rect 3302 2694 3332 2746
rect 3356 2694 3366 2746
rect 3366 2694 3412 2746
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 3276 2692 3332 2694
rect 3356 2692 3412 2694
rect 4666 2202 4722 2204
rect 4746 2202 4802 2204
rect 4826 2202 4882 2204
rect 4906 2202 4962 2204
rect 4666 2150 4712 2202
rect 4712 2150 4722 2202
rect 4746 2150 4776 2202
rect 4776 2150 4788 2202
rect 4788 2150 4802 2202
rect 4826 2150 4840 2202
rect 4840 2150 4852 2202
rect 4852 2150 4882 2202
rect 4906 2150 4916 2202
rect 4916 2150 4962 2202
rect 4666 2148 4722 2150
rect 4746 2148 4802 2150
rect 4826 2148 4882 2150
rect 4906 2148 4962 2150
rect 3116 1658 3172 1660
rect 3196 1658 3252 1660
rect 3276 1658 3332 1660
rect 3356 1658 3412 1660
rect 3116 1606 3162 1658
rect 3162 1606 3172 1658
rect 3196 1606 3226 1658
rect 3226 1606 3238 1658
rect 3238 1606 3252 1658
rect 3276 1606 3290 1658
rect 3290 1606 3302 1658
rect 3302 1606 3332 1658
rect 3356 1606 3366 1658
rect 3366 1606 3412 1658
rect 3116 1604 3172 1606
rect 3196 1604 3252 1606
rect 3276 1604 3332 1606
rect 3356 1604 3412 1606
rect 3606 1264 3662 1320
rect 3116 570 3172 572
rect 3196 570 3252 572
rect 3276 570 3332 572
rect 3356 570 3412 572
rect 3116 518 3162 570
rect 3162 518 3172 570
rect 3196 518 3226 570
rect 3226 518 3238 570
rect 3238 518 3252 570
rect 3276 518 3290 570
rect 3290 518 3302 570
rect 3302 518 3332 570
rect 3356 518 3366 570
rect 3366 518 3412 570
rect 3116 516 3172 518
rect 3196 516 3252 518
rect 3276 516 3332 518
rect 3356 516 3412 518
rect 4666 1114 4722 1116
rect 4746 1114 4802 1116
rect 4826 1114 4882 1116
rect 4906 1114 4962 1116
rect 4666 1062 4712 1114
rect 4712 1062 4722 1114
rect 4746 1062 4776 1114
rect 4776 1062 4788 1114
rect 4788 1062 4802 1114
rect 4826 1062 4840 1114
rect 4840 1062 4852 1114
rect 4852 1062 4882 1114
rect 4906 1062 4916 1114
rect 4916 1062 4962 1114
rect 4666 1060 4722 1062
rect 4746 1060 4802 1062
rect 4826 1060 4882 1062
rect 4906 1060 4962 1062
rect 6216 2746 6272 2748
rect 6296 2746 6352 2748
rect 6376 2746 6432 2748
rect 6456 2746 6512 2748
rect 6216 2694 6262 2746
rect 6262 2694 6272 2746
rect 6296 2694 6326 2746
rect 6326 2694 6338 2746
rect 6338 2694 6352 2746
rect 6376 2694 6390 2746
rect 6390 2694 6402 2746
rect 6402 2694 6432 2746
rect 6456 2694 6466 2746
rect 6466 2694 6512 2746
rect 6216 2692 6272 2694
rect 6296 2692 6352 2694
rect 6376 2692 6432 2694
rect 6456 2692 6512 2694
rect 6216 1658 6272 1660
rect 6296 1658 6352 1660
rect 6376 1658 6432 1660
rect 6456 1658 6512 1660
rect 6216 1606 6262 1658
rect 6262 1606 6272 1658
rect 6296 1606 6326 1658
rect 6326 1606 6338 1658
rect 6338 1606 6352 1658
rect 6376 1606 6390 1658
rect 6390 1606 6402 1658
rect 6402 1606 6432 1658
rect 6456 1606 6466 1658
rect 6466 1606 6512 1658
rect 6216 1604 6272 1606
rect 6296 1604 6352 1606
rect 6376 1604 6432 1606
rect 6456 1604 6512 1606
rect 5538 1264 5594 1320
rect 6366 756 6368 776
rect 6368 756 6420 776
rect 6420 756 6422 776
rect 6366 720 6422 756
rect 6642 720 6698 776
rect 7766 3290 7822 3292
rect 7846 3290 7902 3292
rect 7926 3290 7982 3292
rect 8006 3290 8062 3292
rect 7766 3238 7812 3290
rect 7812 3238 7822 3290
rect 7846 3238 7876 3290
rect 7876 3238 7888 3290
rect 7888 3238 7902 3290
rect 7926 3238 7940 3290
rect 7940 3238 7952 3290
rect 7952 3238 7982 3290
rect 8006 3238 8016 3290
rect 8016 3238 8062 3290
rect 7766 3236 7822 3238
rect 7846 3236 7902 3238
rect 7926 3236 7982 3238
rect 8006 3236 8062 3238
rect 12416 10362 12472 10364
rect 12496 10362 12552 10364
rect 12576 10362 12632 10364
rect 12656 10362 12712 10364
rect 12416 10310 12462 10362
rect 12462 10310 12472 10362
rect 12496 10310 12526 10362
rect 12526 10310 12538 10362
rect 12538 10310 12552 10362
rect 12576 10310 12590 10362
rect 12590 10310 12602 10362
rect 12602 10310 12632 10362
rect 12656 10310 12666 10362
rect 12666 10310 12712 10362
rect 12416 10308 12472 10310
rect 12496 10308 12552 10310
rect 12576 10308 12632 10310
rect 12656 10308 12712 10310
rect 10866 8730 10922 8732
rect 10946 8730 11002 8732
rect 11026 8730 11082 8732
rect 11106 8730 11162 8732
rect 10866 8678 10912 8730
rect 10912 8678 10922 8730
rect 10946 8678 10976 8730
rect 10976 8678 10988 8730
rect 10988 8678 11002 8730
rect 11026 8678 11040 8730
rect 11040 8678 11052 8730
rect 11052 8678 11082 8730
rect 11106 8678 11116 8730
rect 11116 8678 11162 8730
rect 10866 8676 10922 8678
rect 10946 8676 11002 8678
rect 11026 8676 11082 8678
rect 11106 8676 11162 8678
rect 9316 7098 9372 7100
rect 9396 7098 9452 7100
rect 9476 7098 9532 7100
rect 9556 7098 9612 7100
rect 9316 7046 9362 7098
rect 9362 7046 9372 7098
rect 9396 7046 9426 7098
rect 9426 7046 9438 7098
rect 9438 7046 9452 7098
rect 9476 7046 9490 7098
rect 9490 7046 9502 7098
rect 9502 7046 9532 7098
rect 9556 7046 9566 7098
rect 9566 7046 9612 7098
rect 9316 7044 9372 7046
rect 9396 7044 9452 7046
rect 9476 7044 9532 7046
rect 9556 7044 9612 7046
rect 13966 9818 14022 9820
rect 14046 9818 14102 9820
rect 14126 9818 14182 9820
rect 14206 9818 14262 9820
rect 13966 9766 14012 9818
rect 14012 9766 14022 9818
rect 14046 9766 14076 9818
rect 14076 9766 14088 9818
rect 14088 9766 14102 9818
rect 14126 9766 14140 9818
rect 14140 9766 14152 9818
rect 14152 9766 14182 9818
rect 14206 9766 14216 9818
rect 14216 9766 14262 9818
rect 13966 9764 14022 9766
rect 14046 9764 14102 9766
rect 14126 9764 14182 9766
rect 14206 9764 14262 9766
rect 12416 9274 12472 9276
rect 12496 9274 12552 9276
rect 12576 9274 12632 9276
rect 12656 9274 12712 9276
rect 12416 9222 12462 9274
rect 12462 9222 12472 9274
rect 12496 9222 12526 9274
rect 12526 9222 12538 9274
rect 12538 9222 12552 9274
rect 12576 9222 12590 9274
rect 12590 9222 12602 9274
rect 12602 9222 12632 9274
rect 12656 9222 12666 9274
rect 12666 9222 12712 9274
rect 12416 9220 12472 9222
rect 12496 9220 12552 9222
rect 12576 9220 12632 9222
rect 12656 9220 12712 9222
rect 10866 7642 10922 7644
rect 10946 7642 11002 7644
rect 11026 7642 11082 7644
rect 11106 7642 11162 7644
rect 10866 7590 10912 7642
rect 10912 7590 10922 7642
rect 10946 7590 10976 7642
rect 10976 7590 10988 7642
rect 10988 7590 11002 7642
rect 11026 7590 11040 7642
rect 11040 7590 11052 7642
rect 11052 7590 11082 7642
rect 11106 7590 11116 7642
rect 11116 7590 11162 7642
rect 10866 7588 10922 7590
rect 10946 7588 11002 7590
rect 11026 7588 11082 7590
rect 11106 7588 11162 7590
rect 9316 6010 9372 6012
rect 9396 6010 9452 6012
rect 9476 6010 9532 6012
rect 9556 6010 9612 6012
rect 9316 5958 9362 6010
rect 9362 5958 9372 6010
rect 9396 5958 9426 6010
rect 9426 5958 9438 6010
rect 9438 5958 9452 6010
rect 9476 5958 9490 6010
rect 9490 5958 9502 6010
rect 9502 5958 9532 6010
rect 9556 5958 9566 6010
rect 9566 5958 9612 6010
rect 9316 5956 9372 5958
rect 9396 5956 9452 5958
rect 9476 5956 9532 5958
rect 9556 5956 9612 5958
rect 10866 6554 10922 6556
rect 10946 6554 11002 6556
rect 11026 6554 11082 6556
rect 11106 6554 11162 6556
rect 10866 6502 10912 6554
rect 10912 6502 10922 6554
rect 10946 6502 10976 6554
rect 10976 6502 10988 6554
rect 10988 6502 11002 6554
rect 11026 6502 11040 6554
rect 11040 6502 11052 6554
rect 11052 6502 11082 6554
rect 11106 6502 11116 6554
rect 11116 6502 11162 6554
rect 10866 6500 10922 6502
rect 10946 6500 11002 6502
rect 11026 6500 11082 6502
rect 11106 6500 11162 6502
rect 12416 8186 12472 8188
rect 12496 8186 12552 8188
rect 12576 8186 12632 8188
rect 12656 8186 12712 8188
rect 12416 8134 12462 8186
rect 12462 8134 12472 8186
rect 12496 8134 12526 8186
rect 12526 8134 12538 8186
rect 12538 8134 12552 8186
rect 12576 8134 12590 8186
rect 12590 8134 12602 8186
rect 12602 8134 12632 8186
rect 12656 8134 12666 8186
rect 12666 8134 12712 8186
rect 12416 8132 12472 8134
rect 12496 8132 12552 8134
rect 12576 8132 12632 8134
rect 12656 8132 12712 8134
rect 13966 8730 14022 8732
rect 14046 8730 14102 8732
rect 14126 8730 14182 8732
rect 14206 8730 14262 8732
rect 13966 8678 14012 8730
rect 14012 8678 14022 8730
rect 14046 8678 14076 8730
rect 14076 8678 14088 8730
rect 14088 8678 14102 8730
rect 14126 8678 14140 8730
rect 14140 8678 14152 8730
rect 14152 8678 14182 8730
rect 14206 8678 14216 8730
rect 14216 8678 14262 8730
rect 13966 8676 14022 8678
rect 14046 8676 14102 8678
rect 14126 8676 14182 8678
rect 14206 8676 14262 8678
rect 13450 7404 13506 7440
rect 13450 7384 13452 7404
rect 13452 7384 13504 7404
rect 13504 7384 13506 7404
rect 13966 7642 14022 7644
rect 14046 7642 14102 7644
rect 14126 7642 14182 7644
rect 14206 7642 14262 7644
rect 13966 7590 14012 7642
rect 14012 7590 14022 7642
rect 14046 7590 14076 7642
rect 14076 7590 14088 7642
rect 14088 7590 14102 7642
rect 14126 7590 14140 7642
rect 14140 7590 14152 7642
rect 14152 7590 14182 7642
rect 14206 7590 14216 7642
rect 14216 7590 14262 7642
rect 13966 7588 14022 7590
rect 14046 7588 14102 7590
rect 14126 7588 14182 7590
rect 14206 7588 14262 7590
rect 12416 7098 12472 7100
rect 12496 7098 12552 7100
rect 12576 7098 12632 7100
rect 12656 7098 12712 7100
rect 12416 7046 12462 7098
rect 12462 7046 12472 7098
rect 12496 7046 12526 7098
rect 12526 7046 12538 7098
rect 12538 7046 12552 7098
rect 12576 7046 12590 7098
rect 12590 7046 12602 7098
rect 12602 7046 12632 7098
rect 12656 7046 12666 7098
rect 12666 7046 12712 7098
rect 12416 7044 12472 7046
rect 12496 7044 12552 7046
rect 12576 7044 12632 7046
rect 12656 7044 12712 7046
rect 11610 6740 11612 6760
rect 11612 6740 11664 6760
rect 11664 6740 11666 6760
rect 11610 6704 11666 6740
rect 12416 6010 12472 6012
rect 12496 6010 12552 6012
rect 12576 6010 12632 6012
rect 12656 6010 12712 6012
rect 12416 5958 12462 6010
rect 12462 5958 12472 6010
rect 12496 5958 12526 6010
rect 12526 5958 12538 6010
rect 12538 5958 12552 6010
rect 12576 5958 12590 6010
rect 12590 5958 12602 6010
rect 12602 5958 12632 6010
rect 12656 5958 12666 6010
rect 12666 5958 12712 6010
rect 12416 5956 12472 5958
rect 12496 5956 12552 5958
rect 12576 5956 12632 5958
rect 12656 5956 12712 5958
rect 10866 5466 10922 5468
rect 10946 5466 11002 5468
rect 11026 5466 11082 5468
rect 11106 5466 11162 5468
rect 10866 5414 10912 5466
rect 10912 5414 10922 5466
rect 10946 5414 10976 5466
rect 10976 5414 10988 5466
rect 10988 5414 11002 5466
rect 11026 5414 11040 5466
rect 11040 5414 11052 5466
rect 11052 5414 11082 5466
rect 11106 5414 11116 5466
rect 11116 5414 11162 5466
rect 10866 5412 10922 5414
rect 10946 5412 11002 5414
rect 11026 5412 11082 5414
rect 11106 5412 11162 5414
rect 9316 4922 9372 4924
rect 9396 4922 9452 4924
rect 9476 4922 9532 4924
rect 9556 4922 9612 4924
rect 9316 4870 9362 4922
rect 9362 4870 9372 4922
rect 9396 4870 9426 4922
rect 9426 4870 9438 4922
rect 9438 4870 9452 4922
rect 9476 4870 9490 4922
rect 9490 4870 9502 4922
rect 9502 4870 9532 4922
rect 9556 4870 9566 4922
rect 9566 4870 9612 4922
rect 9316 4868 9372 4870
rect 9396 4868 9452 4870
rect 9476 4868 9532 4870
rect 9556 4868 9612 4870
rect 13266 7268 13322 7304
rect 13266 7248 13268 7268
rect 13268 7248 13320 7268
rect 13320 7248 13322 7268
rect 14554 7420 14556 7440
rect 14556 7420 14608 7440
rect 14608 7420 14610 7440
rect 14554 7384 14610 7420
rect 13726 5772 13782 5808
rect 13726 5752 13728 5772
rect 13728 5752 13780 5772
rect 13780 5752 13782 5772
rect 13966 6554 14022 6556
rect 14046 6554 14102 6556
rect 14126 6554 14182 6556
rect 14206 6554 14262 6556
rect 13966 6502 14012 6554
rect 14012 6502 14022 6554
rect 14046 6502 14076 6554
rect 14076 6502 14088 6554
rect 14088 6502 14102 6554
rect 14126 6502 14140 6554
rect 14140 6502 14152 6554
rect 14152 6502 14182 6554
rect 14206 6502 14216 6554
rect 14216 6502 14262 6554
rect 13966 6500 14022 6502
rect 14046 6500 14102 6502
rect 14126 6500 14182 6502
rect 14206 6500 14262 6502
rect 14738 7284 14740 7304
rect 14740 7284 14792 7304
rect 14792 7284 14794 7304
rect 14738 7248 14794 7284
rect 13966 5466 14022 5468
rect 14046 5466 14102 5468
rect 14126 5466 14182 5468
rect 14206 5466 14262 5468
rect 13966 5414 14012 5466
rect 14012 5414 14022 5466
rect 14046 5414 14076 5466
rect 14076 5414 14088 5466
rect 14088 5414 14102 5466
rect 14126 5414 14140 5466
rect 14140 5414 14152 5466
rect 14152 5414 14182 5466
rect 14206 5414 14216 5466
rect 14216 5414 14262 5466
rect 13966 5412 14022 5414
rect 14046 5412 14102 5414
rect 14126 5412 14182 5414
rect 14206 5412 14262 5414
rect 9316 3834 9372 3836
rect 9396 3834 9452 3836
rect 9476 3834 9532 3836
rect 9556 3834 9612 3836
rect 9316 3782 9362 3834
rect 9362 3782 9372 3834
rect 9396 3782 9426 3834
rect 9426 3782 9438 3834
rect 9438 3782 9452 3834
rect 9476 3782 9490 3834
rect 9490 3782 9502 3834
rect 9502 3782 9532 3834
rect 9556 3782 9566 3834
rect 9566 3782 9612 3834
rect 9316 3780 9372 3782
rect 9396 3780 9452 3782
rect 9476 3780 9532 3782
rect 9556 3780 9612 3782
rect 10866 4378 10922 4380
rect 10946 4378 11002 4380
rect 11026 4378 11082 4380
rect 11106 4378 11162 4380
rect 10866 4326 10912 4378
rect 10912 4326 10922 4378
rect 10946 4326 10976 4378
rect 10976 4326 10988 4378
rect 10988 4326 11002 4378
rect 11026 4326 11040 4378
rect 11040 4326 11052 4378
rect 11052 4326 11082 4378
rect 11106 4326 11116 4378
rect 11116 4326 11162 4378
rect 10866 4324 10922 4326
rect 10946 4324 11002 4326
rect 11026 4324 11082 4326
rect 11106 4324 11162 4326
rect 12416 4922 12472 4924
rect 12496 4922 12552 4924
rect 12576 4922 12632 4924
rect 12656 4922 12712 4924
rect 12416 4870 12462 4922
rect 12462 4870 12472 4922
rect 12496 4870 12526 4922
rect 12526 4870 12538 4922
rect 12538 4870 12552 4922
rect 12576 4870 12590 4922
rect 12590 4870 12602 4922
rect 12602 4870 12632 4922
rect 12656 4870 12666 4922
rect 12666 4870 12712 4922
rect 12416 4868 12472 4870
rect 12496 4868 12552 4870
rect 12576 4868 12632 4870
rect 12656 4868 12712 4870
rect 7654 2352 7710 2408
rect 9316 2746 9372 2748
rect 9396 2746 9452 2748
rect 9476 2746 9532 2748
rect 9556 2746 9612 2748
rect 9316 2694 9362 2746
rect 9362 2694 9372 2746
rect 9396 2694 9426 2746
rect 9426 2694 9438 2746
rect 9438 2694 9452 2746
rect 9476 2694 9490 2746
rect 9490 2694 9502 2746
rect 9502 2694 9532 2746
rect 9556 2694 9566 2746
rect 9566 2694 9612 2746
rect 9316 2692 9372 2694
rect 9396 2692 9452 2694
rect 9476 2692 9532 2694
rect 9556 2692 9612 2694
rect 7766 2202 7822 2204
rect 7846 2202 7902 2204
rect 7926 2202 7982 2204
rect 8006 2202 8062 2204
rect 7766 2150 7812 2202
rect 7812 2150 7822 2202
rect 7846 2150 7876 2202
rect 7876 2150 7888 2202
rect 7888 2150 7902 2202
rect 7926 2150 7940 2202
rect 7940 2150 7952 2202
rect 7952 2150 7982 2202
rect 8006 2150 8016 2202
rect 8016 2150 8062 2202
rect 7766 2148 7822 2150
rect 7846 2148 7902 2150
rect 7926 2148 7982 2150
rect 8006 2148 8062 2150
rect 9034 2352 9090 2408
rect 9218 2372 9274 2408
rect 9218 2352 9220 2372
rect 9220 2352 9272 2372
rect 9272 2352 9274 2372
rect 7766 1114 7822 1116
rect 7846 1114 7902 1116
rect 7926 1114 7982 1116
rect 8006 1114 8062 1116
rect 7766 1062 7812 1114
rect 7812 1062 7822 1114
rect 7846 1062 7876 1114
rect 7876 1062 7888 1114
rect 7888 1062 7902 1114
rect 7926 1062 7940 1114
rect 7940 1062 7952 1114
rect 7952 1062 7982 1114
rect 8006 1062 8016 1114
rect 8016 1062 8062 1114
rect 7766 1060 7822 1062
rect 7846 1060 7902 1062
rect 7926 1060 7982 1062
rect 8006 1060 8062 1062
rect 6216 570 6272 572
rect 6296 570 6352 572
rect 6376 570 6432 572
rect 6456 570 6512 572
rect 6216 518 6262 570
rect 6262 518 6272 570
rect 6296 518 6326 570
rect 6326 518 6338 570
rect 6338 518 6352 570
rect 6376 518 6390 570
rect 6390 518 6402 570
rect 6402 518 6432 570
rect 6456 518 6466 570
rect 6466 518 6512 570
rect 6216 516 6272 518
rect 6296 516 6352 518
rect 6376 516 6432 518
rect 6456 516 6512 518
rect 9316 1658 9372 1660
rect 9396 1658 9452 1660
rect 9476 1658 9532 1660
rect 9556 1658 9612 1660
rect 9316 1606 9362 1658
rect 9362 1606 9372 1658
rect 9396 1606 9426 1658
rect 9426 1606 9438 1658
rect 9438 1606 9452 1658
rect 9476 1606 9490 1658
rect 9490 1606 9502 1658
rect 9502 1606 9532 1658
rect 9556 1606 9566 1658
rect 9566 1606 9612 1658
rect 9316 1604 9372 1606
rect 9396 1604 9452 1606
rect 9476 1604 9532 1606
rect 9556 1604 9612 1606
rect 10866 3290 10922 3292
rect 10946 3290 11002 3292
rect 11026 3290 11082 3292
rect 11106 3290 11162 3292
rect 10866 3238 10912 3290
rect 10912 3238 10922 3290
rect 10946 3238 10976 3290
rect 10976 3238 10988 3290
rect 10988 3238 11002 3290
rect 11026 3238 11040 3290
rect 11040 3238 11052 3290
rect 11052 3238 11082 3290
rect 11106 3238 11116 3290
rect 11116 3238 11162 3290
rect 10866 3236 10922 3238
rect 10946 3236 11002 3238
rect 11026 3236 11082 3238
rect 11106 3236 11162 3238
rect 10866 2202 10922 2204
rect 10946 2202 11002 2204
rect 11026 2202 11082 2204
rect 11106 2202 11162 2204
rect 10866 2150 10912 2202
rect 10912 2150 10922 2202
rect 10946 2150 10976 2202
rect 10976 2150 10988 2202
rect 10988 2150 11002 2202
rect 11026 2150 11040 2202
rect 11040 2150 11052 2202
rect 11052 2150 11082 2202
rect 11106 2150 11116 2202
rect 11116 2150 11162 2202
rect 10866 2148 10922 2150
rect 10946 2148 11002 2150
rect 11026 2148 11082 2150
rect 11106 2148 11162 2150
rect 9316 570 9372 572
rect 9396 570 9452 572
rect 9476 570 9532 572
rect 9556 570 9612 572
rect 9316 518 9362 570
rect 9362 518 9372 570
rect 9396 518 9426 570
rect 9426 518 9438 570
rect 9438 518 9452 570
rect 9476 518 9490 570
rect 9490 518 9502 570
rect 9502 518 9532 570
rect 9556 518 9566 570
rect 9566 518 9612 570
rect 9316 516 9372 518
rect 9396 516 9452 518
rect 9476 516 9532 518
rect 9556 516 9612 518
rect 10866 1114 10922 1116
rect 10946 1114 11002 1116
rect 11026 1114 11082 1116
rect 11106 1114 11162 1116
rect 10866 1062 10912 1114
rect 10912 1062 10922 1114
rect 10946 1062 10976 1114
rect 10976 1062 10988 1114
rect 10988 1062 11002 1114
rect 11026 1062 11040 1114
rect 11040 1062 11052 1114
rect 11052 1062 11082 1114
rect 11106 1062 11116 1114
rect 11116 1062 11162 1114
rect 10866 1060 10922 1062
rect 10946 1060 11002 1062
rect 11026 1060 11082 1062
rect 11106 1060 11162 1062
rect 11794 892 11796 912
rect 11796 892 11848 912
rect 11848 892 11850 912
rect 11794 856 11850 892
rect 13966 4378 14022 4380
rect 14046 4378 14102 4380
rect 14126 4378 14182 4380
rect 14206 4378 14262 4380
rect 13966 4326 14012 4378
rect 14012 4326 14022 4378
rect 14046 4326 14076 4378
rect 14076 4326 14088 4378
rect 14088 4326 14102 4378
rect 14126 4326 14140 4378
rect 14140 4326 14152 4378
rect 14152 4326 14182 4378
rect 14206 4326 14216 4378
rect 14216 4326 14262 4378
rect 13966 4324 14022 4326
rect 14046 4324 14102 4326
rect 14126 4324 14182 4326
rect 14206 4324 14262 4326
rect 12416 3834 12472 3836
rect 12496 3834 12552 3836
rect 12576 3834 12632 3836
rect 12656 3834 12712 3836
rect 12416 3782 12462 3834
rect 12462 3782 12472 3834
rect 12496 3782 12526 3834
rect 12526 3782 12538 3834
rect 12538 3782 12552 3834
rect 12576 3782 12590 3834
rect 12590 3782 12602 3834
rect 12602 3782 12632 3834
rect 12656 3782 12666 3834
rect 12666 3782 12712 3834
rect 12416 3780 12472 3782
rect 12496 3780 12552 3782
rect 12576 3780 12632 3782
rect 12656 3780 12712 3782
rect 15014 6704 15070 6760
rect 17066 10906 17122 10908
rect 17146 10906 17202 10908
rect 17226 10906 17282 10908
rect 17306 10906 17362 10908
rect 17066 10854 17112 10906
rect 17112 10854 17122 10906
rect 17146 10854 17176 10906
rect 17176 10854 17188 10906
rect 17188 10854 17202 10906
rect 17226 10854 17240 10906
rect 17240 10854 17252 10906
rect 17252 10854 17282 10906
rect 17306 10854 17316 10906
rect 17316 10854 17362 10906
rect 17066 10852 17122 10854
rect 17146 10852 17202 10854
rect 17226 10852 17282 10854
rect 17306 10852 17362 10854
rect 15516 10362 15572 10364
rect 15596 10362 15652 10364
rect 15676 10362 15732 10364
rect 15756 10362 15812 10364
rect 15516 10310 15562 10362
rect 15562 10310 15572 10362
rect 15596 10310 15626 10362
rect 15626 10310 15638 10362
rect 15638 10310 15652 10362
rect 15676 10310 15690 10362
rect 15690 10310 15702 10362
rect 15702 10310 15732 10362
rect 15756 10310 15766 10362
rect 15766 10310 15812 10362
rect 15516 10308 15572 10310
rect 15596 10308 15652 10310
rect 15676 10308 15732 10310
rect 15756 10308 15812 10310
rect 17066 9818 17122 9820
rect 17146 9818 17202 9820
rect 17226 9818 17282 9820
rect 17306 9818 17362 9820
rect 17066 9766 17112 9818
rect 17112 9766 17122 9818
rect 17146 9766 17176 9818
rect 17176 9766 17188 9818
rect 17188 9766 17202 9818
rect 17226 9766 17240 9818
rect 17240 9766 17252 9818
rect 17252 9766 17282 9818
rect 17306 9766 17316 9818
rect 17316 9766 17362 9818
rect 17066 9764 17122 9766
rect 17146 9764 17202 9766
rect 17226 9764 17282 9766
rect 17306 9764 17362 9766
rect 15516 9274 15572 9276
rect 15596 9274 15652 9276
rect 15676 9274 15732 9276
rect 15756 9274 15812 9276
rect 15516 9222 15562 9274
rect 15562 9222 15572 9274
rect 15596 9222 15626 9274
rect 15626 9222 15638 9274
rect 15638 9222 15652 9274
rect 15676 9222 15690 9274
rect 15690 9222 15702 9274
rect 15702 9222 15732 9274
rect 15756 9222 15766 9274
rect 15766 9222 15812 9274
rect 15516 9220 15572 9222
rect 15596 9220 15652 9222
rect 15676 9220 15732 9222
rect 15756 9220 15812 9222
rect 17066 8730 17122 8732
rect 17146 8730 17202 8732
rect 17226 8730 17282 8732
rect 17306 8730 17362 8732
rect 17066 8678 17112 8730
rect 17112 8678 17122 8730
rect 17146 8678 17176 8730
rect 17176 8678 17188 8730
rect 17188 8678 17202 8730
rect 17226 8678 17240 8730
rect 17240 8678 17252 8730
rect 17252 8678 17282 8730
rect 17306 8678 17316 8730
rect 17316 8678 17362 8730
rect 17066 8676 17122 8678
rect 17146 8676 17202 8678
rect 17226 8676 17282 8678
rect 17306 8676 17362 8678
rect 15516 8186 15572 8188
rect 15596 8186 15652 8188
rect 15676 8186 15732 8188
rect 15756 8186 15812 8188
rect 15516 8134 15562 8186
rect 15562 8134 15572 8186
rect 15596 8134 15626 8186
rect 15626 8134 15638 8186
rect 15638 8134 15652 8186
rect 15676 8134 15690 8186
rect 15690 8134 15702 8186
rect 15702 8134 15732 8186
rect 15756 8134 15766 8186
rect 15766 8134 15812 8186
rect 15516 8132 15572 8134
rect 15596 8132 15652 8134
rect 15676 8132 15732 8134
rect 15756 8132 15812 8134
rect 15516 7098 15572 7100
rect 15596 7098 15652 7100
rect 15676 7098 15732 7100
rect 15756 7098 15812 7100
rect 15516 7046 15562 7098
rect 15562 7046 15572 7098
rect 15596 7046 15626 7098
rect 15626 7046 15638 7098
rect 15638 7046 15652 7098
rect 15676 7046 15690 7098
rect 15690 7046 15702 7098
rect 15702 7046 15732 7098
rect 15756 7046 15766 7098
rect 15766 7046 15812 7098
rect 15516 7044 15572 7046
rect 15596 7044 15652 7046
rect 15676 7044 15732 7046
rect 15756 7044 15812 7046
rect 18786 11192 18842 11248
rect 18602 9696 18658 9752
rect 17066 7642 17122 7644
rect 17146 7642 17202 7644
rect 17226 7642 17282 7644
rect 17306 7642 17362 7644
rect 17066 7590 17112 7642
rect 17112 7590 17122 7642
rect 17146 7590 17176 7642
rect 17176 7590 17188 7642
rect 17188 7590 17202 7642
rect 17226 7590 17240 7642
rect 17240 7590 17252 7642
rect 17252 7590 17282 7642
rect 17306 7590 17316 7642
rect 17316 7590 17362 7642
rect 17066 7588 17122 7590
rect 17146 7588 17202 7590
rect 17226 7588 17282 7590
rect 17306 7588 17362 7590
rect 15516 6010 15572 6012
rect 15596 6010 15652 6012
rect 15676 6010 15732 6012
rect 15756 6010 15812 6012
rect 15516 5958 15562 6010
rect 15562 5958 15572 6010
rect 15596 5958 15626 6010
rect 15626 5958 15638 6010
rect 15638 5958 15652 6010
rect 15676 5958 15690 6010
rect 15690 5958 15702 6010
rect 15702 5958 15732 6010
rect 15756 5958 15766 6010
rect 15766 5958 15812 6010
rect 15516 5956 15572 5958
rect 15596 5956 15652 5958
rect 15676 5956 15732 5958
rect 15756 5956 15812 5958
rect 17066 6554 17122 6556
rect 17146 6554 17202 6556
rect 17226 6554 17282 6556
rect 17306 6554 17362 6556
rect 17066 6502 17112 6554
rect 17112 6502 17122 6554
rect 17146 6502 17176 6554
rect 17176 6502 17188 6554
rect 17188 6502 17202 6554
rect 17226 6502 17240 6554
rect 17240 6502 17252 6554
rect 17252 6502 17282 6554
rect 17306 6502 17316 6554
rect 17316 6502 17362 6554
rect 17066 6500 17122 6502
rect 17146 6500 17202 6502
rect 17226 6500 17282 6502
rect 17306 6500 17362 6502
rect 12416 2746 12472 2748
rect 12496 2746 12552 2748
rect 12576 2746 12632 2748
rect 12656 2746 12712 2748
rect 12416 2694 12462 2746
rect 12462 2694 12472 2746
rect 12496 2694 12526 2746
rect 12526 2694 12538 2746
rect 12538 2694 12552 2746
rect 12576 2694 12590 2746
rect 12590 2694 12602 2746
rect 12602 2694 12632 2746
rect 12656 2694 12666 2746
rect 12666 2694 12712 2746
rect 12416 2692 12472 2694
rect 12496 2692 12552 2694
rect 12576 2692 12632 2694
rect 12656 2692 12712 2694
rect 12416 1658 12472 1660
rect 12496 1658 12552 1660
rect 12576 1658 12632 1660
rect 12656 1658 12712 1660
rect 12416 1606 12462 1658
rect 12462 1606 12472 1658
rect 12496 1606 12526 1658
rect 12526 1606 12538 1658
rect 12538 1606 12552 1658
rect 12576 1606 12590 1658
rect 12590 1606 12602 1658
rect 12602 1606 12632 1658
rect 12656 1606 12666 1658
rect 12666 1606 12712 1658
rect 12416 1604 12472 1606
rect 12496 1604 12552 1606
rect 12576 1604 12632 1606
rect 12656 1604 12712 1606
rect 13966 3290 14022 3292
rect 14046 3290 14102 3292
rect 14126 3290 14182 3292
rect 14206 3290 14262 3292
rect 13966 3238 14012 3290
rect 14012 3238 14022 3290
rect 14046 3238 14076 3290
rect 14076 3238 14088 3290
rect 14088 3238 14102 3290
rect 14126 3238 14140 3290
rect 14140 3238 14152 3290
rect 14152 3238 14182 3290
rect 14206 3238 14216 3290
rect 14216 3238 14262 3290
rect 13966 3236 14022 3238
rect 14046 3236 14102 3238
rect 14126 3236 14182 3238
rect 14206 3236 14262 3238
rect 18602 8200 18658 8256
rect 18510 6740 18512 6760
rect 18512 6740 18564 6760
rect 18564 6740 18566 6760
rect 18510 6704 18566 6740
rect 17406 5752 17462 5808
rect 17066 5466 17122 5468
rect 17146 5466 17202 5468
rect 17226 5466 17282 5468
rect 17306 5466 17362 5468
rect 17066 5414 17112 5466
rect 17112 5414 17122 5466
rect 17146 5414 17176 5466
rect 17176 5414 17188 5466
rect 17188 5414 17202 5466
rect 17226 5414 17240 5466
rect 17240 5414 17252 5466
rect 17252 5414 17282 5466
rect 17306 5414 17316 5466
rect 17316 5414 17362 5466
rect 17066 5412 17122 5414
rect 17146 5412 17202 5414
rect 17226 5412 17282 5414
rect 17306 5412 17362 5414
rect 18510 5208 18566 5264
rect 15516 4922 15572 4924
rect 15596 4922 15652 4924
rect 15676 4922 15732 4924
rect 15756 4922 15812 4924
rect 15516 4870 15562 4922
rect 15562 4870 15572 4922
rect 15596 4870 15626 4922
rect 15626 4870 15638 4922
rect 15638 4870 15652 4922
rect 15676 4870 15690 4922
rect 15690 4870 15702 4922
rect 15702 4870 15732 4922
rect 15756 4870 15766 4922
rect 15766 4870 15812 4922
rect 15516 4868 15572 4870
rect 15596 4868 15652 4870
rect 15676 4868 15732 4870
rect 15756 4868 15812 4870
rect 13966 2202 14022 2204
rect 14046 2202 14102 2204
rect 14126 2202 14182 2204
rect 14206 2202 14262 2204
rect 13966 2150 14012 2202
rect 14012 2150 14022 2202
rect 14046 2150 14076 2202
rect 14076 2150 14088 2202
rect 14088 2150 14102 2202
rect 14126 2150 14140 2202
rect 14140 2150 14152 2202
rect 14152 2150 14182 2202
rect 14206 2150 14216 2202
rect 14216 2150 14262 2202
rect 13966 2148 14022 2150
rect 14046 2148 14102 2150
rect 14126 2148 14182 2150
rect 14206 2148 14262 2150
rect 10966 720 11022 776
rect 13966 1114 14022 1116
rect 14046 1114 14102 1116
rect 14126 1114 14182 1116
rect 14206 1114 14262 1116
rect 13966 1062 14012 1114
rect 14012 1062 14022 1114
rect 14046 1062 14076 1114
rect 14076 1062 14088 1114
rect 14088 1062 14102 1114
rect 14126 1062 14140 1114
rect 14140 1062 14152 1114
rect 14152 1062 14182 1114
rect 14206 1062 14216 1114
rect 14216 1062 14262 1114
rect 13966 1060 14022 1062
rect 14046 1060 14102 1062
rect 14126 1060 14182 1062
rect 14206 1060 14262 1062
rect 13818 856 13874 912
rect 12416 570 12472 572
rect 12496 570 12552 572
rect 12576 570 12632 572
rect 12656 570 12712 572
rect 12416 518 12462 570
rect 12462 518 12472 570
rect 12496 518 12526 570
rect 12526 518 12538 570
rect 12538 518 12552 570
rect 12576 518 12590 570
rect 12590 518 12602 570
rect 12602 518 12632 570
rect 12656 518 12666 570
rect 12666 518 12712 570
rect 12416 516 12472 518
rect 12496 516 12552 518
rect 12576 516 12632 518
rect 12656 516 12712 518
rect 17066 4378 17122 4380
rect 17146 4378 17202 4380
rect 17226 4378 17282 4380
rect 17306 4378 17362 4380
rect 17066 4326 17112 4378
rect 17112 4326 17122 4378
rect 17146 4326 17176 4378
rect 17176 4326 17188 4378
rect 17188 4326 17202 4378
rect 17226 4326 17240 4378
rect 17240 4326 17252 4378
rect 17252 4326 17282 4378
rect 17306 4326 17316 4378
rect 17316 4326 17362 4378
rect 17066 4324 17122 4326
rect 17146 4324 17202 4326
rect 17226 4324 17282 4326
rect 17306 4324 17362 4326
rect 15516 3834 15572 3836
rect 15596 3834 15652 3836
rect 15676 3834 15732 3836
rect 15756 3834 15812 3836
rect 15516 3782 15562 3834
rect 15562 3782 15572 3834
rect 15596 3782 15626 3834
rect 15626 3782 15638 3834
rect 15638 3782 15652 3834
rect 15676 3782 15690 3834
rect 15690 3782 15702 3834
rect 15702 3782 15732 3834
rect 15756 3782 15766 3834
rect 15766 3782 15812 3834
rect 15516 3780 15572 3782
rect 15596 3780 15652 3782
rect 15676 3780 15732 3782
rect 15756 3780 15812 3782
rect 17066 3290 17122 3292
rect 17146 3290 17202 3292
rect 17226 3290 17282 3292
rect 17306 3290 17362 3292
rect 17066 3238 17112 3290
rect 17112 3238 17122 3290
rect 17146 3238 17176 3290
rect 17176 3238 17188 3290
rect 17188 3238 17202 3290
rect 17226 3238 17240 3290
rect 17240 3238 17252 3290
rect 17252 3238 17282 3290
rect 17306 3238 17316 3290
rect 17316 3238 17362 3290
rect 17066 3236 17122 3238
rect 17146 3236 17202 3238
rect 17226 3236 17282 3238
rect 17306 3236 17362 3238
rect 15516 2746 15572 2748
rect 15596 2746 15652 2748
rect 15676 2746 15732 2748
rect 15756 2746 15812 2748
rect 15516 2694 15562 2746
rect 15562 2694 15572 2746
rect 15596 2694 15626 2746
rect 15626 2694 15638 2746
rect 15638 2694 15652 2746
rect 15676 2694 15690 2746
rect 15690 2694 15702 2746
rect 15702 2694 15732 2746
rect 15756 2694 15766 2746
rect 15766 2694 15812 2746
rect 15516 2692 15572 2694
rect 15596 2692 15652 2694
rect 15676 2692 15732 2694
rect 15756 2692 15812 2694
rect 15516 1658 15572 1660
rect 15596 1658 15652 1660
rect 15676 1658 15732 1660
rect 15756 1658 15812 1660
rect 15516 1606 15562 1658
rect 15562 1606 15572 1658
rect 15596 1606 15626 1658
rect 15626 1606 15638 1658
rect 15638 1606 15652 1658
rect 15676 1606 15690 1658
rect 15690 1606 15702 1658
rect 15702 1606 15732 1658
rect 15756 1606 15766 1658
rect 15766 1606 15812 1658
rect 15516 1604 15572 1606
rect 15596 1604 15652 1606
rect 15676 1604 15732 1606
rect 15756 1604 15812 1606
rect 17066 2202 17122 2204
rect 17146 2202 17202 2204
rect 17226 2202 17282 2204
rect 17306 2202 17362 2204
rect 17066 2150 17112 2202
rect 17112 2150 17122 2202
rect 17146 2150 17176 2202
rect 17176 2150 17188 2202
rect 17188 2150 17202 2202
rect 17226 2150 17240 2202
rect 17240 2150 17252 2202
rect 17252 2150 17282 2202
rect 17306 2150 17316 2202
rect 17316 2150 17362 2202
rect 17066 2148 17122 2150
rect 17146 2148 17202 2150
rect 17226 2148 17282 2150
rect 17306 2148 17362 2150
rect 15516 570 15572 572
rect 15596 570 15652 572
rect 15676 570 15732 572
rect 15756 570 15812 572
rect 15516 518 15562 570
rect 15562 518 15572 570
rect 15596 518 15626 570
rect 15626 518 15638 570
rect 15638 518 15652 570
rect 15676 518 15690 570
rect 15690 518 15702 570
rect 15702 518 15732 570
rect 15756 518 15766 570
rect 15766 518 15812 570
rect 15516 516 15572 518
rect 15596 516 15652 518
rect 15676 516 15732 518
rect 15756 516 15812 518
rect 14646 312 14702 368
rect 8666 212 8668 232
rect 8668 212 8720 232
rect 8720 212 8722 232
rect 8666 176 8722 212
rect 17066 1114 17122 1116
rect 17146 1114 17202 1116
rect 17226 1114 17282 1116
rect 17306 1114 17362 1116
rect 17066 1062 17112 1114
rect 17112 1062 17122 1114
rect 17146 1062 17176 1114
rect 17176 1062 17188 1114
rect 17188 1062 17202 1114
rect 17226 1062 17240 1114
rect 17240 1062 17252 1114
rect 17252 1062 17282 1114
rect 17306 1062 17316 1114
rect 17316 1062 17362 1114
rect 17066 1060 17122 1062
rect 17146 1060 17202 1062
rect 17226 1060 17282 1062
rect 17306 1060 17362 1062
rect 18510 3712 18566 3768
rect 18510 2216 18566 2272
rect 18142 720 18198 776
rect 17958 312 18014 368
rect 18510 720 18566 776
rect 12622 176 12678 232
rect 4666 26 4722 28
rect 4746 26 4802 28
rect 4826 26 4882 28
rect 4906 26 4962 28
rect 4666 -26 4712 26
rect 4712 -26 4722 26
rect 4746 -26 4776 26
rect 4776 -26 4788 26
rect 4788 -26 4802 26
rect 4826 -26 4840 26
rect 4840 -26 4852 26
rect 4852 -26 4882 26
rect 4906 -26 4916 26
rect 4916 -26 4962 26
rect 4666 -28 4722 -26
rect 4746 -28 4802 -26
rect 4826 -28 4882 -26
rect 4906 -28 4962 -26
rect 7766 26 7822 28
rect 7846 26 7902 28
rect 7926 26 7982 28
rect 8006 26 8062 28
rect 7766 -26 7812 26
rect 7812 -26 7822 26
rect 7846 -26 7876 26
rect 7876 -26 7888 26
rect 7888 -26 7902 26
rect 7926 -26 7940 26
rect 7940 -26 7952 26
rect 7952 -26 7982 26
rect 8006 -26 8016 26
rect 8016 -26 8062 26
rect 7766 -28 7822 -26
rect 7846 -28 7902 -26
rect 7926 -28 7982 -26
rect 8006 -28 8062 -26
rect 10866 26 10922 28
rect 10946 26 11002 28
rect 11026 26 11082 28
rect 11106 26 11162 28
rect 10866 -26 10912 26
rect 10912 -26 10922 26
rect 10946 -26 10976 26
rect 10976 -26 10988 26
rect 10988 -26 11002 26
rect 11026 -26 11040 26
rect 11040 -26 11052 26
rect 11052 -26 11082 26
rect 11106 -26 11116 26
rect 11116 -26 11162 26
rect 10866 -28 10922 -26
rect 10946 -28 11002 -26
rect 11026 -28 11082 -26
rect 11106 -28 11162 -26
rect 13966 26 14022 28
rect 14046 26 14102 28
rect 14126 26 14182 28
rect 14206 26 14262 28
rect 13966 -26 14012 26
rect 14012 -26 14022 26
rect 14046 -26 14076 26
rect 14076 -26 14088 26
rect 14088 -26 14102 26
rect 14126 -26 14140 26
rect 14140 -26 14152 26
rect 14152 -26 14182 26
rect 14206 -26 14216 26
rect 14216 -26 14262 26
rect 13966 -28 14022 -26
rect 14046 -28 14102 -26
rect 14126 -28 14182 -26
rect 14206 -28 14262 -26
rect 17066 26 17122 28
rect 17146 26 17202 28
rect 17226 26 17282 28
rect 17306 26 17362 28
rect 17066 -26 17112 26
rect 17112 -26 17122 26
rect 17146 -26 17176 26
rect 17176 -26 17188 26
rect 17188 -26 17202 26
rect 17226 -26 17240 26
rect 17240 -26 17252 26
rect 17252 -26 17282 26
rect 17306 -26 17316 26
rect 17316 -26 17362 26
rect 17066 -28 17122 -26
rect 17146 -28 17202 -26
rect 17226 -28 17282 -26
rect 17306 -28 17362 -26
<< metal3 >>
rect 18781 11250 18847 11253
rect 19200 11250 20000 11280
rect 18781 11248 20000 11250
rect 18781 11192 18786 11248
rect 18842 11192 20000 11248
rect 18781 11190 20000 11192
rect 18781 11187 18847 11190
rect 19200 11160 20000 11190
rect 4654 10912 4974 10913
rect 4654 10848 4662 10912
rect 4726 10848 4742 10912
rect 4806 10848 4822 10912
rect 4886 10848 4902 10912
rect 4966 10848 4974 10912
rect 4654 10847 4974 10848
rect 7754 10912 8074 10913
rect 7754 10848 7762 10912
rect 7826 10848 7842 10912
rect 7906 10848 7922 10912
rect 7986 10848 8002 10912
rect 8066 10848 8074 10912
rect 7754 10847 8074 10848
rect 10854 10912 11174 10913
rect 10854 10848 10862 10912
rect 10926 10848 10942 10912
rect 11006 10848 11022 10912
rect 11086 10848 11102 10912
rect 11166 10848 11174 10912
rect 10854 10847 11174 10848
rect 13954 10912 14274 10913
rect 13954 10848 13962 10912
rect 14026 10848 14042 10912
rect 14106 10848 14122 10912
rect 14186 10848 14202 10912
rect 14266 10848 14274 10912
rect 13954 10847 14274 10848
rect 17054 10912 17374 10913
rect 17054 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17222 10912
rect 17286 10848 17302 10912
rect 17366 10848 17374 10912
rect 17054 10847 17374 10848
rect 3104 10368 3424 10369
rect 3104 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3272 10368
rect 3336 10304 3352 10368
rect 3416 10304 3424 10368
rect 3104 10303 3424 10304
rect 6204 10368 6524 10369
rect 6204 10304 6212 10368
rect 6276 10304 6292 10368
rect 6356 10304 6372 10368
rect 6436 10304 6452 10368
rect 6516 10304 6524 10368
rect 6204 10303 6524 10304
rect 9304 10368 9624 10369
rect 9304 10304 9312 10368
rect 9376 10304 9392 10368
rect 9456 10304 9472 10368
rect 9536 10304 9552 10368
rect 9616 10304 9624 10368
rect 9304 10303 9624 10304
rect 12404 10368 12724 10369
rect 12404 10304 12412 10368
rect 12476 10304 12492 10368
rect 12556 10304 12572 10368
rect 12636 10304 12652 10368
rect 12716 10304 12724 10368
rect 12404 10303 12724 10304
rect 15504 10368 15824 10369
rect 15504 10304 15512 10368
rect 15576 10304 15592 10368
rect 15656 10304 15672 10368
rect 15736 10304 15752 10368
rect 15816 10304 15824 10368
rect 15504 10303 15824 10304
rect 3141 10162 3207 10165
rect 3969 10162 4035 10165
rect 3141 10160 4035 10162
rect 3141 10104 3146 10160
rect 3202 10104 3974 10160
rect 4030 10104 4035 10160
rect 3141 10102 4035 10104
rect 3141 10099 3207 10102
rect 3969 10099 4035 10102
rect 3233 10026 3299 10029
rect 3969 10026 4035 10029
rect 3233 10024 4035 10026
rect 3233 9968 3238 10024
rect 3294 9968 3974 10024
rect 4030 9968 4035 10024
rect 3233 9966 4035 9968
rect 3233 9963 3299 9966
rect 3969 9963 4035 9966
rect 4654 9824 4974 9825
rect 4654 9760 4662 9824
rect 4726 9760 4742 9824
rect 4806 9760 4822 9824
rect 4886 9760 4902 9824
rect 4966 9760 4974 9824
rect 4654 9759 4974 9760
rect 7754 9824 8074 9825
rect 7754 9760 7762 9824
rect 7826 9760 7842 9824
rect 7906 9760 7922 9824
rect 7986 9760 8002 9824
rect 8066 9760 8074 9824
rect 7754 9759 8074 9760
rect 10854 9824 11174 9825
rect 10854 9760 10862 9824
rect 10926 9760 10942 9824
rect 11006 9760 11022 9824
rect 11086 9760 11102 9824
rect 11166 9760 11174 9824
rect 10854 9759 11174 9760
rect 13954 9824 14274 9825
rect 13954 9760 13962 9824
rect 14026 9760 14042 9824
rect 14106 9760 14122 9824
rect 14186 9760 14202 9824
rect 14266 9760 14274 9824
rect 13954 9759 14274 9760
rect 17054 9824 17374 9825
rect 17054 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17222 9824
rect 17286 9760 17302 9824
rect 17366 9760 17374 9824
rect 17054 9759 17374 9760
rect 18597 9754 18663 9757
rect 19200 9754 20000 9784
rect 18597 9752 20000 9754
rect 18597 9696 18602 9752
rect 18658 9696 20000 9752
rect 18597 9694 20000 9696
rect 18597 9691 18663 9694
rect 19200 9664 20000 9694
rect 2405 9482 2471 9485
rect 3325 9482 3391 9485
rect 2405 9480 3391 9482
rect 2405 9424 2410 9480
rect 2466 9424 3330 9480
rect 3386 9424 3391 9480
rect 2405 9422 3391 9424
rect 2405 9419 2471 9422
rect 3325 9419 3391 9422
rect 3104 9280 3424 9281
rect 3104 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3272 9280
rect 3336 9216 3352 9280
rect 3416 9216 3424 9280
rect 3104 9215 3424 9216
rect 6204 9280 6524 9281
rect 6204 9216 6212 9280
rect 6276 9216 6292 9280
rect 6356 9216 6372 9280
rect 6436 9216 6452 9280
rect 6516 9216 6524 9280
rect 6204 9215 6524 9216
rect 9304 9280 9624 9281
rect 9304 9216 9312 9280
rect 9376 9216 9392 9280
rect 9456 9216 9472 9280
rect 9536 9216 9552 9280
rect 9616 9216 9624 9280
rect 9304 9215 9624 9216
rect 12404 9280 12724 9281
rect 12404 9216 12412 9280
rect 12476 9216 12492 9280
rect 12556 9216 12572 9280
rect 12636 9216 12652 9280
rect 12716 9216 12724 9280
rect 12404 9215 12724 9216
rect 15504 9280 15824 9281
rect 15504 9216 15512 9280
rect 15576 9216 15592 9280
rect 15656 9216 15672 9280
rect 15736 9216 15752 9280
rect 15816 9216 15824 9280
rect 15504 9215 15824 9216
rect 4654 8736 4974 8737
rect 4654 8672 4662 8736
rect 4726 8672 4742 8736
rect 4806 8672 4822 8736
rect 4886 8672 4902 8736
rect 4966 8672 4974 8736
rect 4654 8671 4974 8672
rect 7754 8736 8074 8737
rect 7754 8672 7762 8736
rect 7826 8672 7842 8736
rect 7906 8672 7922 8736
rect 7986 8672 8002 8736
rect 8066 8672 8074 8736
rect 7754 8671 8074 8672
rect 10854 8736 11174 8737
rect 10854 8672 10862 8736
rect 10926 8672 10942 8736
rect 11006 8672 11022 8736
rect 11086 8672 11102 8736
rect 11166 8672 11174 8736
rect 10854 8671 11174 8672
rect 13954 8736 14274 8737
rect 13954 8672 13962 8736
rect 14026 8672 14042 8736
rect 14106 8672 14122 8736
rect 14186 8672 14202 8736
rect 14266 8672 14274 8736
rect 13954 8671 14274 8672
rect 17054 8736 17374 8737
rect 17054 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17222 8736
rect 17286 8672 17302 8736
rect 17366 8672 17374 8736
rect 17054 8671 17374 8672
rect 18597 8258 18663 8261
rect 19200 8258 20000 8288
rect 18597 8256 20000 8258
rect 18597 8200 18602 8256
rect 18658 8200 20000 8256
rect 18597 8198 20000 8200
rect 18597 8195 18663 8198
rect 3104 8192 3424 8193
rect 3104 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3272 8192
rect 3336 8128 3352 8192
rect 3416 8128 3424 8192
rect 3104 8127 3424 8128
rect 6204 8192 6524 8193
rect 6204 8128 6212 8192
rect 6276 8128 6292 8192
rect 6356 8128 6372 8192
rect 6436 8128 6452 8192
rect 6516 8128 6524 8192
rect 6204 8127 6524 8128
rect 9304 8192 9624 8193
rect 9304 8128 9312 8192
rect 9376 8128 9392 8192
rect 9456 8128 9472 8192
rect 9536 8128 9552 8192
rect 9616 8128 9624 8192
rect 9304 8127 9624 8128
rect 12404 8192 12724 8193
rect 12404 8128 12412 8192
rect 12476 8128 12492 8192
rect 12556 8128 12572 8192
rect 12636 8128 12652 8192
rect 12716 8128 12724 8192
rect 12404 8127 12724 8128
rect 15504 8192 15824 8193
rect 15504 8128 15512 8192
rect 15576 8128 15592 8192
rect 15656 8128 15672 8192
rect 15736 8128 15752 8192
rect 15816 8128 15824 8192
rect 19200 8168 20000 8198
rect 15504 8127 15824 8128
rect 4654 7648 4974 7649
rect 4654 7584 4662 7648
rect 4726 7584 4742 7648
rect 4806 7584 4822 7648
rect 4886 7584 4902 7648
rect 4966 7584 4974 7648
rect 4654 7583 4974 7584
rect 7754 7648 8074 7649
rect 7754 7584 7762 7648
rect 7826 7584 7842 7648
rect 7906 7584 7922 7648
rect 7986 7584 8002 7648
rect 8066 7584 8074 7648
rect 7754 7583 8074 7584
rect 10854 7648 11174 7649
rect 10854 7584 10862 7648
rect 10926 7584 10942 7648
rect 11006 7584 11022 7648
rect 11086 7584 11102 7648
rect 11166 7584 11174 7648
rect 10854 7583 11174 7584
rect 13954 7648 14274 7649
rect 13954 7584 13962 7648
rect 14026 7584 14042 7648
rect 14106 7584 14122 7648
rect 14186 7584 14202 7648
rect 14266 7584 14274 7648
rect 13954 7583 14274 7584
rect 17054 7648 17374 7649
rect 17054 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17222 7648
rect 17286 7584 17302 7648
rect 17366 7584 17374 7648
rect 17054 7583 17374 7584
rect 13445 7442 13511 7445
rect 14549 7442 14615 7445
rect 13445 7440 14615 7442
rect 13445 7384 13450 7440
rect 13506 7384 14554 7440
rect 14610 7384 14615 7440
rect 13445 7382 14615 7384
rect 13445 7379 13511 7382
rect 14549 7379 14615 7382
rect 13261 7306 13327 7309
rect 14733 7306 14799 7309
rect 13261 7304 14799 7306
rect 13261 7248 13266 7304
rect 13322 7248 14738 7304
rect 14794 7248 14799 7304
rect 13261 7246 14799 7248
rect 13261 7243 13327 7246
rect 14733 7243 14799 7246
rect 3104 7104 3424 7105
rect 3104 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3272 7104
rect 3336 7040 3352 7104
rect 3416 7040 3424 7104
rect 3104 7039 3424 7040
rect 6204 7104 6524 7105
rect 6204 7040 6212 7104
rect 6276 7040 6292 7104
rect 6356 7040 6372 7104
rect 6436 7040 6452 7104
rect 6516 7040 6524 7104
rect 6204 7039 6524 7040
rect 9304 7104 9624 7105
rect 9304 7040 9312 7104
rect 9376 7040 9392 7104
rect 9456 7040 9472 7104
rect 9536 7040 9552 7104
rect 9616 7040 9624 7104
rect 9304 7039 9624 7040
rect 12404 7104 12724 7105
rect 12404 7040 12412 7104
rect 12476 7040 12492 7104
rect 12556 7040 12572 7104
rect 12636 7040 12652 7104
rect 12716 7040 12724 7104
rect 12404 7039 12724 7040
rect 15504 7104 15824 7105
rect 15504 7040 15512 7104
rect 15576 7040 15592 7104
rect 15656 7040 15672 7104
rect 15736 7040 15752 7104
rect 15816 7040 15824 7104
rect 15504 7039 15824 7040
rect 11605 6762 11671 6765
rect 15009 6762 15075 6765
rect 11605 6760 15075 6762
rect 11605 6704 11610 6760
rect 11666 6704 15014 6760
rect 15070 6704 15075 6760
rect 11605 6702 15075 6704
rect 11605 6699 11671 6702
rect 15009 6699 15075 6702
rect 18505 6762 18571 6765
rect 19200 6762 20000 6792
rect 18505 6760 20000 6762
rect 18505 6704 18510 6760
rect 18566 6704 20000 6760
rect 18505 6702 20000 6704
rect 18505 6699 18571 6702
rect 19200 6672 20000 6702
rect 4654 6560 4974 6561
rect 4654 6496 4662 6560
rect 4726 6496 4742 6560
rect 4806 6496 4822 6560
rect 4886 6496 4902 6560
rect 4966 6496 4974 6560
rect 4654 6495 4974 6496
rect 7754 6560 8074 6561
rect 7754 6496 7762 6560
rect 7826 6496 7842 6560
rect 7906 6496 7922 6560
rect 7986 6496 8002 6560
rect 8066 6496 8074 6560
rect 7754 6495 8074 6496
rect 10854 6560 11174 6561
rect 10854 6496 10862 6560
rect 10926 6496 10942 6560
rect 11006 6496 11022 6560
rect 11086 6496 11102 6560
rect 11166 6496 11174 6560
rect 10854 6495 11174 6496
rect 13954 6560 14274 6561
rect 13954 6496 13962 6560
rect 14026 6496 14042 6560
rect 14106 6496 14122 6560
rect 14186 6496 14202 6560
rect 14266 6496 14274 6560
rect 13954 6495 14274 6496
rect 17054 6560 17374 6561
rect 17054 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17222 6560
rect 17286 6496 17302 6560
rect 17366 6496 17374 6560
rect 17054 6495 17374 6496
rect 3104 6016 3424 6017
rect 3104 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3272 6016
rect 3336 5952 3352 6016
rect 3416 5952 3424 6016
rect 3104 5951 3424 5952
rect 6204 6016 6524 6017
rect 6204 5952 6212 6016
rect 6276 5952 6292 6016
rect 6356 5952 6372 6016
rect 6436 5952 6452 6016
rect 6516 5952 6524 6016
rect 6204 5951 6524 5952
rect 9304 6016 9624 6017
rect 9304 5952 9312 6016
rect 9376 5952 9392 6016
rect 9456 5952 9472 6016
rect 9536 5952 9552 6016
rect 9616 5952 9624 6016
rect 9304 5951 9624 5952
rect 12404 6016 12724 6017
rect 12404 5952 12412 6016
rect 12476 5952 12492 6016
rect 12556 5952 12572 6016
rect 12636 5952 12652 6016
rect 12716 5952 12724 6016
rect 12404 5951 12724 5952
rect 15504 6016 15824 6017
rect 15504 5952 15512 6016
rect 15576 5952 15592 6016
rect 15656 5952 15672 6016
rect 15736 5952 15752 6016
rect 15816 5952 15824 6016
rect 15504 5951 15824 5952
rect 13721 5810 13787 5813
rect 17401 5810 17467 5813
rect 13721 5808 17467 5810
rect 13721 5752 13726 5808
rect 13782 5752 17406 5808
rect 17462 5752 17467 5808
rect 13721 5750 17467 5752
rect 13721 5747 13787 5750
rect 17401 5747 17467 5750
rect 4654 5472 4974 5473
rect 4654 5408 4662 5472
rect 4726 5408 4742 5472
rect 4806 5408 4822 5472
rect 4886 5408 4902 5472
rect 4966 5408 4974 5472
rect 4654 5407 4974 5408
rect 7754 5472 8074 5473
rect 7754 5408 7762 5472
rect 7826 5408 7842 5472
rect 7906 5408 7922 5472
rect 7986 5408 8002 5472
rect 8066 5408 8074 5472
rect 7754 5407 8074 5408
rect 10854 5472 11174 5473
rect 10854 5408 10862 5472
rect 10926 5408 10942 5472
rect 11006 5408 11022 5472
rect 11086 5408 11102 5472
rect 11166 5408 11174 5472
rect 10854 5407 11174 5408
rect 13954 5472 14274 5473
rect 13954 5408 13962 5472
rect 14026 5408 14042 5472
rect 14106 5408 14122 5472
rect 14186 5408 14202 5472
rect 14266 5408 14274 5472
rect 13954 5407 14274 5408
rect 17054 5472 17374 5473
rect 17054 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17222 5472
rect 17286 5408 17302 5472
rect 17366 5408 17374 5472
rect 17054 5407 17374 5408
rect 18505 5266 18571 5269
rect 19200 5266 20000 5296
rect 18505 5264 20000 5266
rect 18505 5208 18510 5264
rect 18566 5208 20000 5264
rect 18505 5206 20000 5208
rect 18505 5203 18571 5206
rect 19200 5176 20000 5206
rect 3104 4928 3424 4929
rect 3104 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3272 4928
rect 3336 4864 3352 4928
rect 3416 4864 3424 4928
rect 3104 4863 3424 4864
rect 6204 4928 6524 4929
rect 6204 4864 6212 4928
rect 6276 4864 6292 4928
rect 6356 4864 6372 4928
rect 6436 4864 6452 4928
rect 6516 4864 6524 4928
rect 6204 4863 6524 4864
rect 9304 4928 9624 4929
rect 9304 4864 9312 4928
rect 9376 4864 9392 4928
rect 9456 4864 9472 4928
rect 9536 4864 9552 4928
rect 9616 4864 9624 4928
rect 9304 4863 9624 4864
rect 12404 4928 12724 4929
rect 12404 4864 12412 4928
rect 12476 4864 12492 4928
rect 12556 4864 12572 4928
rect 12636 4864 12652 4928
rect 12716 4864 12724 4928
rect 12404 4863 12724 4864
rect 15504 4928 15824 4929
rect 15504 4864 15512 4928
rect 15576 4864 15592 4928
rect 15656 4864 15672 4928
rect 15736 4864 15752 4928
rect 15816 4864 15824 4928
rect 15504 4863 15824 4864
rect 4654 4384 4974 4385
rect 4654 4320 4662 4384
rect 4726 4320 4742 4384
rect 4806 4320 4822 4384
rect 4886 4320 4902 4384
rect 4966 4320 4974 4384
rect 4654 4319 4974 4320
rect 7754 4384 8074 4385
rect 7754 4320 7762 4384
rect 7826 4320 7842 4384
rect 7906 4320 7922 4384
rect 7986 4320 8002 4384
rect 8066 4320 8074 4384
rect 7754 4319 8074 4320
rect 10854 4384 11174 4385
rect 10854 4320 10862 4384
rect 10926 4320 10942 4384
rect 11006 4320 11022 4384
rect 11086 4320 11102 4384
rect 11166 4320 11174 4384
rect 10854 4319 11174 4320
rect 13954 4384 14274 4385
rect 13954 4320 13962 4384
rect 14026 4320 14042 4384
rect 14106 4320 14122 4384
rect 14186 4320 14202 4384
rect 14266 4320 14274 4384
rect 13954 4319 14274 4320
rect 17054 4384 17374 4385
rect 17054 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17222 4384
rect 17286 4320 17302 4384
rect 17366 4320 17374 4384
rect 17054 4319 17374 4320
rect 3049 4178 3115 4181
rect 3509 4178 3575 4181
rect 4981 4178 5047 4181
rect 3049 4176 5047 4178
rect 3049 4120 3054 4176
rect 3110 4120 3514 4176
rect 3570 4120 4986 4176
rect 5042 4120 5047 4176
rect 3049 4118 5047 4120
rect 3049 4115 3115 4118
rect 3509 4115 3575 4118
rect 4981 4115 5047 4118
rect 3104 3840 3424 3841
rect 3104 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3272 3840
rect 3336 3776 3352 3840
rect 3416 3776 3424 3840
rect 3104 3775 3424 3776
rect 6204 3840 6524 3841
rect 6204 3776 6212 3840
rect 6276 3776 6292 3840
rect 6356 3776 6372 3840
rect 6436 3776 6452 3840
rect 6516 3776 6524 3840
rect 6204 3775 6524 3776
rect 9304 3840 9624 3841
rect 9304 3776 9312 3840
rect 9376 3776 9392 3840
rect 9456 3776 9472 3840
rect 9536 3776 9552 3840
rect 9616 3776 9624 3840
rect 9304 3775 9624 3776
rect 12404 3840 12724 3841
rect 12404 3776 12412 3840
rect 12476 3776 12492 3840
rect 12556 3776 12572 3840
rect 12636 3776 12652 3840
rect 12716 3776 12724 3840
rect 12404 3775 12724 3776
rect 15504 3840 15824 3841
rect 15504 3776 15512 3840
rect 15576 3776 15592 3840
rect 15656 3776 15672 3840
rect 15736 3776 15752 3840
rect 15816 3776 15824 3840
rect 15504 3775 15824 3776
rect 18505 3770 18571 3773
rect 19200 3770 20000 3800
rect 18505 3768 20000 3770
rect 18505 3712 18510 3768
rect 18566 3712 20000 3768
rect 18505 3710 20000 3712
rect 18505 3707 18571 3710
rect 19200 3680 20000 3710
rect 4654 3296 4974 3297
rect 4654 3232 4662 3296
rect 4726 3232 4742 3296
rect 4806 3232 4822 3296
rect 4886 3232 4902 3296
rect 4966 3232 4974 3296
rect 4654 3231 4974 3232
rect 7754 3296 8074 3297
rect 7754 3232 7762 3296
rect 7826 3232 7842 3296
rect 7906 3232 7922 3296
rect 7986 3232 8002 3296
rect 8066 3232 8074 3296
rect 7754 3231 8074 3232
rect 10854 3296 11174 3297
rect 10854 3232 10862 3296
rect 10926 3232 10942 3296
rect 11006 3232 11022 3296
rect 11086 3232 11102 3296
rect 11166 3232 11174 3296
rect 10854 3231 11174 3232
rect 13954 3296 14274 3297
rect 13954 3232 13962 3296
rect 14026 3232 14042 3296
rect 14106 3232 14122 3296
rect 14186 3232 14202 3296
rect 14266 3232 14274 3296
rect 13954 3231 14274 3232
rect 17054 3296 17374 3297
rect 17054 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17222 3296
rect 17286 3232 17302 3296
rect 17366 3232 17374 3296
rect 17054 3231 17374 3232
rect 3104 2752 3424 2753
rect 3104 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3272 2752
rect 3336 2688 3352 2752
rect 3416 2688 3424 2752
rect 3104 2687 3424 2688
rect 6204 2752 6524 2753
rect 6204 2688 6212 2752
rect 6276 2688 6292 2752
rect 6356 2688 6372 2752
rect 6436 2688 6452 2752
rect 6516 2688 6524 2752
rect 6204 2687 6524 2688
rect 9304 2752 9624 2753
rect 9304 2688 9312 2752
rect 9376 2688 9392 2752
rect 9456 2688 9472 2752
rect 9536 2688 9552 2752
rect 9616 2688 9624 2752
rect 9304 2687 9624 2688
rect 12404 2752 12724 2753
rect 12404 2688 12412 2752
rect 12476 2688 12492 2752
rect 12556 2688 12572 2752
rect 12636 2688 12652 2752
rect 12716 2688 12724 2752
rect 12404 2687 12724 2688
rect 15504 2752 15824 2753
rect 15504 2688 15512 2752
rect 15576 2688 15592 2752
rect 15656 2688 15672 2752
rect 15736 2688 15752 2752
rect 15816 2688 15824 2752
rect 15504 2687 15824 2688
rect 7649 2410 7715 2413
rect 9029 2410 9095 2413
rect 9213 2410 9279 2413
rect 7649 2408 9279 2410
rect 7649 2352 7654 2408
rect 7710 2352 9034 2408
rect 9090 2352 9218 2408
rect 9274 2352 9279 2408
rect 7649 2350 9279 2352
rect 7649 2347 7715 2350
rect 9029 2347 9095 2350
rect 9213 2347 9279 2350
rect 18505 2274 18571 2277
rect 19200 2274 20000 2304
rect 18505 2272 20000 2274
rect 18505 2216 18510 2272
rect 18566 2216 20000 2272
rect 18505 2214 20000 2216
rect 18505 2211 18571 2214
rect 4654 2208 4974 2209
rect 4654 2144 4662 2208
rect 4726 2144 4742 2208
rect 4806 2144 4822 2208
rect 4886 2144 4902 2208
rect 4966 2144 4974 2208
rect 4654 2143 4974 2144
rect 7754 2208 8074 2209
rect 7754 2144 7762 2208
rect 7826 2144 7842 2208
rect 7906 2144 7922 2208
rect 7986 2144 8002 2208
rect 8066 2144 8074 2208
rect 7754 2143 8074 2144
rect 10854 2208 11174 2209
rect 10854 2144 10862 2208
rect 10926 2144 10942 2208
rect 11006 2144 11022 2208
rect 11086 2144 11102 2208
rect 11166 2144 11174 2208
rect 10854 2143 11174 2144
rect 13954 2208 14274 2209
rect 13954 2144 13962 2208
rect 14026 2144 14042 2208
rect 14106 2144 14122 2208
rect 14186 2144 14202 2208
rect 14266 2144 14274 2208
rect 13954 2143 14274 2144
rect 17054 2208 17374 2209
rect 17054 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17222 2208
rect 17286 2144 17302 2208
rect 17366 2144 17374 2208
rect 19200 2184 20000 2214
rect 17054 2143 17374 2144
rect 3104 1664 3424 1665
rect 3104 1600 3112 1664
rect 3176 1600 3192 1664
rect 3256 1600 3272 1664
rect 3336 1600 3352 1664
rect 3416 1600 3424 1664
rect 3104 1599 3424 1600
rect 6204 1664 6524 1665
rect 6204 1600 6212 1664
rect 6276 1600 6292 1664
rect 6356 1600 6372 1664
rect 6436 1600 6452 1664
rect 6516 1600 6524 1664
rect 6204 1599 6524 1600
rect 9304 1664 9624 1665
rect 9304 1600 9312 1664
rect 9376 1600 9392 1664
rect 9456 1600 9472 1664
rect 9536 1600 9552 1664
rect 9616 1600 9624 1664
rect 9304 1599 9624 1600
rect 12404 1664 12724 1665
rect 12404 1600 12412 1664
rect 12476 1600 12492 1664
rect 12556 1600 12572 1664
rect 12636 1600 12652 1664
rect 12716 1600 12724 1664
rect 12404 1599 12724 1600
rect 15504 1664 15824 1665
rect 15504 1600 15512 1664
rect 15576 1600 15592 1664
rect 15656 1600 15672 1664
rect 15736 1600 15752 1664
rect 15816 1600 15824 1664
rect 15504 1599 15824 1600
rect 3601 1322 3667 1325
rect 5533 1322 5599 1325
rect 3601 1320 5599 1322
rect 3601 1264 3606 1320
rect 3662 1264 5538 1320
rect 5594 1264 5599 1320
rect 3601 1262 5599 1264
rect 3601 1259 3667 1262
rect 5533 1259 5599 1262
rect 4654 1120 4974 1121
rect 4654 1056 4662 1120
rect 4726 1056 4742 1120
rect 4806 1056 4822 1120
rect 4886 1056 4902 1120
rect 4966 1056 4974 1120
rect 4654 1055 4974 1056
rect 7754 1120 8074 1121
rect 7754 1056 7762 1120
rect 7826 1056 7842 1120
rect 7906 1056 7922 1120
rect 7986 1056 8002 1120
rect 8066 1056 8074 1120
rect 7754 1055 8074 1056
rect 10854 1120 11174 1121
rect 10854 1056 10862 1120
rect 10926 1056 10942 1120
rect 11006 1056 11022 1120
rect 11086 1056 11102 1120
rect 11166 1056 11174 1120
rect 10854 1055 11174 1056
rect 13954 1120 14274 1121
rect 13954 1056 13962 1120
rect 14026 1056 14042 1120
rect 14106 1056 14122 1120
rect 14186 1056 14202 1120
rect 14266 1056 14274 1120
rect 13954 1055 14274 1056
rect 17054 1120 17374 1121
rect 17054 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17222 1120
rect 17286 1056 17302 1120
rect 17366 1056 17374 1120
rect 17054 1055 17374 1056
rect 11789 914 11855 917
rect 13813 914 13879 917
rect 11789 912 13879 914
rect 11789 856 11794 912
rect 11850 856 13818 912
rect 13874 856 13879 912
rect 11789 854 13879 856
rect 11789 851 11855 854
rect 13813 851 13879 854
rect 6361 778 6427 781
rect 6637 778 6703 781
rect 10961 778 11027 781
rect 18137 778 18203 781
rect 6361 776 18203 778
rect 6361 720 6366 776
rect 6422 720 6642 776
rect 6698 720 10966 776
rect 11022 720 18142 776
rect 18198 720 18203 776
rect 6361 718 18203 720
rect 6361 715 6427 718
rect 6637 715 6703 718
rect 10961 715 11027 718
rect 18137 715 18203 718
rect 18505 778 18571 781
rect 19200 778 20000 808
rect 18505 776 20000 778
rect 18505 720 18510 776
rect 18566 720 20000 776
rect 18505 718 20000 720
rect 18505 715 18571 718
rect 19200 688 20000 718
rect 3104 576 3424 577
rect 3104 512 3112 576
rect 3176 512 3192 576
rect 3256 512 3272 576
rect 3336 512 3352 576
rect 3416 512 3424 576
rect 3104 511 3424 512
rect 6204 576 6524 577
rect 6204 512 6212 576
rect 6276 512 6292 576
rect 6356 512 6372 576
rect 6436 512 6452 576
rect 6516 512 6524 576
rect 6204 511 6524 512
rect 9304 576 9624 577
rect 9304 512 9312 576
rect 9376 512 9392 576
rect 9456 512 9472 576
rect 9536 512 9552 576
rect 9616 512 9624 576
rect 9304 511 9624 512
rect 12404 576 12724 577
rect 12404 512 12412 576
rect 12476 512 12492 576
rect 12556 512 12572 576
rect 12636 512 12652 576
rect 12716 512 12724 576
rect 12404 511 12724 512
rect 15504 576 15824 577
rect 15504 512 15512 576
rect 15576 512 15592 576
rect 15656 512 15672 576
rect 15736 512 15752 576
rect 15816 512 15824 576
rect 15504 511 15824 512
rect 14641 370 14707 373
rect 17953 370 18019 373
rect 14641 368 18019 370
rect 14641 312 14646 368
rect 14702 312 17958 368
rect 18014 312 18019 368
rect 14641 310 18019 312
rect 14641 307 14707 310
rect 17953 307 18019 310
rect 8661 234 8727 237
rect 12617 234 12683 237
rect 8661 232 12683 234
rect 8661 176 8666 232
rect 8722 176 12622 232
rect 12678 176 12683 232
rect 8661 174 12683 176
rect 8661 171 8727 174
rect 12617 171 12683 174
rect 4654 32 4974 33
rect 4654 -32 4662 32
rect 4726 -32 4742 32
rect 4806 -32 4822 32
rect 4886 -32 4902 32
rect 4966 -32 4974 32
rect 4654 -33 4974 -32
rect 7754 32 8074 33
rect 7754 -32 7762 32
rect 7826 -32 7842 32
rect 7906 -32 7922 32
rect 7986 -32 8002 32
rect 8066 -32 8074 32
rect 7754 -33 8074 -32
rect 10854 32 11174 33
rect 10854 -32 10862 32
rect 10926 -32 10942 32
rect 11006 -32 11022 32
rect 11086 -32 11102 32
rect 11166 -32 11174 32
rect 10854 -33 11174 -32
rect 13954 32 14274 33
rect 13954 -32 13962 32
rect 14026 -32 14042 32
rect 14106 -32 14122 32
rect 14186 -32 14202 32
rect 14266 -32 14274 32
rect 13954 -33 14274 -32
rect 17054 32 17374 33
rect 17054 -32 17062 32
rect 17126 -32 17142 32
rect 17206 -32 17222 32
rect 17286 -32 17302 32
rect 17366 -32 17374 32
rect 17054 -33 17374 -32
<< via3 >>
rect 4662 10908 4726 10912
rect 4662 10852 4666 10908
rect 4666 10852 4722 10908
rect 4722 10852 4726 10908
rect 4662 10848 4726 10852
rect 4742 10908 4806 10912
rect 4742 10852 4746 10908
rect 4746 10852 4802 10908
rect 4802 10852 4806 10908
rect 4742 10848 4806 10852
rect 4822 10908 4886 10912
rect 4822 10852 4826 10908
rect 4826 10852 4882 10908
rect 4882 10852 4886 10908
rect 4822 10848 4886 10852
rect 4902 10908 4966 10912
rect 4902 10852 4906 10908
rect 4906 10852 4962 10908
rect 4962 10852 4966 10908
rect 4902 10848 4966 10852
rect 7762 10908 7826 10912
rect 7762 10852 7766 10908
rect 7766 10852 7822 10908
rect 7822 10852 7826 10908
rect 7762 10848 7826 10852
rect 7842 10908 7906 10912
rect 7842 10852 7846 10908
rect 7846 10852 7902 10908
rect 7902 10852 7906 10908
rect 7842 10848 7906 10852
rect 7922 10908 7986 10912
rect 7922 10852 7926 10908
rect 7926 10852 7982 10908
rect 7982 10852 7986 10908
rect 7922 10848 7986 10852
rect 8002 10908 8066 10912
rect 8002 10852 8006 10908
rect 8006 10852 8062 10908
rect 8062 10852 8066 10908
rect 8002 10848 8066 10852
rect 10862 10908 10926 10912
rect 10862 10852 10866 10908
rect 10866 10852 10922 10908
rect 10922 10852 10926 10908
rect 10862 10848 10926 10852
rect 10942 10908 11006 10912
rect 10942 10852 10946 10908
rect 10946 10852 11002 10908
rect 11002 10852 11006 10908
rect 10942 10848 11006 10852
rect 11022 10908 11086 10912
rect 11022 10852 11026 10908
rect 11026 10852 11082 10908
rect 11082 10852 11086 10908
rect 11022 10848 11086 10852
rect 11102 10908 11166 10912
rect 11102 10852 11106 10908
rect 11106 10852 11162 10908
rect 11162 10852 11166 10908
rect 11102 10848 11166 10852
rect 13962 10908 14026 10912
rect 13962 10852 13966 10908
rect 13966 10852 14022 10908
rect 14022 10852 14026 10908
rect 13962 10848 14026 10852
rect 14042 10908 14106 10912
rect 14042 10852 14046 10908
rect 14046 10852 14102 10908
rect 14102 10852 14106 10908
rect 14042 10848 14106 10852
rect 14122 10908 14186 10912
rect 14122 10852 14126 10908
rect 14126 10852 14182 10908
rect 14182 10852 14186 10908
rect 14122 10848 14186 10852
rect 14202 10908 14266 10912
rect 14202 10852 14206 10908
rect 14206 10852 14262 10908
rect 14262 10852 14266 10908
rect 14202 10848 14266 10852
rect 17062 10908 17126 10912
rect 17062 10852 17066 10908
rect 17066 10852 17122 10908
rect 17122 10852 17126 10908
rect 17062 10848 17126 10852
rect 17142 10908 17206 10912
rect 17142 10852 17146 10908
rect 17146 10852 17202 10908
rect 17202 10852 17206 10908
rect 17142 10848 17206 10852
rect 17222 10908 17286 10912
rect 17222 10852 17226 10908
rect 17226 10852 17282 10908
rect 17282 10852 17286 10908
rect 17222 10848 17286 10852
rect 17302 10908 17366 10912
rect 17302 10852 17306 10908
rect 17306 10852 17362 10908
rect 17362 10852 17366 10908
rect 17302 10848 17366 10852
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 3272 10364 3336 10368
rect 3272 10308 3276 10364
rect 3276 10308 3332 10364
rect 3332 10308 3336 10364
rect 3272 10304 3336 10308
rect 3352 10364 3416 10368
rect 3352 10308 3356 10364
rect 3356 10308 3412 10364
rect 3412 10308 3416 10364
rect 3352 10304 3416 10308
rect 6212 10364 6276 10368
rect 6212 10308 6216 10364
rect 6216 10308 6272 10364
rect 6272 10308 6276 10364
rect 6212 10304 6276 10308
rect 6292 10364 6356 10368
rect 6292 10308 6296 10364
rect 6296 10308 6352 10364
rect 6352 10308 6356 10364
rect 6292 10304 6356 10308
rect 6372 10364 6436 10368
rect 6372 10308 6376 10364
rect 6376 10308 6432 10364
rect 6432 10308 6436 10364
rect 6372 10304 6436 10308
rect 6452 10364 6516 10368
rect 6452 10308 6456 10364
rect 6456 10308 6512 10364
rect 6512 10308 6516 10364
rect 6452 10304 6516 10308
rect 9312 10364 9376 10368
rect 9312 10308 9316 10364
rect 9316 10308 9372 10364
rect 9372 10308 9376 10364
rect 9312 10304 9376 10308
rect 9392 10364 9456 10368
rect 9392 10308 9396 10364
rect 9396 10308 9452 10364
rect 9452 10308 9456 10364
rect 9392 10304 9456 10308
rect 9472 10364 9536 10368
rect 9472 10308 9476 10364
rect 9476 10308 9532 10364
rect 9532 10308 9536 10364
rect 9472 10304 9536 10308
rect 9552 10364 9616 10368
rect 9552 10308 9556 10364
rect 9556 10308 9612 10364
rect 9612 10308 9616 10364
rect 9552 10304 9616 10308
rect 12412 10364 12476 10368
rect 12412 10308 12416 10364
rect 12416 10308 12472 10364
rect 12472 10308 12476 10364
rect 12412 10304 12476 10308
rect 12492 10364 12556 10368
rect 12492 10308 12496 10364
rect 12496 10308 12552 10364
rect 12552 10308 12556 10364
rect 12492 10304 12556 10308
rect 12572 10364 12636 10368
rect 12572 10308 12576 10364
rect 12576 10308 12632 10364
rect 12632 10308 12636 10364
rect 12572 10304 12636 10308
rect 12652 10364 12716 10368
rect 12652 10308 12656 10364
rect 12656 10308 12712 10364
rect 12712 10308 12716 10364
rect 12652 10304 12716 10308
rect 15512 10364 15576 10368
rect 15512 10308 15516 10364
rect 15516 10308 15572 10364
rect 15572 10308 15576 10364
rect 15512 10304 15576 10308
rect 15592 10364 15656 10368
rect 15592 10308 15596 10364
rect 15596 10308 15652 10364
rect 15652 10308 15656 10364
rect 15592 10304 15656 10308
rect 15672 10364 15736 10368
rect 15672 10308 15676 10364
rect 15676 10308 15732 10364
rect 15732 10308 15736 10364
rect 15672 10304 15736 10308
rect 15752 10364 15816 10368
rect 15752 10308 15756 10364
rect 15756 10308 15812 10364
rect 15812 10308 15816 10364
rect 15752 10304 15816 10308
rect 4662 9820 4726 9824
rect 4662 9764 4666 9820
rect 4666 9764 4722 9820
rect 4722 9764 4726 9820
rect 4662 9760 4726 9764
rect 4742 9820 4806 9824
rect 4742 9764 4746 9820
rect 4746 9764 4802 9820
rect 4802 9764 4806 9820
rect 4742 9760 4806 9764
rect 4822 9820 4886 9824
rect 4822 9764 4826 9820
rect 4826 9764 4882 9820
rect 4882 9764 4886 9820
rect 4822 9760 4886 9764
rect 4902 9820 4966 9824
rect 4902 9764 4906 9820
rect 4906 9764 4962 9820
rect 4962 9764 4966 9820
rect 4902 9760 4966 9764
rect 7762 9820 7826 9824
rect 7762 9764 7766 9820
rect 7766 9764 7822 9820
rect 7822 9764 7826 9820
rect 7762 9760 7826 9764
rect 7842 9820 7906 9824
rect 7842 9764 7846 9820
rect 7846 9764 7902 9820
rect 7902 9764 7906 9820
rect 7842 9760 7906 9764
rect 7922 9820 7986 9824
rect 7922 9764 7926 9820
rect 7926 9764 7982 9820
rect 7982 9764 7986 9820
rect 7922 9760 7986 9764
rect 8002 9820 8066 9824
rect 8002 9764 8006 9820
rect 8006 9764 8062 9820
rect 8062 9764 8066 9820
rect 8002 9760 8066 9764
rect 10862 9820 10926 9824
rect 10862 9764 10866 9820
rect 10866 9764 10922 9820
rect 10922 9764 10926 9820
rect 10862 9760 10926 9764
rect 10942 9820 11006 9824
rect 10942 9764 10946 9820
rect 10946 9764 11002 9820
rect 11002 9764 11006 9820
rect 10942 9760 11006 9764
rect 11022 9820 11086 9824
rect 11022 9764 11026 9820
rect 11026 9764 11082 9820
rect 11082 9764 11086 9820
rect 11022 9760 11086 9764
rect 11102 9820 11166 9824
rect 11102 9764 11106 9820
rect 11106 9764 11162 9820
rect 11162 9764 11166 9820
rect 11102 9760 11166 9764
rect 13962 9820 14026 9824
rect 13962 9764 13966 9820
rect 13966 9764 14022 9820
rect 14022 9764 14026 9820
rect 13962 9760 14026 9764
rect 14042 9820 14106 9824
rect 14042 9764 14046 9820
rect 14046 9764 14102 9820
rect 14102 9764 14106 9820
rect 14042 9760 14106 9764
rect 14122 9820 14186 9824
rect 14122 9764 14126 9820
rect 14126 9764 14182 9820
rect 14182 9764 14186 9820
rect 14122 9760 14186 9764
rect 14202 9820 14266 9824
rect 14202 9764 14206 9820
rect 14206 9764 14262 9820
rect 14262 9764 14266 9820
rect 14202 9760 14266 9764
rect 17062 9820 17126 9824
rect 17062 9764 17066 9820
rect 17066 9764 17122 9820
rect 17122 9764 17126 9820
rect 17062 9760 17126 9764
rect 17142 9820 17206 9824
rect 17142 9764 17146 9820
rect 17146 9764 17202 9820
rect 17202 9764 17206 9820
rect 17142 9760 17206 9764
rect 17222 9820 17286 9824
rect 17222 9764 17226 9820
rect 17226 9764 17282 9820
rect 17282 9764 17286 9820
rect 17222 9760 17286 9764
rect 17302 9820 17366 9824
rect 17302 9764 17306 9820
rect 17306 9764 17362 9820
rect 17362 9764 17366 9820
rect 17302 9760 17366 9764
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 3272 9276 3336 9280
rect 3272 9220 3276 9276
rect 3276 9220 3332 9276
rect 3332 9220 3336 9276
rect 3272 9216 3336 9220
rect 3352 9276 3416 9280
rect 3352 9220 3356 9276
rect 3356 9220 3412 9276
rect 3412 9220 3416 9276
rect 3352 9216 3416 9220
rect 6212 9276 6276 9280
rect 6212 9220 6216 9276
rect 6216 9220 6272 9276
rect 6272 9220 6276 9276
rect 6212 9216 6276 9220
rect 6292 9276 6356 9280
rect 6292 9220 6296 9276
rect 6296 9220 6352 9276
rect 6352 9220 6356 9276
rect 6292 9216 6356 9220
rect 6372 9276 6436 9280
rect 6372 9220 6376 9276
rect 6376 9220 6432 9276
rect 6432 9220 6436 9276
rect 6372 9216 6436 9220
rect 6452 9276 6516 9280
rect 6452 9220 6456 9276
rect 6456 9220 6512 9276
rect 6512 9220 6516 9276
rect 6452 9216 6516 9220
rect 9312 9276 9376 9280
rect 9312 9220 9316 9276
rect 9316 9220 9372 9276
rect 9372 9220 9376 9276
rect 9312 9216 9376 9220
rect 9392 9276 9456 9280
rect 9392 9220 9396 9276
rect 9396 9220 9452 9276
rect 9452 9220 9456 9276
rect 9392 9216 9456 9220
rect 9472 9276 9536 9280
rect 9472 9220 9476 9276
rect 9476 9220 9532 9276
rect 9532 9220 9536 9276
rect 9472 9216 9536 9220
rect 9552 9276 9616 9280
rect 9552 9220 9556 9276
rect 9556 9220 9612 9276
rect 9612 9220 9616 9276
rect 9552 9216 9616 9220
rect 12412 9276 12476 9280
rect 12412 9220 12416 9276
rect 12416 9220 12472 9276
rect 12472 9220 12476 9276
rect 12412 9216 12476 9220
rect 12492 9276 12556 9280
rect 12492 9220 12496 9276
rect 12496 9220 12552 9276
rect 12552 9220 12556 9276
rect 12492 9216 12556 9220
rect 12572 9276 12636 9280
rect 12572 9220 12576 9276
rect 12576 9220 12632 9276
rect 12632 9220 12636 9276
rect 12572 9216 12636 9220
rect 12652 9276 12716 9280
rect 12652 9220 12656 9276
rect 12656 9220 12712 9276
rect 12712 9220 12716 9276
rect 12652 9216 12716 9220
rect 15512 9276 15576 9280
rect 15512 9220 15516 9276
rect 15516 9220 15572 9276
rect 15572 9220 15576 9276
rect 15512 9216 15576 9220
rect 15592 9276 15656 9280
rect 15592 9220 15596 9276
rect 15596 9220 15652 9276
rect 15652 9220 15656 9276
rect 15592 9216 15656 9220
rect 15672 9276 15736 9280
rect 15672 9220 15676 9276
rect 15676 9220 15732 9276
rect 15732 9220 15736 9276
rect 15672 9216 15736 9220
rect 15752 9276 15816 9280
rect 15752 9220 15756 9276
rect 15756 9220 15812 9276
rect 15812 9220 15816 9276
rect 15752 9216 15816 9220
rect 4662 8732 4726 8736
rect 4662 8676 4666 8732
rect 4666 8676 4722 8732
rect 4722 8676 4726 8732
rect 4662 8672 4726 8676
rect 4742 8732 4806 8736
rect 4742 8676 4746 8732
rect 4746 8676 4802 8732
rect 4802 8676 4806 8732
rect 4742 8672 4806 8676
rect 4822 8732 4886 8736
rect 4822 8676 4826 8732
rect 4826 8676 4882 8732
rect 4882 8676 4886 8732
rect 4822 8672 4886 8676
rect 4902 8732 4966 8736
rect 4902 8676 4906 8732
rect 4906 8676 4962 8732
rect 4962 8676 4966 8732
rect 4902 8672 4966 8676
rect 7762 8732 7826 8736
rect 7762 8676 7766 8732
rect 7766 8676 7822 8732
rect 7822 8676 7826 8732
rect 7762 8672 7826 8676
rect 7842 8732 7906 8736
rect 7842 8676 7846 8732
rect 7846 8676 7902 8732
rect 7902 8676 7906 8732
rect 7842 8672 7906 8676
rect 7922 8732 7986 8736
rect 7922 8676 7926 8732
rect 7926 8676 7982 8732
rect 7982 8676 7986 8732
rect 7922 8672 7986 8676
rect 8002 8732 8066 8736
rect 8002 8676 8006 8732
rect 8006 8676 8062 8732
rect 8062 8676 8066 8732
rect 8002 8672 8066 8676
rect 10862 8732 10926 8736
rect 10862 8676 10866 8732
rect 10866 8676 10922 8732
rect 10922 8676 10926 8732
rect 10862 8672 10926 8676
rect 10942 8732 11006 8736
rect 10942 8676 10946 8732
rect 10946 8676 11002 8732
rect 11002 8676 11006 8732
rect 10942 8672 11006 8676
rect 11022 8732 11086 8736
rect 11022 8676 11026 8732
rect 11026 8676 11082 8732
rect 11082 8676 11086 8732
rect 11022 8672 11086 8676
rect 11102 8732 11166 8736
rect 11102 8676 11106 8732
rect 11106 8676 11162 8732
rect 11162 8676 11166 8732
rect 11102 8672 11166 8676
rect 13962 8732 14026 8736
rect 13962 8676 13966 8732
rect 13966 8676 14022 8732
rect 14022 8676 14026 8732
rect 13962 8672 14026 8676
rect 14042 8732 14106 8736
rect 14042 8676 14046 8732
rect 14046 8676 14102 8732
rect 14102 8676 14106 8732
rect 14042 8672 14106 8676
rect 14122 8732 14186 8736
rect 14122 8676 14126 8732
rect 14126 8676 14182 8732
rect 14182 8676 14186 8732
rect 14122 8672 14186 8676
rect 14202 8732 14266 8736
rect 14202 8676 14206 8732
rect 14206 8676 14262 8732
rect 14262 8676 14266 8732
rect 14202 8672 14266 8676
rect 17062 8732 17126 8736
rect 17062 8676 17066 8732
rect 17066 8676 17122 8732
rect 17122 8676 17126 8732
rect 17062 8672 17126 8676
rect 17142 8732 17206 8736
rect 17142 8676 17146 8732
rect 17146 8676 17202 8732
rect 17202 8676 17206 8732
rect 17142 8672 17206 8676
rect 17222 8732 17286 8736
rect 17222 8676 17226 8732
rect 17226 8676 17282 8732
rect 17282 8676 17286 8732
rect 17222 8672 17286 8676
rect 17302 8732 17366 8736
rect 17302 8676 17306 8732
rect 17306 8676 17362 8732
rect 17362 8676 17366 8732
rect 17302 8672 17366 8676
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 3272 8188 3336 8192
rect 3272 8132 3276 8188
rect 3276 8132 3332 8188
rect 3332 8132 3336 8188
rect 3272 8128 3336 8132
rect 3352 8188 3416 8192
rect 3352 8132 3356 8188
rect 3356 8132 3412 8188
rect 3412 8132 3416 8188
rect 3352 8128 3416 8132
rect 6212 8188 6276 8192
rect 6212 8132 6216 8188
rect 6216 8132 6272 8188
rect 6272 8132 6276 8188
rect 6212 8128 6276 8132
rect 6292 8188 6356 8192
rect 6292 8132 6296 8188
rect 6296 8132 6352 8188
rect 6352 8132 6356 8188
rect 6292 8128 6356 8132
rect 6372 8188 6436 8192
rect 6372 8132 6376 8188
rect 6376 8132 6432 8188
rect 6432 8132 6436 8188
rect 6372 8128 6436 8132
rect 6452 8188 6516 8192
rect 6452 8132 6456 8188
rect 6456 8132 6512 8188
rect 6512 8132 6516 8188
rect 6452 8128 6516 8132
rect 9312 8188 9376 8192
rect 9312 8132 9316 8188
rect 9316 8132 9372 8188
rect 9372 8132 9376 8188
rect 9312 8128 9376 8132
rect 9392 8188 9456 8192
rect 9392 8132 9396 8188
rect 9396 8132 9452 8188
rect 9452 8132 9456 8188
rect 9392 8128 9456 8132
rect 9472 8188 9536 8192
rect 9472 8132 9476 8188
rect 9476 8132 9532 8188
rect 9532 8132 9536 8188
rect 9472 8128 9536 8132
rect 9552 8188 9616 8192
rect 9552 8132 9556 8188
rect 9556 8132 9612 8188
rect 9612 8132 9616 8188
rect 9552 8128 9616 8132
rect 12412 8188 12476 8192
rect 12412 8132 12416 8188
rect 12416 8132 12472 8188
rect 12472 8132 12476 8188
rect 12412 8128 12476 8132
rect 12492 8188 12556 8192
rect 12492 8132 12496 8188
rect 12496 8132 12552 8188
rect 12552 8132 12556 8188
rect 12492 8128 12556 8132
rect 12572 8188 12636 8192
rect 12572 8132 12576 8188
rect 12576 8132 12632 8188
rect 12632 8132 12636 8188
rect 12572 8128 12636 8132
rect 12652 8188 12716 8192
rect 12652 8132 12656 8188
rect 12656 8132 12712 8188
rect 12712 8132 12716 8188
rect 12652 8128 12716 8132
rect 15512 8188 15576 8192
rect 15512 8132 15516 8188
rect 15516 8132 15572 8188
rect 15572 8132 15576 8188
rect 15512 8128 15576 8132
rect 15592 8188 15656 8192
rect 15592 8132 15596 8188
rect 15596 8132 15652 8188
rect 15652 8132 15656 8188
rect 15592 8128 15656 8132
rect 15672 8188 15736 8192
rect 15672 8132 15676 8188
rect 15676 8132 15732 8188
rect 15732 8132 15736 8188
rect 15672 8128 15736 8132
rect 15752 8188 15816 8192
rect 15752 8132 15756 8188
rect 15756 8132 15812 8188
rect 15812 8132 15816 8188
rect 15752 8128 15816 8132
rect 4662 7644 4726 7648
rect 4662 7588 4666 7644
rect 4666 7588 4722 7644
rect 4722 7588 4726 7644
rect 4662 7584 4726 7588
rect 4742 7644 4806 7648
rect 4742 7588 4746 7644
rect 4746 7588 4802 7644
rect 4802 7588 4806 7644
rect 4742 7584 4806 7588
rect 4822 7644 4886 7648
rect 4822 7588 4826 7644
rect 4826 7588 4882 7644
rect 4882 7588 4886 7644
rect 4822 7584 4886 7588
rect 4902 7644 4966 7648
rect 4902 7588 4906 7644
rect 4906 7588 4962 7644
rect 4962 7588 4966 7644
rect 4902 7584 4966 7588
rect 7762 7644 7826 7648
rect 7762 7588 7766 7644
rect 7766 7588 7822 7644
rect 7822 7588 7826 7644
rect 7762 7584 7826 7588
rect 7842 7644 7906 7648
rect 7842 7588 7846 7644
rect 7846 7588 7902 7644
rect 7902 7588 7906 7644
rect 7842 7584 7906 7588
rect 7922 7644 7986 7648
rect 7922 7588 7926 7644
rect 7926 7588 7982 7644
rect 7982 7588 7986 7644
rect 7922 7584 7986 7588
rect 8002 7644 8066 7648
rect 8002 7588 8006 7644
rect 8006 7588 8062 7644
rect 8062 7588 8066 7644
rect 8002 7584 8066 7588
rect 10862 7644 10926 7648
rect 10862 7588 10866 7644
rect 10866 7588 10922 7644
rect 10922 7588 10926 7644
rect 10862 7584 10926 7588
rect 10942 7644 11006 7648
rect 10942 7588 10946 7644
rect 10946 7588 11002 7644
rect 11002 7588 11006 7644
rect 10942 7584 11006 7588
rect 11022 7644 11086 7648
rect 11022 7588 11026 7644
rect 11026 7588 11082 7644
rect 11082 7588 11086 7644
rect 11022 7584 11086 7588
rect 11102 7644 11166 7648
rect 11102 7588 11106 7644
rect 11106 7588 11162 7644
rect 11162 7588 11166 7644
rect 11102 7584 11166 7588
rect 13962 7644 14026 7648
rect 13962 7588 13966 7644
rect 13966 7588 14022 7644
rect 14022 7588 14026 7644
rect 13962 7584 14026 7588
rect 14042 7644 14106 7648
rect 14042 7588 14046 7644
rect 14046 7588 14102 7644
rect 14102 7588 14106 7644
rect 14042 7584 14106 7588
rect 14122 7644 14186 7648
rect 14122 7588 14126 7644
rect 14126 7588 14182 7644
rect 14182 7588 14186 7644
rect 14122 7584 14186 7588
rect 14202 7644 14266 7648
rect 14202 7588 14206 7644
rect 14206 7588 14262 7644
rect 14262 7588 14266 7644
rect 14202 7584 14266 7588
rect 17062 7644 17126 7648
rect 17062 7588 17066 7644
rect 17066 7588 17122 7644
rect 17122 7588 17126 7644
rect 17062 7584 17126 7588
rect 17142 7644 17206 7648
rect 17142 7588 17146 7644
rect 17146 7588 17202 7644
rect 17202 7588 17206 7644
rect 17142 7584 17206 7588
rect 17222 7644 17286 7648
rect 17222 7588 17226 7644
rect 17226 7588 17282 7644
rect 17282 7588 17286 7644
rect 17222 7584 17286 7588
rect 17302 7644 17366 7648
rect 17302 7588 17306 7644
rect 17306 7588 17362 7644
rect 17362 7588 17366 7644
rect 17302 7584 17366 7588
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 3272 7100 3336 7104
rect 3272 7044 3276 7100
rect 3276 7044 3332 7100
rect 3332 7044 3336 7100
rect 3272 7040 3336 7044
rect 3352 7100 3416 7104
rect 3352 7044 3356 7100
rect 3356 7044 3412 7100
rect 3412 7044 3416 7100
rect 3352 7040 3416 7044
rect 6212 7100 6276 7104
rect 6212 7044 6216 7100
rect 6216 7044 6272 7100
rect 6272 7044 6276 7100
rect 6212 7040 6276 7044
rect 6292 7100 6356 7104
rect 6292 7044 6296 7100
rect 6296 7044 6352 7100
rect 6352 7044 6356 7100
rect 6292 7040 6356 7044
rect 6372 7100 6436 7104
rect 6372 7044 6376 7100
rect 6376 7044 6432 7100
rect 6432 7044 6436 7100
rect 6372 7040 6436 7044
rect 6452 7100 6516 7104
rect 6452 7044 6456 7100
rect 6456 7044 6512 7100
rect 6512 7044 6516 7100
rect 6452 7040 6516 7044
rect 9312 7100 9376 7104
rect 9312 7044 9316 7100
rect 9316 7044 9372 7100
rect 9372 7044 9376 7100
rect 9312 7040 9376 7044
rect 9392 7100 9456 7104
rect 9392 7044 9396 7100
rect 9396 7044 9452 7100
rect 9452 7044 9456 7100
rect 9392 7040 9456 7044
rect 9472 7100 9536 7104
rect 9472 7044 9476 7100
rect 9476 7044 9532 7100
rect 9532 7044 9536 7100
rect 9472 7040 9536 7044
rect 9552 7100 9616 7104
rect 9552 7044 9556 7100
rect 9556 7044 9612 7100
rect 9612 7044 9616 7100
rect 9552 7040 9616 7044
rect 12412 7100 12476 7104
rect 12412 7044 12416 7100
rect 12416 7044 12472 7100
rect 12472 7044 12476 7100
rect 12412 7040 12476 7044
rect 12492 7100 12556 7104
rect 12492 7044 12496 7100
rect 12496 7044 12552 7100
rect 12552 7044 12556 7100
rect 12492 7040 12556 7044
rect 12572 7100 12636 7104
rect 12572 7044 12576 7100
rect 12576 7044 12632 7100
rect 12632 7044 12636 7100
rect 12572 7040 12636 7044
rect 12652 7100 12716 7104
rect 12652 7044 12656 7100
rect 12656 7044 12712 7100
rect 12712 7044 12716 7100
rect 12652 7040 12716 7044
rect 15512 7100 15576 7104
rect 15512 7044 15516 7100
rect 15516 7044 15572 7100
rect 15572 7044 15576 7100
rect 15512 7040 15576 7044
rect 15592 7100 15656 7104
rect 15592 7044 15596 7100
rect 15596 7044 15652 7100
rect 15652 7044 15656 7100
rect 15592 7040 15656 7044
rect 15672 7100 15736 7104
rect 15672 7044 15676 7100
rect 15676 7044 15732 7100
rect 15732 7044 15736 7100
rect 15672 7040 15736 7044
rect 15752 7100 15816 7104
rect 15752 7044 15756 7100
rect 15756 7044 15812 7100
rect 15812 7044 15816 7100
rect 15752 7040 15816 7044
rect 4662 6556 4726 6560
rect 4662 6500 4666 6556
rect 4666 6500 4722 6556
rect 4722 6500 4726 6556
rect 4662 6496 4726 6500
rect 4742 6556 4806 6560
rect 4742 6500 4746 6556
rect 4746 6500 4802 6556
rect 4802 6500 4806 6556
rect 4742 6496 4806 6500
rect 4822 6556 4886 6560
rect 4822 6500 4826 6556
rect 4826 6500 4882 6556
rect 4882 6500 4886 6556
rect 4822 6496 4886 6500
rect 4902 6556 4966 6560
rect 4902 6500 4906 6556
rect 4906 6500 4962 6556
rect 4962 6500 4966 6556
rect 4902 6496 4966 6500
rect 7762 6556 7826 6560
rect 7762 6500 7766 6556
rect 7766 6500 7822 6556
rect 7822 6500 7826 6556
rect 7762 6496 7826 6500
rect 7842 6556 7906 6560
rect 7842 6500 7846 6556
rect 7846 6500 7902 6556
rect 7902 6500 7906 6556
rect 7842 6496 7906 6500
rect 7922 6556 7986 6560
rect 7922 6500 7926 6556
rect 7926 6500 7982 6556
rect 7982 6500 7986 6556
rect 7922 6496 7986 6500
rect 8002 6556 8066 6560
rect 8002 6500 8006 6556
rect 8006 6500 8062 6556
rect 8062 6500 8066 6556
rect 8002 6496 8066 6500
rect 10862 6556 10926 6560
rect 10862 6500 10866 6556
rect 10866 6500 10922 6556
rect 10922 6500 10926 6556
rect 10862 6496 10926 6500
rect 10942 6556 11006 6560
rect 10942 6500 10946 6556
rect 10946 6500 11002 6556
rect 11002 6500 11006 6556
rect 10942 6496 11006 6500
rect 11022 6556 11086 6560
rect 11022 6500 11026 6556
rect 11026 6500 11082 6556
rect 11082 6500 11086 6556
rect 11022 6496 11086 6500
rect 11102 6556 11166 6560
rect 11102 6500 11106 6556
rect 11106 6500 11162 6556
rect 11162 6500 11166 6556
rect 11102 6496 11166 6500
rect 13962 6556 14026 6560
rect 13962 6500 13966 6556
rect 13966 6500 14022 6556
rect 14022 6500 14026 6556
rect 13962 6496 14026 6500
rect 14042 6556 14106 6560
rect 14042 6500 14046 6556
rect 14046 6500 14102 6556
rect 14102 6500 14106 6556
rect 14042 6496 14106 6500
rect 14122 6556 14186 6560
rect 14122 6500 14126 6556
rect 14126 6500 14182 6556
rect 14182 6500 14186 6556
rect 14122 6496 14186 6500
rect 14202 6556 14266 6560
rect 14202 6500 14206 6556
rect 14206 6500 14262 6556
rect 14262 6500 14266 6556
rect 14202 6496 14266 6500
rect 17062 6556 17126 6560
rect 17062 6500 17066 6556
rect 17066 6500 17122 6556
rect 17122 6500 17126 6556
rect 17062 6496 17126 6500
rect 17142 6556 17206 6560
rect 17142 6500 17146 6556
rect 17146 6500 17202 6556
rect 17202 6500 17206 6556
rect 17142 6496 17206 6500
rect 17222 6556 17286 6560
rect 17222 6500 17226 6556
rect 17226 6500 17282 6556
rect 17282 6500 17286 6556
rect 17222 6496 17286 6500
rect 17302 6556 17366 6560
rect 17302 6500 17306 6556
rect 17306 6500 17362 6556
rect 17362 6500 17366 6556
rect 17302 6496 17366 6500
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 3272 6012 3336 6016
rect 3272 5956 3276 6012
rect 3276 5956 3332 6012
rect 3332 5956 3336 6012
rect 3272 5952 3336 5956
rect 3352 6012 3416 6016
rect 3352 5956 3356 6012
rect 3356 5956 3412 6012
rect 3412 5956 3416 6012
rect 3352 5952 3416 5956
rect 6212 6012 6276 6016
rect 6212 5956 6216 6012
rect 6216 5956 6272 6012
rect 6272 5956 6276 6012
rect 6212 5952 6276 5956
rect 6292 6012 6356 6016
rect 6292 5956 6296 6012
rect 6296 5956 6352 6012
rect 6352 5956 6356 6012
rect 6292 5952 6356 5956
rect 6372 6012 6436 6016
rect 6372 5956 6376 6012
rect 6376 5956 6432 6012
rect 6432 5956 6436 6012
rect 6372 5952 6436 5956
rect 6452 6012 6516 6016
rect 6452 5956 6456 6012
rect 6456 5956 6512 6012
rect 6512 5956 6516 6012
rect 6452 5952 6516 5956
rect 9312 6012 9376 6016
rect 9312 5956 9316 6012
rect 9316 5956 9372 6012
rect 9372 5956 9376 6012
rect 9312 5952 9376 5956
rect 9392 6012 9456 6016
rect 9392 5956 9396 6012
rect 9396 5956 9452 6012
rect 9452 5956 9456 6012
rect 9392 5952 9456 5956
rect 9472 6012 9536 6016
rect 9472 5956 9476 6012
rect 9476 5956 9532 6012
rect 9532 5956 9536 6012
rect 9472 5952 9536 5956
rect 9552 6012 9616 6016
rect 9552 5956 9556 6012
rect 9556 5956 9612 6012
rect 9612 5956 9616 6012
rect 9552 5952 9616 5956
rect 12412 6012 12476 6016
rect 12412 5956 12416 6012
rect 12416 5956 12472 6012
rect 12472 5956 12476 6012
rect 12412 5952 12476 5956
rect 12492 6012 12556 6016
rect 12492 5956 12496 6012
rect 12496 5956 12552 6012
rect 12552 5956 12556 6012
rect 12492 5952 12556 5956
rect 12572 6012 12636 6016
rect 12572 5956 12576 6012
rect 12576 5956 12632 6012
rect 12632 5956 12636 6012
rect 12572 5952 12636 5956
rect 12652 6012 12716 6016
rect 12652 5956 12656 6012
rect 12656 5956 12712 6012
rect 12712 5956 12716 6012
rect 12652 5952 12716 5956
rect 15512 6012 15576 6016
rect 15512 5956 15516 6012
rect 15516 5956 15572 6012
rect 15572 5956 15576 6012
rect 15512 5952 15576 5956
rect 15592 6012 15656 6016
rect 15592 5956 15596 6012
rect 15596 5956 15652 6012
rect 15652 5956 15656 6012
rect 15592 5952 15656 5956
rect 15672 6012 15736 6016
rect 15672 5956 15676 6012
rect 15676 5956 15732 6012
rect 15732 5956 15736 6012
rect 15672 5952 15736 5956
rect 15752 6012 15816 6016
rect 15752 5956 15756 6012
rect 15756 5956 15812 6012
rect 15812 5956 15816 6012
rect 15752 5952 15816 5956
rect 4662 5468 4726 5472
rect 4662 5412 4666 5468
rect 4666 5412 4722 5468
rect 4722 5412 4726 5468
rect 4662 5408 4726 5412
rect 4742 5468 4806 5472
rect 4742 5412 4746 5468
rect 4746 5412 4802 5468
rect 4802 5412 4806 5468
rect 4742 5408 4806 5412
rect 4822 5468 4886 5472
rect 4822 5412 4826 5468
rect 4826 5412 4882 5468
rect 4882 5412 4886 5468
rect 4822 5408 4886 5412
rect 4902 5468 4966 5472
rect 4902 5412 4906 5468
rect 4906 5412 4962 5468
rect 4962 5412 4966 5468
rect 4902 5408 4966 5412
rect 7762 5468 7826 5472
rect 7762 5412 7766 5468
rect 7766 5412 7822 5468
rect 7822 5412 7826 5468
rect 7762 5408 7826 5412
rect 7842 5468 7906 5472
rect 7842 5412 7846 5468
rect 7846 5412 7902 5468
rect 7902 5412 7906 5468
rect 7842 5408 7906 5412
rect 7922 5468 7986 5472
rect 7922 5412 7926 5468
rect 7926 5412 7982 5468
rect 7982 5412 7986 5468
rect 7922 5408 7986 5412
rect 8002 5468 8066 5472
rect 8002 5412 8006 5468
rect 8006 5412 8062 5468
rect 8062 5412 8066 5468
rect 8002 5408 8066 5412
rect 10862 5468 10926 5472
rect 10862 5412 10866 5468
rect 10866 5412 10922 5468
rect 10922 5412 10926 5468
rect 10862 5408 10926 5412
rect 10942 5468 11006 5472
rect 10942 5412 10946 5468
rect 10946 5412 11002 5468
rect 11002 5412 11006 5468
rect 10942 5408 11006 5412
rect 11022 5468 11086 5472
rect 11022 5412 11026 5468
rect 11026 5412 11082 5468
rect 11082 5412 11086 5468
rect 11022 5408 11086 5412
rect 11102 5468 11166 5472
rect 11102 5412 11106 5468
rect 11106 5412 11162 5468
rect 11162 5412 11166 5468
rect 11102 5408 11166 5412
rect 13962 5468 14026 5472
rect 13962 5412 13966 5468
rect 13966 5412 14022 5468
rect 14022 5412 14026 5468
rect 13962 5408 14026 5412
rect 14042 5468 14106 5472
rect 14042 5412 14046 5468
rect 14046 5412 14102 5468
rect 14102 5412 14106 5468
rect 14042 5408 14106 5412
rect 14122 5468 14186 5472
rect 14122 5412 14126 5468
rect 14126 5412 14182 5468
rect 14182 5412 14186 5468
rect 14122 5408 14186 5412
rect 14202 5468 14266 5472
rect 14202 5412 14206 5468
rect 14206 5412 14262 5468
rect 14262 5412 14266 5468
rect 14202 5408 14266 5412
rect 17062 5468 17126 5472
rect 17062 5412 17066 5468
rect 17066 5412 17122 5468
rect 17122 5412 17126 5468
rect 17062 5408 17126 5412
rect 17142 5468 17206 5472
rect 17142 5412 17146 5468
rect 17146 5412 17202 5468
rect 17202 5412 17206 5468
rect 17142 5408 17206 5412
rect 17222 5468 17286 5472
rect 17222 5412 17226 5468
rect 17226 5412 17282 5468
rect 17282 5412 17286 5468
rect 17222 5408 17286 5412
rect 17302 5468 17366 5472
rect 17302 5412 17306 5468
rect 17306 5412 17362 5468
rect 17362 5412 17366 5468
rect 17302 5408 17366 5412
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 3272 4924 3336 4928
rect 3272 4868 3276 4924
rect 3276 4868 3332 4924
rect 3332 4868 3336 4924
rect 3272 4864 3336 4868
rect 3352 4924 3416 4928
rect 3352 4868 3356 4924
rect 3356 4868 3412 4924
rect 3412 4868 3416 4924
rect 3352 4864 3416 4868
rect 6212 4924 6276 4928
rect 6212 4868 6216 4924
rect 6216 4868 6272 4924
rect 6272 4868 6276 4924
rect 6212 4864 6276 4868
rect 6292 4924 6356 4928
rect 6292 4868 6296 4924
rect 6296 4868 6352 4924
rect 6352 4868 6356 4924
rect 6292 4864 6356 4868
rect 6372 4924 6436 4928
rect 6372 4868 6376 4924
rect 6376 4868 6432 4924
rect 6432 4868 6436 4924
rect 6372 4864 6436 4868
rect 6452 4924 6516 4928
rect 6452 4868 6456 4924
rect 6456 4868 6512 4924
rect 6512 4868 6516 4924
rect 6452 4864 6516 4868
rect 9312 4924 9376 4928
rect 9312 4868 9316 4924
rect 9316 4868 9372 4924
rect 9372 4868 9376 4924
rect 9312 4864 9376 4868
rect 9392 4924 9456 4928
rect 9392 4868 9396 4924
rect 9396 4868 9452 4924
rect 9452 4868 9456 4924
rect 9392 4864 9456 4868
rect 9472 4924 9536 4928
rect 9472 4868 9476 4924
rect 9476 4868 9532 4924
rect 9532 4868 9536 4924
rect 9472 4864 9536 4868
rect 9552 4924 9616 4928
rect 9552 4868 9556 4924
rect 9556 4868 9612 4924
rect 9612 4868 9616 4924
rect 9552 4864 9616 4868
rect 12412 4924 12476 4928
rect 12412 4868 12416 4924
rect 12416 4868 12472 4924
rect 12472 4868 12476 4924
rect 12412 4864 12476 4868
rect 12492 4924 12556 4928
rect 12492 4868 12496 4924
rect 12496 4868 12552 4924
rect 12552 4868 12556 4924
rect 12492 4864 12556 4868
rect 12572 4924 12636 4928
rect 12572 4868 12576 4924
rect 12576 4868 12632 4924
rect 12632 4868 12636 4924
rect 12572 4864 12636 4868
rect 12652 4924 12716 4928
rect 12652 4868 12656 4924
rect 12656 4868 12712 4924
rect 12712 4868 12716 4924
rect 12652 4864 12716 4868
rect 15512 4924 15576 4928
rect 15512 4868 15516 4924
rect 15516 4868 15572 4924
rect 15572 4868 15576 4924
rect 15512 4864 15576 4868
rect 15592 4924 15656 4928
rect 15592 4868 15596 4924
rect 15596 4868 15652 4924
rect 15652 4868 15656 4924
rect 15592 4864 15656 4868
rect 15672 4924 15736 4928
rect 15672 4868 15676 4924
rect 15676 4868 15732 4924
rect 15732 4868 15736 4924
rect 15672 4864 15736 4868
rect 15752 4924 15816 4928
rect 15752 4868 15756 4924
rect 15756 4868 15812 4924
rect 15812 4868 15816 4924
rect 15752 4864 15816 4868
rect 4662 4380 4726 4384
rect 4662 4324 4666 4380
rect 4666 4324 4722 4380
rect 4722 4324 4726 4380
rect 4662 4320 4726 4324
rect 4742 4380 4806 4384
rect 4742 4324 4746 4380
rect 4746 4324 4802 4380
rect 4802 4324 4806 4380
rect 4742 4320 4806 4324
rect 4822 4380 4886 4384
rect 4822 4324 4826 4380
rect 4826 4324 4882 4380
rect 4882 4324 4886 4380
rect 4822 4320 4886 4324
rect 4902 4380 4966 4384
rect 4902 4324 4906 4380
rect 4906 4324 4962 4380
rect 4962 4324 4966 4380
rect 4902 4320 4966 4324
rect 7762 4380 7826 4384
rect 7762 4324 7766 4380
rect 7766 4324 7822 4380
rect 7822 4324 7826 4380
rect 7762 4320 7826 4324
rect 7842 4380 7906 4384
rect 7842 4324 7846 4380
rect 7846 4324 7902 4380
rect 7902 4324 7906 4380
rect 7842 4320 7906 4324
rect 7922 4380 7986 4384
rect 7922 4324 7926 4380
rect 7926 4324 7982 4380
rect 7982 4324 7986 4380
rect 7922 4320 7986 4324
rect 8002 4380 8066 4384
rect 8002 4324 8006 4380
rect 8006 4324 8062 4380
rect 8062 4324 8066 4380
rect 8002 4320 8066 4324
rect 10862 4380 10926 4384
rect 10862 4324 10866 4380
rect 10866 4324 10922 4380
rect 10922 4324 10926 4380
rect 10862 4320 10926 4324
rect 10942 4380 11006 4384
rect 10942 4324 10946 4380
rect 10946 4324 11002 4380
rect 11002 4324 11006 4380
rect 10942 4320 11006 4324
rect 11022 4380 11086 4384
rect 11022 4324 11026 4380
rect 11026 4324 11082 4380
rect 11082 4324 11086 4380
rect 11022 4320 11086 4324
rect 11102 4380 11166 4384
rect 11102 4324 11106 4380
rect 11106 4324 11162 4380
rect 11162 4324 11166 4380
rect 11102 4320 11166 4324
rect 13962 4380 14026 4384
rect 13962 4324 13966 4380
rect 13966 4324 14022 4380
rect 14022 4324 14026 4380
rect 13962 4320 14026 4324
rect 14042 4380 14106 4384
rect 14042 4324 14046 4380
rect 14046 4324 14102 4380
rect 14102 4324 14106 4380
rect 14042 4320 14106 4324
rect 14122 4380 14186 4384
rect 14122 4324 14126 4380
rect 14126 4324 14182 4380
rect 14182 4324 14186 4380
rect 14122 4320 14186 4324
rect 14202 4380 14266 4384
rect 14202 4324 14206 4380
rect 14206 4324 14262 4380
rect 14262 4324 14266 4380
rect 14202 4320 14266 4324
rect 17062 4380 17126 4384
rect 17062 4324 17066 4380
rect 17066 4324 17122 4380
rect 17122 4324 17126 4380
rect 17062 4320 17126 4324
rect 17142 4380 17206 4384
rect 17142 4324 17146 4380
rect 17146 4324 17202 4380
rect 17202 4324 17206 4380
rect 17142 4320 17206 4324
rect 17222 4380 17286 4384
rect 17222 4324 17226 4380
rect 17226 4324 17282 4380
rect 17282 4324 17286 4380
rect 17222 4320 17286 4324
rect 17302 4380 17366 4384
rect 17302 4324 17306 4380
rect 17306 4324 17362 4380
rect 17362 4324 17366 4380
rect 17302 4320 17366 4324
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 3272 3836 3336 3840
rect 3272 3780 3276 3836
rect 3276 3780 3332 3836
rect 3332 3780 3336 3836
rect 3272 3776 3336 3780
rect 3352 3836 3416 3840
rect 3352 3780 3356 3836
rect 3356 3780 3412 3836
rect 3412 3780 3416 3836
rect 3352 3776 3416 3780
rect 6212 3836 6276 3840
rect 6212 3780 6216 3836
rect 6216 3780 6272 3836
rect 6272 3780 6276 3836
rect 6212 3776 6276 3780
rect 6292 3836 6356 3840
rect 6292 3780 6296 3836
rect 6296 3780 6352 3836
rect 6352 3780 6356 3836
rect 6292 3776 6356 3780
rect 6372 3836 6436 3840
rect 6372 3780 6376 3836
rect 6376 3780 6432 3836
rect 6432 3780 6436 3836
rect 6372 3776 6436 3780
rect 6452 3836 6516 3840
rect 6452 3780 6456 3836
rect 6456 3780 6512 3836
rect 6512 3780 6516 3836
rect 6452 3776 6516 3780
rect 9312 3836 9376 3840
rect 9312 3780 9316 3836
rect 9316 3780 9372 3836
rect 9372 3780 9376 3836
rect 9312 3776 9376 3780
rect 9392 3836 9456 3840
rect 9392 3780 9396 3836
rect 9396 3780 9452 3836
rect 9452 3780 9456 3836
rect 9392 3776 9456 3780
rect 9472 3836 9536 3840
rect 9472 3780 9476 3836
rect 9476 3780 9532 3836
rect 9532 3780 9536 3836
rect 9472 3776 9536 3780
rect 9552 3836 9616 3840
rect 9552 3780 9556 3836
rect 9556 3780 9612 3836
rect 9612 3780 9616 3836
rect 9552 3776 9616 3780
rect 12412 3836 12476 3840
rect 12412 3780 12416 3836
rect 12416 3780 12472 3836
rect 12472 3780 12476 3836
rect 12412 3776 12476 3780
rect 12492 3836 12556 3840
rect 12492 3780 12496 3836
rect 12496 3780 12552 3836
rect 12552 3780 12556 3836
rect 12492 3776 12556 3780
rect 12572 3836 12636 3840
rect 12572 3780 12576 3836
rect 12576 3780 12632 3836
rect 12632 3780 12636 3836
rect 12572 3776 12636 3780
rect 12652 3836 12716 3840
rect 12652 3780 12656 3836
rect 12656 3780 12712 3836
rect 12712 3780 12716 3836
rect 12652 3776 12716 3780
rect 15512 3836 15576 3840
rect 15512 3780 15516 3836
rect 15516 3780 15572 3836
rect 15572 3780 15576 3836
rect 15512 3776 15576 3780
rect 15592 3836 15656 3840
rect 15592 3780 15596 3836
rect 15596 3780 15652 3836
rect 15652 3780 15656 3836
rect 15592 3776 15656 3780
rect 15672 3836 15736 3840
rect 15672 3780 15676 3836
rect 15676 3780 15732 3836
rect 15732 3780 15736 3836
rect 15672 3776 15736 3780
rect 15752 3836 15816 3840
rect 15752 3780 15756 3836
rect 15756 3780 15812 3836
rect 15812 3780 15816 3836
rect 15752 3776 15816 3780
rect 4662 3292 4726 3296
rect 4662 3236 4666 3292
rect 4666 3236 4722 3292
rect 4722 3236 4726 3292
rect 4662 3232 4726 3236
rect 4742 3292 4806 3296
rect 4742 3236 4746 3292
rect 4746 3236 4802 3292
rect 4802 3236 4806 3292
rect 4742 3232 4806 3236
rect 4822 3292 4886 3296
rect 4822 3236 4826 3292
rect 4826 3236 4882 3292
rect 4882 3236 4886 3292
rect 4822 3232 4886 3236
rect 4902 3292 4966 3296
rect 4902 3236 4906 3292
rect 4906 3236 4962 3292
rect 4962 3236 4966 3292
rect 4902 3232 4966 3236
rect 7762 3292 7826 3296
rect 7762 3236 7766 3292
rect 7766 3236 7822 3292
rect 7822 3236 7826 3292
rect 7762 3232 7826 3236
rect 7842 3292 7906 3296
rect 7842 3236 7846 3292
rect 7846 3236 7902 3292
rect 7902 3236 7906 3292
rect 7842 3232 7906 3236
rect 7922 3292 7986 3296
rect 7922 3236 7926 3292
rect 7926 3236 7982 3292
rect 7982 3236 7986 3292
rect 7922 3232 7986 3236
rect 8002 3292 8066 3296
rect 8002 3236 8006 3292
rect 8006 3236 8062 3292
rect 8062 3236 8066 3292
rect 8002 3232 8066 3236
rect 10862 3292 10926 3296
rect 10862 3236 10866 3292
rect 10866 3236 10922 3292
rect 10922 3236 10926 3292
rect 10862 3232 10926 3236
rect 10942 3292 11006 3296
rect 10942 3236 10946 3292
rect 10946 3236 11002 3292
rect 11002 3236 11006 3292
rect 10942 3232 11006 3236
rect 11022 3292 11086 3296
rect 11022 3236 11026 3292
rect 11026 3236 11082 3292
rect 11082 3236 11086 3292
rect 11022 3232 11086 3236
rect 11102 3292 11166 3296
rect 11102 3236 11106 3292
rect 11106 3236 11162 3292
rect 11162 3236 11166 3292
rect 11102 3232 11166 3236
rect 13962 3292 14026 3296
rect 13962 3236 13966 3292
rect 13966 3236 14022 3292
rect 14022 3236 14026 3292
rect 13962 3232 14026 3236
rect 14042 3292 14106 3296
rect 14042 3236 14046 3292
rect 14046 3236 14102 3292
rect 14102 3236 14106 3292
rect 14042 3232 14106 3236
rect 14122 3292 14186 3296
rect 14122 3236 14126 3292
rect 14126 3236 14182 3292
rect 14182 3236 14186 3292
rect 14122 3232 14186 3236
rect 14202 3292 14266 3296
rect 14202 3236 14206 3292
rect 14206 3236 14262 3292
rect 14262 3236 14266 3292
rect 14202 3232 14266 3236
rect 17062 3292 17126 3296
rect 17062 3236 17066 3292
rect 17066 3236 17122 3292
rect 17122 3236 17126 3292
rect 17062 3232 17126 3236
rect 17142 3292 17206 3296
rect 17142 3236 17146 3292
rect 17146 3236 17202 3292
rect 17202 3236 17206 3292
rect 17142 3232 17206 3236
rect 17222 3292 17286 3296
rect 17222 3236 17226 3292
rect 17226 3236 17282 3292
rect 17282 3236 17286 3292
rect 17222 3232 17286 3236
rect 17302 3292 17366 3296
rect 17302 3236 17306 3292
rect 17306 3236 17362 3292
rect 17362 3236 17366 3292
rect 17302 3232 17366 3236
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 3272 2748 3336 2752
rect 3272 2692 3276 2748
rect 3276 2692 3332 2748
rect 3332 2692 3336 2748
rect 3272 2688 3336 2692
rect 3352 2748 3416 2752
rect 3352 2692 3356 2748
rect 3356 2692 3412 2748
rect 3412 2692 3416 2748
rect 3352 2688 3416 2692
rect 6212 2748 6276 2752
rect 6212 2692 6216 2748
rect 6216 2692 6272 2748
rect 6272 2692 6276 2748
rect 6212 2688 6276 2692
rect 6292 2748 6356 2752
rect 6292 2692 6296 2748
rect 6296 2692 6352 2748
rect 6352 2692 6356 2748
rect 6292 2688 6356 2692
rect 6372 2748 6436 2752
rect 6372 2692 6376 2748
rect 6376 2692 6432 2748
rect 6432 2692 6436 2748
rect 6372 2688 6436 2692
rect 6452 2748 6516 2752
rect 6452 2692 6456 2748
rect 6456 2692 6512 2748
rect 6512 2692 6516 2748
rect 6452 2688 6516 2692
rect 9312 2748 9376 2752
rect 9312 2692 9316 2748
rect 9316 2692 9372 2748
rect 9372 2692 9376 2748
rect 9312 2688 9376 2692
rect 9392 2748 9456 2752
rect 9392 2692 9396 2748
rect 9396 2692 9452 2748
rect 9452 2692 9456 2748
rect 9392 2688 9456 2692
rect 9472 2748 9536 2752
rect 9472 2692 9476 2748
rect 9476 2692 9532 2748
rect 9532 2692 9536 2748
rect 9472 2688 9536 2692
rect 9552 2748 9616 2752
rect 9552 2692 9556 2748
rect 9556 2692 9612 2748
rect 9612 2692 9616 2748
rect 9552 2688 9616 2692
rect 12412 2748 12476 2752
rect 12412 2692 12416 2748
rect 12416 2692 12472 2748
rect 12472 2692 12476 2748
rect 12412 2688 12476 2692
rect 12492 2748 12556 2752
rect 12492 2692 12496 2748
rect 12496 2692 12552 2748
rect 12552 2692 12556 2748
rect 12492 2688 12556 2692
rect 12572 2748 12636 2752
rect 12572 2692 12576 2748
rect 12576 2692 12632 2748
rect 12632 2692 12636 2748
rect 12572 2688 12636 2692
rect 12652 2748 12716 2752
rect 12652 2692 12656 2748
rect 12656 2692 12712 2748
rect 12712 2692 12716 2748
rect 12652 2688 12716 2692
rect 15512 2748 15576 2752
rect 15512 2692 15516 2748
rect 15516 2692 15572 2748
rect 15572 2692 15576 2748
rect 15512 2688 15576 2692
rect 15592 2748 15656 2752
rect 15592 2692 15596 2748
rect 15596 2692 15652 2748
rect 15652 2692 15656 2748
rect 15592 2688 15656 2692
rect 15672 2748 15736 2752
rect 15672 2692 15676 2748
rect 15676 2692 15732 2748
rect 15732 2692 15736 2748
rect 15672 2688 15736 2692
rect 15752 2748 15816 2752
rect 15752 2692 15756 2748
rect 15756 2692 15812 2748
rect 15812 2692 15816 2748
rect 15752 2688 15816 2692
rect 4662 2204 4726 2208
rect 4662 2148 4666 2204
rect 4666 2148 4722 2204
rect 4722 2148 4726 2204
rect 4662 2144 4726 2148
rect 4742 2204 4806 2208
rect 4742 2148 4746 2204
rect 4746 2148 4802 2204
rect 4802 2148 4806 2204
rect 4742 2144 4806 2148
rect 4822 2204 4886 2208
rect 4822 2148 4826 2204
rect 4826 2148 4882 2204
rect 4882 2148 4886 2204
rect 4822 2144 4886 2148
rect 4902 2204 4966 2208
rect 4902 2148 4906 2204
rect 4906 2148 4962 2204
rect 4962 2148 4966 2204
rect 4902 2144 4966 2148
rect 7762 2204 7826 2208
rect 7762 2148 7766 2204
rect 7766 2148 7822 2204
rect 7822 2148 7826 2204
rect 7762 2144 7826 2148
rect 7842 2204 7906 2208
rect 7842 2148 7846 2204
rect 7846 2148 7902 2204
rect 7902 2148 7906 2204
rect 7842 2144 7906 2148
rect 7922 2204 7986 2208
rect 7922 2148 7926 2204
rect 7926 2148 7982 2204
rect 7982 2148 7986 2204
rect 7922 2144 7986 2148
rect 8002 2204 8066 2208
rect 8002 2148 8006 2204
rect 8006 2148 8062 2204
rect 8062 2148 8066 2204
rect 8002 2144 8066 2148
rect 10862 2204 10926 2208
rect 10862 2148 10866 2204
rect 10866 2148 10922 2204
rect 10922 2148 10926 2204
rect 10862 2144 10926 2148
rect 10942 2204 11006 2208
rect 10942 2148 10946 2204
rect 10946 2148 11002 2204
rect 11002 2148 11006 2204
rect 10942 2144 11006 2148
rect 11022 2204 11086 2208
rect 11022 2148 11026 2204
rect 11026 2148 11082 2204
rect 11082 2148 11086 2204
rect 11022 2144 11086 2148
rect 11102 2204 11166 2208
rect 11102 2148 11106 2204
rect 11106 2148 11162 2204
rect 11162 2148 11166 2204
rect 11102 2144 11166 2148
rect 13962 2204 14026 2208
rect 13962 2148 13966 2204
rect 13966 2148 14022 2204
rect 14022 2148 14026 2204
rect 13962 2144 14026 2148
rect 14042 2204 14106 2208
rect 14042 2148 14046 2204
rect 14046 2148 14102 2204
rect 14102 2148 14106 2204
rect 14042 2144 14106 2148
rect 14122 2204 14186 2208
rect 14122 2148 14126 2204
rect 14126 2148 14182 2204
rect 14182 2148 14186 2204
rect 14122 2144 14186 2148
rect 14202 2204 14266 2208
rect 14202 2148 14206 2204
rect 14206 2148 14262 2204
rect 14262 2148 14266 2204
rect 14202 2144 14266 2148
rect 17062 2204 17126 2208
rect 17062 2148 17066 2204
rect 17066 2148 17122 2204
rect 17122 2148 17126 2204
rect 17062 2144 17126 2148
rect 17142 2204 17206 2208
rect 17142 2148 17146 2204
rect 17146 2148 17202 2204
rect 17202 2148 17206 2204
rect 17142 2144 17206 2148
rect 17222 2204 17286 2208
rect 17222 2148 17226 2204
rect 17226 2148 17282 2204
rect 17282 2148 17286 2204
rect 17222 2144 17286 2148
rect 17302 2204 17366 2208
rect 17302 2148 17306 2204
rect 17306 2148 17362 2204
rect 17362 2148 17366 2204
rect 17302 2144 17366 2148
rect 3112 1660 3176 1664
rect 3112 1604 3116 1660
rect 3116 1604 3172 1660
rect 3172 1604 3176 1660
rect 3112 1600 3176 1604
rect 3192 1660 3256 1664
rect 3192 1604 3196 1660
rect 3196 1604 3252 1660
rect 3252 1604 3256 1660
rect 3192 1600 3256 1604
rect 3272 1660 3336 1664
rect 3272 1604 3276 1660
rect 3276 1604 3332 1660
rect 3332 1604 3336 1660
rect 3272 1600 3336 1604
rect 3352 1660 3416 1664
rect 3352 1604 3356 1660
rect 3356 1604 3412 1660
rect 3412 1604 3416 1660
rect 3352 1600 3416 1604
rect 6212 1660 6276 1664
rect 6212 1604 6216 1660
rect 6216 1604 6272 1660
rect 6272 1604 6276 1660
rect 6212 1600 6276 1604
rect 6292 1660 6356 1664
rect 6292 1604 6296 1660
rect 6296 1604 6352 1660
rect 6352 1604 6356 1660
rect 6292 1600 6356 1604
rect 6372 1660 6436 1664
rect 6372 1604 6376 1660
rect 6376 1604 6432 1660
rect 6432 1604 6436 1660
rect 6372 1600 6436 1604
rect 6452 1660 6516 1664
rect 6452 1604 6456 1660
rect 6456 1604 6512 1660
rect 6512 1604 6516 1660
rect 6452 1600 6516 1604
rect 9312 1660 9376 1664
rect 9312 1604 9316 1660
rect 9316 1604 9372 1660
rect 9372 1604 9376 1660
rect 9312 1600 9376 1604
rect 9392 1660 9456 1664
rect 9392 1604 9396 1660
rect 9396 1604 9452 1660
rect 9452 1604 9456 1660
rect 9392 1600 9456 1604
rect 9472 1660 9536 1664
rect 9472 1604 9476 1660
rect 9476 1604 9532 1660
rect 9532 1604 9536 1660
rect 9472 1600 9536 1604
rect 9552 1660 9616 1664
rect 9552 1604 9556 1660
rect 9556 1604 9612 1660
rect 9612 1604 9616 1660
rect 9552 1600 9616 1604
rect 12412 1660 12476 1664
rect 12412 1604 12416 1660
rect 12416 1604 12472 1660
rect 12472 1604 12476 1660
rect 12412 1600 12476 1604
rect 12492 1660 12556 1664
rect 12492 1604 12496 1660
rect 12496 1604 12552 1660
rect 12552 1604 12556 1660
rect 12492 1600 12556 1604
rect 12572 1660 12636 1664
rect 12572 1604 12576 1660
rect 12576 1604 12632 1660
rect 12632 1604 12636 1660
rect 12572 1600 12636 1604
rect 12652 1660 12716 1664
rect 12652 1604 12656 1660
rect 12656 1604 12712 1660
rect 12712 1604 12716 1660
rect 12652 1600 12716 1604
rect 15512 1660 15576 1664
rect 15512 1604 15516 1660
rect 15516 1604 15572 1660
rect 15572 1604 15576 1660
rect 15512 1600 15576 1604
rect 15592 1660 15656 1664
rect 15592 1604 15596 1660
rect 15596 1604 15652 1660
rect 15652 1604 15656 1660
rect 15592 1600 15656 1604
rect 15672 1660 15736 1664
rect 15672 1604 15676 1660
rect 15676 1604 15732 1660
rect 15732 1604 15736 1660
rect 15672 1600 15736 1604
rect 15752 1660 15816 1664
rect 15752 1604 15756 1660
rect 15756 1604 15812 1660
rect 15812 1604 15816 1660
rect 15752 1600 15816 1604
rect 4662 1116 4726 1120
rect 4662 1060 4666 1116
rect 4666 1060 4722 1116
rect 4722 1060 4726 1116
rect 4662 1056 4726 1060
rect 4742 1116 4806 1120
rect 4742 1060 4746 1116
rect 4746 1060 4802 1116
rect 4802 1060 4806 1116
rect 4742 1056 4806 1060
rect 4822 1116 4886 1120
rect 4822 1060 4826 1116
rect 4826 1060 4882 1116
rect 4882 1060 4886 1116
rect 4822 1056 4886 1060
rect 4902 1116 4966 1120
rect 4902 1060 4906 1116
rect 4906 1060 4962 1116
rect 4962 1060 4966 1116
rect 4902 1056 4966 1060
rect 7762 1116 7826 1120
rect 7762 1060 7766 1116
rect 7766 1060 7822 1116
rect 7822 1060 7826 1116
rect 7762 1056 7826 1060
rect 7842 1116 7906 1120
rect 7842 1060 7846 1116
rect 7846 1060 7902 1116
rect 7902 1060 7906 1116
rect 7842 1056 7906 1060
rect 7922 1116 7986 1120
rect 7922 1060 7926 1116
rect 7926 1060 7982 1116
rect 7982 1060 7986 1116
rect 7922 1056 7986 1060
rect 8002 1116 8066 1120
rect 8002 1060 8006 1116
rect 8006 1060 8062 1116
rect 8062 1060 8066 1116
rect 8002 1056 8066 1060
rect 10862 1116 10926 1120
rect 10862 1060 10866 1116
rect 10866 1060 10922 1116
rect 10922 1060 10926 1116
rect 10862 1056 10926 1060
rect 10942 1116 11006 1120
rect 10942 1060 10946 1116
rect 10946 1060 11002 1116
rect 11002 1060 11006 1116
rect 10942 1056 11006 1060
rect 11022 1116 11086 1120
rect 11022 1060 11026 1116
rect 11026 1060 11082 1116
rect 11082 1060 11086 1116
rect 11022 1056 11086 1060
rect 11102 1116 11166 1120
rect 11102 1060 11106 1116
rect 11106 1060 11162 1116
rect 11162 1060 11166 1116
rect 11102 1056 11166 1060
rect 13962 1116 14026 1120
rect 13962 1060 13966 1116
rect 13966 1060 14022 1116
rect 14022 1060 14026 1116
rect 13962 1056 14026 1060
rect 14042 1116 14106 1120
rect 14042 1060 14046 1116
rect 14046 1060 14102 1116
rect 14102 1060 14106 1116
rect 14042 1056 14106 1060
rect 14122 1116 14186 1120
rect 14122 1060 14126 1116
rect 14126 1060 14182 1116
rect 14182 1060 14186 1116
rect 14122 1056 14186 1060
rect 14202 1116 14266 1120
rect 14202 1060 14206 1116
rect 14206 1060 14262 1116
rect 14262 1060 14266 1116
rect 14202 1056 14266 1060
rect 17062 1116 17126 1120
rect 17062 1060 17066 1116
rect 17066 1060 17122 1116
rect 17122 1060 17126 1116
rect 17062 1056 17126 1060
rect 17142 1116 17206 1120
rect 17142 1060 17146 1116
rect 17146 1060 17202 1116
rect 17202 1060 17206 1116
rect 17142 1056 17206 1060
rect 17222 1116 17286 1120
rect 17222 1060 17226 1116
rect 17226 1060 17282 1116
rect 17282 1060 17286 1116
rect 17222 1056 17286 1060
rect 17302 1116 17366 1120
rect 17302 1060 17306 1116
rect 17306 1060 17362 1116
rect 17362 1060 17366 1116
rect 17302 1056 17366 1060
rect 3112 572 3176 576
rect 3112 516 3116 572
rect 3116 516 3172 572
rect 3172 516 3176 572
rect 3112 512 3176 516
rect 3192 572 3256 576
rect 3192 516 3196 572
rect 3196 516 3252 572
rect 3252 516 3256 572
rect 3192 512 3256 516
rect 3272 572 3336 576
rect 3272 516 3276 572
rect 3276 516 3332 572
rect 3332 516 3336 572
rect 3272 512 3336 516
rect 3352 572 3416 576
rect 3352 516 3356 572
rect 3356 516 3412 572
rect 3412 516 3416 572
rect 3352 512 3416 516
rect 6212 572 6276 576
rect 6212 516 6216 572
rect 6216 516 6272 572
rect 6272 516 6276 572
rect 6212 512 6276 516
rect 6292 572 6356 576
rect 6292 516 6296 572
rect 6296 516 6352 572
rect 6352 516 6356 572
rect 6292 512 6356 516
rect 6372 572 6436 576
rect 6372 516 6376 572
rect 6376 516 6432 572
rect 6432 516 6436 572
rect 6372 512 6436 516
rect 6452 572 6516 576
rect 6452 516 6456 572
rect 6456 516 6512 572
rect 6512 516 6516 572
rect 6452 512 6516 516
rect 9312 572 9376 576
rect 9312 516 9316 572
rect 9316 516 9372 572
rect 9372 516 9376 572
rect 9312 512 9376 516
rect 9392 572 9456 576
rect 9392 516 9396 572
rect 9396 516 9452 572
rect 9452 516 9456 572
rect 9392 512 9456 516
rect 9472 572 9536 576
rect 9472 516 9476 572
rect 9476 516 9532 572
rect 9532 516 9536 572
rect 9472 512 9536 516
rect 9552 572 9616 576
rect 9552 516 9556 572
rect 9556 516 9612 572
rect 9612 516 9616 572
rect 9552 512 9616 516
rect 12412 572 12476 576
rect 12412 516 12416 572
rect 12416 516 12472 572
rect 12472 516 12476 572
rect 12412 512 12476 516
rect 12492 572 12556 576
rect 12492 516 12496 572
rect 12496 516 12552 572
rect 12552 516 12556 572
rect 12492 512 12556 516
rect 12572 572 12636 576
rect 12572 516 12576 572
rect 12576 516 12632 572
rect 12632 516 12636 572
rect 12572 512 12636 516
rect 12652 572 12716 576
rect 12652 516 12656 572
rect 12656 516 12712 572
rect 12712 516 12716 572
rect 12652 512 12716 516
rect 15512 572 15576 576
rect 15512 516 15516 572
rect 15516 516 15572 572
rect 15572 516 15576 572
rect 15512 512 15576 516
rect 15592 572 15656 576
rect 15592 516 15596 572
rect 15596 516 15652 572
rect 15652 516 15656 572
rect 15592 512 15656 516
rect 15672 572 15736 576
rect 15672 516 15676 572
rect 15676 516 15732 572
rect 15732 516 15736 572
rect 15672 512 15736 516
rect 15752 572 15816 576
rect 15752 516 15756 572
rect 15756 516 15812 572
rect 15812 516 15816 572
rect 15752 512 15816 516
rect 4662 28 4726 32
rect 4662 -28 4666 28
rect 4666 -28 4722 28
rect 4722 -28 4726 28
rect 4662 -32 4726 -28
rect 4742 28 4806 32
rect 4742 -28 4746 28
rect 4746 -28 4802 28
rect 4802 -28 4806 28
rect 4742 -32 4806 -28
rect 4822 28 4886 32
rect 4822 -28 4826 28
rect 4826 -28 4882 28
rect 4882 -28 4886 28
rect 4822 -32 4886 -28
rect 4902 28 4966 32
rect 4902 -28 4906 28
rect 4906 -28 4962 28
rect 4962 -28 4966 28
rect 4902 -32 4966 -28
rect 7762 28 7826 32
rect 7762 -28 7766 28
rect 7766 -28 7822 28
rect 7822 -28 7826 28
rect 7762 -32 7826 -28
rect 7842 28 7906 32
rect 7842 -28 7846 28
rect 7846 -28 7902 28
rect 7902 -28 7906 28
rect 7842 -32 7906 -28
rect 7922 28 7986 32
rect 7922 -28 7926 28
rect 7926 -28 7982 28
rect 7982 -28 7986 28
rect 7922 -32 7986 -28
rect 8002 28 8066 32
rect 8002 -28 8006 28
rect 8006 -28 8062 28
rect 8062 -28 8066 28
rect 8002 -32 8066 -28
rect 10862 28 10926 32
rect 10862 -28 10866 28
rect 10866 -28 10922 28
rect 10922 -28 10926 28
rect 10862 -32 10926 -28
rect 10942 28 11006 32
rect 10942 -28 10946 28
rect 10946 -28 11002 28
rect 11002 -28 11006 28
rect 10942 -32 11006 -28
rect 11022 28 11086 32
rect 11022 -28 11026 28
rect 11026 -28 11082 28
rect 11082 -28 11086 28
rect 11022 -32 11086 -28
rect 11102 28 11166 32
rect 11102 -28 11106 28
rect 11106 -28 11162 28
rect 11162 -28 11166 28
rect 11102 -32 11166 -28
rect 13962 28 14026 32
rect 13962 -28 13966 28
rect 13966 -28 14022 28
rect 14022 -28 14026 28
rect 13962 -32 14026 -28
rect 14042 28 14106 32
rect 14042 -28 14046 28
rect 14046 -28 14102 28
rect 14102 -28 14106 28
rect 14042 -32 14106 -28
rect 14122 28 14186 32
rect 14122 -28 14126 28
rect 14126 -28 14182 28
rect 14182 -28 14186 28
rect 14122 -32 14186 -28
rect 14202 28 14266 32
rect 14202 -28 14206 28
rect 14206 -28 14262 28
rect 14262 -28 14266 28
rect 14202 -32 14266 -28
rect 17062 28 17126 32
rect 17062 -28 17066 28
rect 17066 -28 17122 28
rect 17122 -28 17126 28
rect 17062 -32 17126 -28
rect 17142 28 17206 32
rect 17142 -28 17146 28
rect 17146 -28 17202 28
rect 17202 -28 17206 28
rect 17142 -32 17206 -28
rect 17222 28 17286 32
rect 17222 -28 17226 28
rect 17226 -28 17282 28
rect 17282 -28 17286 28
rect 17222 -32 17286 -28
rect 17302 28 17366 32
rect 17302 -28 17306 28
rect 17306 -28 17362 28
rect 17362 -28 17366 28
rect 17302 -32 17366 -28
<< metal4 >>
rect 3104 10368 3424 10928
rect 3104 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3272 10368
rect 3336 10304 3352 10368
rect 3416 10304 3424 10368
rect 3104 10160 3424 10304
rect 3104 9924 3146 10160
rect 3382 9924 3424 10160
rect 3104 9280 3424 9924
rect 3104 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3272 9280
rect 3336 9216 3352 9280
rect 3416 9216 3424 9280
rect 3104 8192 3424 9216
rect 3104 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3272 8192
rect 3336 8128 3352 8192
rect 3416 8128 3424 8192
rect 3104 7104 3424 8128
rect 3104 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3272 7104
rect 3336 7040 3352 7104
rect 3416 7040 3424 7104
rect 3104 6780 3424 7040
rect 3104 6544 3146 6780
rect 3382 6544 3424 6780
rect 3104 6016 3424 6544
rect 3104 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3272 6016
rect 3336 5952 3352 6016
rect 3416 5952 3424 6016
rect 3104 4928 3424 5952
rect 3104 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3272 4928
rect 3336 4864 3352 4928
rect 3416 4864 3424 4928
rect 3104 3840 3424 4864
rect 3104 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3272 3840
rect 3336 3776 3352 3840
rect 3416 3776 3424 3840
rect 3104 3400 3424 3776
rect 3104 3164 3146 3400
rect 3382 3164 3424 3400
rect 3104 2752 3424 3164
rect 3104 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3272 2752
rect 3336 2688 3352 2752
rect 3416 2688 3424 2752
rect 3104 1664 3424 2688
rect 3104 1600 3112 1664
rect 3176 1600 3192 1664
rect 3256 1600 3272 1664
rect 3336 1600 3352 1664
rect 3416 1600 3424 1664
rect 3104 576 3424 1600
rect 3104 512 3112 576
rect 3176 512 3192 576
rect 3256 512 3272 576
rect 3336 512 3352 576
rect 3416 512 3424 576
rect 3104 -48 3424 512
rect 4654 10912 4974 10928
rect 4654 10848 4662 10912
rect 4726 10848 4742 10912
rect 4806 10848 4822 10912
rect 4886 10848 4902 10912
rect 4966 10848 4974 10912
rect 4654 9824 4974 10848
rect 4654 9760 4662 9824
rect 4726 9760 4742 9824
rect 4806 9760 4822 9824
rect 4886 9760 4902 9824
rect 4966 9760 4974 9824
rect 4654 8736 4974 9760
rect 4654 8672 4662 8736
rect 4726 8672 4742 8736
rect 4806 8672 4822 8736
rect 4886 8672 4902 8736
rect 4966 8672 4974 8736
rect 4654 8470 4974 8672
rect 4654 8234 4696 8470
rect 4932 8234 4974 8470
rect 4654 7648 4974 8234
rect 4654 7584 4662 7648
rect 4726 7584 4742 7648
rect 4806 7584 4822 7648
rect 4886 7584 4902 7648
rect 4966 7584 4974 7648
rect 4654 6560 4974 7584
rect 4654 6496 4662 6560
rect 4726 6496 4742 6560
rect 4806 6496 4822 6560
rect 4886 6496 4902 6560
rect 4966 6496 4974 6560
rect 4654 5472 4974 6496
rect 4654 5408 4662 5472
rect 4726 5408 4742 5472
rect 4806 5408 4822 5472
rect 4886 5408 4902 5472
rect 4966 5408 4974 5472
rect 4654 5090 4974 5408
rect 4654 4854 4696 5090
rect 4932 4854 4974 5090
rect 4654 4384 4974 4854
rect 4654 4320 4662 4384
rect 4726 4320 4742 4384
rect 4806 4320 4822 4384
rect 4886 4320 4902 4384
rect 4966 4320 4974 4384
rect 4654 3296 4974 4320
rect 4654 3232 4662 3296
rect 4726 3232 4742 3296
rect 4806 3232 4822 3296
rect 4886 3232 4902 3296
rect 4966 3232 4974 3296
rect 4654 2208 4974 3232
rect 4654 2144 4662 2208
rect 4726 2144 4742 2208
rect 4806 2144 4822 2208
rect 4886 2144 4902 2208
rect 4966 2144 4974 2208
rect 4654 1120 4974 2144
rect 4654 1056 4662 1120
rect 4726 1056 4742 1120
rect 4806 1056 4822 1120
rect 4886 1056 4902 1120
rect 4966 1056 4974 1120
rect 4654 32 4974 1056
rect 4654 -32 4662 32
rect 4726 -32 4742 32
rect 4806 -32 4822 32
rect 4886 -32 4902 32
rect 4966 -32 4974 32
rect 4654 -48 4974 -32
rect 6204 10368 6524 10928
rect 6204 10304 6212 10368
rect 6276 10304 6292 10368
rect 6356 10304 6372 10368
rect 6436 10304 6452 10368
rect 6516 10304 6524 10368
rect 6204 10160 6524 10304
rect 6204 9924 6246 10160
rect 6482 9924 6524 10160
rect 6204 9280 6524 9924
rect 6204 9216 6212 9280
rect 6276 9216 6292 9280
rect 6356 9216 6372 9280
rect 6436 9216 6452 9280
rect 6516 9216 6524 9280
rect 6204 8192 6524 9216
rect 6204 8128 6212 8192
rect 6276 8128 6292 8192
rect 6356 8128 6372 8192
rect 6436 8128 6452 8192
rect 6516 8128 6524 8192
rect 6204 7104 6524 8128
rect 6204 7040 6212 7104
rect 6276 7040 6292 7104
rect 6356 7040 6372 7104
rect 6436 7040 6452 7104
rect 6516 7040 6524 7104
rect 6204 6780 6524 7040
rect 6204 6544 6246 6780
rect 6482 6544 6524 6780
rect 6204 6016 6524 6544
rect 6204 5952 6212 6016
rect 6276 5952 6292 6016
rect 6356 5952 6372 6016
rect 6436 5952 6452 6016
rect 6516 5952 6524 6016
rect 6204 4928 6524 5952
rect 6204 4864 6212 4928
rect 6276 4864 6292 4928
rect 6356 4864 6372 4928
rect 6436 4864 6452 4928
rect 6516 4864 6524 4928
rect 6204 3840 6524 4864
rect 6204 3776 6212 3840
rect 6276 3776 6292 3840
rect 6356 3776 6372 3840
rect 6436 3776 6452 3840
rect 6516 3776 6524 3840
rect 6204 3400 6524 3776
rect 6204 3164 6246 3400
rect 6482 3164 6524 3400
rect 6204 2752 6524 3164
rect 6204 2688 6212 2752
rect 6276 2688 6292 2752
rect 6356 2688 6372 2752
rect 6436 2688 6452 2752
rect 6516 2688 6524 2752
rect 6204 1664 6524 2688
rect 6204 1600 6212 1664
rect 6276 1600 6292 1664
rect 6356 1600 6372 1664
rect 6436 1600 6452 1664
rect 6516 1600 6524 1664
rect 6204 576 6524 1600
rect 6204 512 6212 576
rect 6276 512 6292 576
rect 6356 512 6372 576
rect 6436 512 6452 576
rect 6516 512 6524 576
rect 6204 -48 6524 512
rect 7754 10912 8074 10928
rect 7754 10848 7762 10912
rect 7826 10848 7842 10912
rect 7906 10848 7922 10912
rect 7986 10848 8002 10912
rect 8066 10848 8074 10912
rect 7754 9824 8074 10848
rect 7754 9760 7762 9824
rect 7826 9760 7842 9824
rect 7906 9760 7922 9824
rect 7986 9760 8002 9824
rect 8066 9760 8074 9824
rect 7754 8736 8074 9760
rect 7754 8672 7762 8736
rect 7826 8672 7842 8736
rect 7906 8672 7922 8736
rect 7986 8672 8002 8736
rect 8066 8672 8074 8736
rect 7754 8470 8074 8672
rect 7754 8234 7796 8470
rect 8032 8234 8074 8470
rect 7754 7648 8074 8234
rect 7754 7584 7762 7648
rect 7826 7584 7842 7648
rect 7906 7584 7922 7648
rect 7986 7584 8002 7648
rect 8066 7584 8074 7648
rect 7754 6560 8074 7584
rect 7754 6496 7762 6560
rect 7826 6496 7842 6560
rect 7906 6496 7922 6560
rect 7986 6496 8002 6560
rect 8066 6496 8074 6560
rect 7754 5472 8074 6496
rect 7754 5408 7762 5472
rect 7826 5408 7842 5472
rect 7906 5408 7922 5472
rect 7986 5408 8002 5472
rect 8066 5408 8074 5472
rect 7754 5090 8074 5408
rect 7754 4854 7796 5090
rect 8032 4854 8074 5090
rect 7754 4384 8074 4854
rect 7754 4320 7762 4384
rect 7826 4320 7842 4384
rect 7906 4320 7922 4384
rect 7986 4320 8002 4384
rect 8066 4320 8074 4384
rect 7754 3296 8074 4320
rect 7754 3232 7762 3296
rect 7826 3232 7842 3296
rect 7906 3232 7922 3296
rect 7986 3232 8002 3296
rect 8066 3232 8074 3296
rect 7754 2208 8074 3232
rect 7754 2144 7762 2208
rect 7826 2144 7842 2208
rect 7906 2144 7922 2208
rect 7986 2144 8002 2208
rect 8066 2144 8074 2208
rect 7754 1120 8074 2144
rect 7754 1056 7762 1120
rect 7826 1056 7842 1120
rect 7906 1056 7922 1120
rect 7986 1056 8002 1120
rect 8066 1056 8074 1120
rect 7754 32 8074 1056
rect 7754 -32 7762 32
rect 7826 -32 7842 32
rect 7906 -32 7922 32
rect 7986 -32 8002 32
rect 8066 -32 8074 32
rect 7754 -48 8074 -32
rect 9304 10368 9624 10928
rect 9304 10304 9312 10368
rect 9376 10304 9392 10368
rect 9456 10304 9472 10368
rect 9536 10304 9552 10368
rect 9616 10304 9624 10368
rect 9304 10160 9624 10304
rect 9304 9924 9346 10160
rect 9582 9924 9624 10160
rect 9304 9280 9624 9924
rect 9304 9216 9312 9280
rect 9376 9216 9392 9280
rect 9456 9216 9472 9280
rect 9536 9216 9552 9280
rect 9616 9216 9624 9280
rect 9304 8192 9624 9216
rect 9304 8128 9312 8192
rect 9376 8128 9392 8192
rect 9456 8128 9472 8192
rect 9536 8128 9552 8192
rect 9616 8128 9624 8192
rect 9304 7104 9624 8128
rect 9304 7040 9312 7104
rect 9376 7040 9392 7104
rect 9456 7040 9472 7104
rect 9536 7040 9552 7104
rect 9616 7040 9624 7104
rect 9304 6780 9624 7040
rect 9304 6544 9346 6780
rect 9582 6544 9624 6780
rect 9304 6016 9624 6544
rect 9304 5952 9312 6016
rect 9376 5952 9392 6016
rect 9456 5952 9472 6016
rect 9536 5952 9552 6016
rect 9616 5952 9624 6016
rect 9304 4928 9624 5952
rect 9304 4864 9312 4928
rect 9376 4864 9392 4928
rect 9456 4864 9472 4928
rect 9536 4864 9552 4928
rect 9616 4864 9624 4928
rect 9304 3840 9624 4864
rect 9304 3776 9312 3840
rect 9376 3776 9392 3840
rect 9456 3776 9472 3840
rect 9536 3776 9552 3840
rect 9616 3776 9624 3840
rect 9304 3400 9624 3776
rect 9304 3164 9346 3400
rect 9582 3164 9624 3400
rect 9304 2752 9624 3164
rect 9304 2688 9312 2752
rect 9376 2688 9392 2752
rect 9456 2688 9472 2752
rect 9536 2688 9552 2752
rect 9616 2688 9624 2752
rect 9304 1664 9624 2688
rect 9304 1600 9312 1664
rect 9376 1600 9392 1664
rect 9456 1600 9472 1664
rect 9536 1600 9552 1664
rect 9616 1600 9624 1664
rect 9304 576 9624 1600
rect 9304 512 9312 576
rect 9376 512 9392 576
rect 9456 512 9472 576
rect 9536 512 9552 576
rect 9616 512 9624 576
rect 9304 -48 9624 512
rect 10854 10912 11174 10928
rect 10854 10848 10862 10912
rect 10926 10848 10942 10912
rect 11006 10848 11022 10912
rect 11086 10848 11102 10912
rect 11166 10848 11174 10912
rect 10854 9824 11174 10848
rect 10854 9760 10862 9824
rect 10926 9760 10942 9824
rect 11006 9760 11022 9824
rect 11086 9760 11102 9824
rect 11166 9760 11174 9824
rect 10854 8736 11174 9760
rect 10854 8672 10862 8736
rect 10926 8672 10942 8736
rect 11006 8672 11022 8736
rect 11086 8672 11102 8736
rect 11166 8672 11174 8736
rect 10854 8470 11174 8672
rect 10854 8234 10896 8470
rect 11132 8234 11174 8470
rect 10854 7648 11174 8234
rect 10854 7584 10862 7648
rect 10926 7584 10942 7648
rect 11006 7584 11022 7648
rect 11086 7584 11102 7648
rect 11166 7584 11174 7648
rect 10854 6560 11174 7584
rect 10854 6496 10862 6560
rect 10926 6496 10942 6560
rect 11006 6496 11022 6560
rect 11086 6496 11102 6560
rect 11166 6496 11174 6560
rect 10854 5472 11174 6496
rect 10854 5408 10862 5472
rect 10926 5408 10942 5472
rect 11006 5408 11022 5472
rect 11086 5408 11102 5472
rect 11166 5408 11174 5472
rect 10854 5090 11174 5408
rect 10854 4854 10896 5090
rect 11132 4854 11174 5090
rect 10854 4384 11174 4854
rect 10854 4320 10862 4384
rect 10926 4320 10942 4384
rect 11006 4320 11022 4384
rect 11086 4320 11102 4384
rect 11166 4320 11174 4384
rect 10854 3296 11174 4320
rect 10854 3232 10862 3296
rect 10926 3232 10942 3296
rect 11006 3232 11022 3296
rect 11086 3232 11102 3296
rect 11166 3232 11174 3296
rect 10854 2208 11174 3232
rect 10854 2144 10862 2208
rect 10926 2144 10942 2208
rect 11006 2144 11022 2208
rect 11086 2144 11102 2208
rect 11166 2144 11174 2208
rect 10854 1120 11174 2144
rect 10854 1056 10862 1120
rect 10926 1056 10942 1120
rect 11006 1056 11022 1120
rect 11086 1056 11102 1120
rect 11166 1056 11174 1120
rect 10854 32 11174 1056
rect 10854 -32 10862 32
rect 10926 -32 10942 32
rect 11006 -32 11022 32
rect 11086 -32 11102 32
rect 11166 -32 11174 32
rect 10854 -48 11174 -32
rect 12404 10368 12724 10928
rect 12404 10304 12412 10368
rect 12476 10304 12492 10368
rect 12556 10304 12572 10368
rect 12636 10304 12652 10368
rect 12716 10304 12724 10368
rect 12404 10160 12724 10304
rect 12404 9924 12446 10160
rect 12682 9924 12724 10160
rect 12404 9280 12724 9924
rect 12404 9216 12412 9280
rect 12476 9216 12492 9280
rect 12556 9216 12572 9280
rect 12636 9216 12652 9280
rect 12716 9216 12724 9280
rect 12404 8192 12724 9216
rect 12404 8128 12412 8192
rect 12476 8128 12492 8192
rect 12556 8128 12572 8192
rect 12636 8128 12652 8192
rect 12716 8128 12724 8192
rect 12404 7104 12724 8128
rect 12404 7040 12412 7104
rect 12476 7040 12492 7104
rect 12556 7040 12572 7104
rect 12636 7040 12652 7104
rect 12716 7040 12724 7104
rect 12404 6780 12724 7040
rect 12404 6544 12446 6780
rect 12682 6544 12724 6780
rect 12404 6016 12724 6544
rect 12404 5952 12412 6016
rect 12476 5952 12492 6016
rect 12556 5952 12572 6016
rect 12636 5952 12652 6016
rect 12716 5952 12724 6016
rect 12404 4928 12724 5952
rect 12404 4864 12412 4928
rect 12476 4864 12492 4928
rect 12556 4864 12572 4928
rect 12636 4864 12652 4928
rect 12716 4864 12724 4928
rect 12404 3840 12724 4864
rect 12404 3776 12412 3840
rect 12476 3776 12492 3840
rect 12556 3776 12572 3840
rect 12636 3776 12652 3840
rect 12716 3776 12724 3840
rect 12404 3400 12724 3776
rect 12404 3164 12446 3400
rect 12682 3164 12724 3400
rect 12404 2752 12724 3164
rect 12404 2688 12412 2752
rect 12476 2688 12492 2752
rect 12556 2688 12572 2752
rect 12636 2688 12652 2752
rect 12716 2688 12724 2752
rect 12404 1664 12724 2688
rect 12404 1600 12412 1664
rect 12476 1600 12492 1664
rect 12556 1600 12572 1664
rect 12636 1600 12652 1664
rect 12716 1600 12724 1664
rect 12404 576 12724 1600
rect 12404 512 12412 576
rect 12476 512 12492 576
rect 12556 512 12572 576
rect 12636 512 12652 576
rect 12716 512 12724 576
rect 12404 -48 12724 512
rect 13954 10912 14274 10928
rect 13954 10848 13962 10912
rect 14026 10848 14042 10912
rect 14106 10848 14122 10912
rect 14186 10848 14202 10912
rect 14266 10848 14274 10912
rect 13954 9824 14274 10848
rect 13954 9760 13962 9824
rect 14026 9760 14042 9824
rect 14106 9760 14122 9824
rect 14186 9760 14202 9824
rect 14266 9760 14274 9824
rect 13954 8736 14274 9760
rect 13954 8672 13962 8736
rect 14026 8672 14042 8736
rect 14106 8672 14122 8736
rect 14186 8672 14202 8736
rect 14266 8672 14274 8736
rect 13954 8470 14274 8672
rect 13954 8234 13996 8470
rect 14232 8234 14274 8470
rect 13954 7648 14274 8234
rect 13954 7584 13962 7648
rect 14026 7584 14042 7648
rect 14106 7584 14122 7648
rect 14186 7584 14202 7648
rect 14266 7584 14274 7648
rect 13954 6560 14274 7584
rect 13954 6496 13962 6560
rect 14026 6496 14042 6560
rect 14106 6496 14122 6560
rect 14186 6496 14202 6560
rect 14266 6496 14274 6560
rect 13954 5472 14274 6496
rect 13954 5408 13962 5472
rect 14026 5408 14042 5472
rect 14106 5408 14122 5472
rect 14186 5408 14202 5472
rect 14266 5408 14274 5472
rect 13954 5090 14274 5408
rect 13954 4854 13996 5090
rect 14232 4854 14274 5090
rect 13954 4384 14274 4854
rect 13954 4320 13962 4384
rect 14026 4320 14042 4384
rect 14106 4320 14122 4384
rect 14186 4320 14202 4384
rect 14266 4320 14274 4384
rect 13954 3296 14274 4320
rect 13954 3232 13962 3296
rect 14026 3232 14042 3296
rect 14106 3232 14122 3296
rect 14186 3232 14202 3296
rect 14266 3232 14274 3296
rect 13954 2208 14274 3232
rect 13954 2144 13962 2208
rect 14026 2144 14042 2208
rect 14106 2144 14122 2208
rect 14186 2144 14202 2208
rect 14266 2144 14274 2208
rect 13954 1120 14274 2144
rect 13954 1056 13962 1120
rect 14026 1056 14042 1120
rect 14106 1056 14122 1120
rect 14186 1056 14202 1120
rect 14266 1056 14274 1120
rect 13954 32 14274 1056
rect 13954 -32 13962 32
rect 14026 -32 14042 32
rect 14106 -32 14122 32
rect 14186 -32 14202 32
rect 14266 -32 14274 32
rect 13954 -48 14274 -32
rect 15504 10368 15824 10928
rect 15504 10304 15512 10368
rect 15576 10304 15592 10368
rect 15656 10304 15672 10368
rect 15736 10304 15752 10368
rect 15816 10304 15824 10368
rect 15504 10160 15824 10304
rect 15504 9924 15546 10160
rect 15782 9924 15824 10160
rect 15504 9280 15824 9924
rect 15504 9216 15512 9280
rect 15576 9216 15592 9280
rect 15656 9216 15672 9280
rect 15736 9216 15752 9280
rect 15816 9216 15824 9280
rect 15504 8192 15824 9216
rect 15504 8128 15512 8192
rect 15576 8128 15592 8192
rect 15656 8128 15672 8192
rect 15736 8128 15752 8192
rect 15816 8128 15824 8192
rect 15504 7104 15824 8128
rect 15504 7040 15512 7104
rect 15576 7040 15592 7104
rect 15656 7040 15672 7104
rect 15736 7040 15752 7104
rect 15816 7040 15824 7104
rect 15504 6780 15824 7040
rect 15504 6544 15546 6780
rect 15782 6544 15824 6780
rect 15504 6016 15824 6544
rect 15504 5952 15512 6016
rect 15576 5952 15592 6016
rect 15656 5952 15672 6016
rect 15736 5952 15752 6016
rect 15816 5952 15824 6016
rect 15504 4928 15824 5952
rect 15504 4864 15512 4928
rect 15576 4864 15592 4928
rect 15656 4864 15672 4928
rect 15736 4864 15752 4928
rect 15816 4864 15824 4928
rect 15504 3840 15824 4864
rect 15504 3776 15512 3840
rect 15576 3776 15592 3840
rect 15656 3776 15672 3840
rect 15736 3776 15752 3840
rect 15816 3776 15824 3840
rect 15504 3400 15824 3776
rect 15504 3164 15546 3400
rect 15782 3164 15824 3400
rect 15504 2752 15824 3164
rect 15504 2688 15512 2752
rect 15576 2688 15592 2752
rect 15656 2688 15672 2752
rect 15736 2688 15752 2752
rect 15816 2688 15824 2752
rect 15504 1664 15824 2688
rect 15504 1600 15512 1664
rect 15576 1600 15592 1664
rect 15656 1600 15672 1664
rect 15736 1600 15752 1664
rect 15816 1600 15824 1664
rect 15504 576 15824 1600
rect 15504 512 15512 576
rect 15576 512 15592 576
rect 15656 512 15672 576
rect 15736 512 15752 576
rect 15816 512 15824 576
rect 15504 -48 15824 512
rect 17054 10912 17374 10928
rect 17054 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17222 10912
rect 17286 10848 17302 10912
rect 17366 10848 17374 10912
rect 17054 9824 17374 10848
rect 17054 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17222 9824
rect 17286 9760 17302 9824
rect 17366 9760 17374 9824
rect 17054 8736 17374 9760
rect 17054 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17222 8736
rect 17286 8672 17302 8736
rect 17366 8672 17374 8736
rect 17054 8470 17374 8672
rect 17054 8234 17096 8470
rect 17332 8234 17374 8470
rect 17054 7648 17374 8234
rect 17054 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17222 7648
rect 17286 7584 17302 7648
rect 17366 7584 17374 7648
rect 17054 6560 17374 7584
rect 17054 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17222 6560
rect 17286 6496 17302 6560
rect 17366 6496 17374 6560
rect 17054 5472 17374 6496
rect 17054 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17222 5472
rect 17286 5408 17302 5472
rect 17366 5408 17374 5472
rect 17054 5090 17374 5408
rect 17054 4854 17096 5090
rect 17332 4854 17374 5090
rect 17054 4384 17374 4854
rect 17054 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17222 4384
rect 17286 4320 17302 4384
rect 17366 4320 17374 4384
rect 17054 3296 17374 4320
rect 17054 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17222 3296
rect 17286 3232 17302 3296
rect 17366 3232 17374 3296
rect 17054 2208 17374 3232
rect 17054 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17222 2208
rect 17286 2144 17302 2208
rect 17366 2144 17374 2208
rect 17054 1120 17374 2144
rect 17054 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17222 1120
rect 17286 1056 17302 1120
rect 17366 1056 17374 1120
rect 17054 32 17374 1056
rect 17054 -32 17062 32
rect 17126 -32 17142 32
rect 17206 -32 17222 32
rect 17286 -32 17302 32
rect 17366 -32 17374 32
rect 17054 -48 17374 -32
<< via4 >>
rect 3146 9924 3382 10160
rect 3146 6544 3382 6780
rect 3146 3164 3382 3400
rect 4696 8234 4932 8470
rect 4696 4854 4932 5090
rect 6246 9924 6482 10160
rect 6246 6544 6482 6780
rect 6246 3164 6482 3400
rect 7796 8234 8032 8470
rect 7796 4854 8032 5090
rect 9346 9924 9582 10160
rect 9346 6544 9582 6780
rect 9346 3164 9582 3400
rect 10896 8234 11132 8470
rect 10896 4854 11132 5090
rect 12446 9924 12682 10160
rect 12446 6544 12682 6780
rect 12446 3164 12682 3400
rect 13996 8234 14232 8470
rect 13996 4854 14232 5090
rect 15546 9924 15782 10160
rect 15546 6544 15782 6780
rect 15546 3164 15782 3400
rect 17096 8234 17332 8470
rect 17096 4854 17332 5090
<< metal5 >>
rect 0 10160 18860 10202
rect 0 9924 3146 10160
rect 3382 9924 6246 10160
rect 6482 9924 9346 10160
rect 9582 9924 12446 10160
rect 12682 9924 15546 10160
rect 15782 9924 18860 10160
rect 0 9882 18860 9924
rect 0 8470 18860 8512
rect 0 8234 4696 8470
rect 4932 8234 7796 8470
rect 8032 8234 10896 8470
rect 11132 8234 13996 8470
rect 14232 8234 17096 8470
rect 17332 8234 18860 8470
rect 0 8192 18860 8234
rect 0 6780 18860 6822
rect 0 6544 3146 6780
rect 3382 6544 6246 6780
rect 6482 6544 9346 6780
rect 9582 6544 12446 6780
rect 12682 6544 15546 6780
rect 15782 6544 18860 6780
rect 0 6502 18860 6544
rect 0 5090 18860 5132
rect 0 4854 4696 5090
rect 4932 4854 7796 5090
rect 8032 4854 10896 5090
rect 11132 4854 13996 5090
rect 14232 4854 17096 5090
rect 17332 4854 18860 5090
rect 0 4812 18860 4854
rect 0 3400 18860 3442
rect 0 3164 3146 3400
rect 3382 3164 6246 3400
rect 6482 3164 9346 3400
rect 9582 3164 12446 3400
rect 12682 3164 15546 3400
rect 15782 3164 18860 3400
rect 0 3122 18860 3164
use sky130_fd_sc_hd__decap_3  PHY_2 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 0 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1636915332
transform 1 0 0 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 276 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1012 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1196 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_23 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2116 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15
timestamp 1636915332
transform 1 0 1380 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__SET_B OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 2392 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 276 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_14
timestamp 1636915332
transform 1 0 1288 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _339_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 3404 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1636915332
transform 1 0 2392 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1636915332
transform 1 0 2392 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37
timestamp 1636915332
transform 1 0 3404 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2484 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _338_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 3956 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 4692 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1636915332
transform 1 0 3588 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43
timestamp 1636915332
transform 1 0 3956 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_1  _447_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2484 0 -1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _361_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5244 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_2  _311_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4876 0 -1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1636915332
transform 1 0 4784 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1636915332
transform 1 0 4784 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_51
timestamp 1636915332
transform 1 0 4692 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4876 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51
timestamp 1636915332
transform 1 0 4692 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _388_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 6072 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _387_
timestamp 1636915332
transform -1 0 6900 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _362_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5796 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1636915332
transform 1 0 5980 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64
timestamp 1636915332
transform 1 0 5888 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1636915332
transform 1 0 7176 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1636915332
transform 1 0 7176 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_79
timestamp 1636915332
transform 1 0 7268 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_75
timestamp 1636915332
transform 1 0 6900 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75
timestamp 1636915332
transform 1 0 6900 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__SET_B
timestamp 1636915332
transform -1 0 7176 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_1  _293_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 9200 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1636915332
transform 1 0 8372 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _458_
timestamp 1636915332
transform 1 0 7360 0 -1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_0_79
timestamp 1636915332
transform 1 0 7268 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_1  _365_
timestamp 1636915332
transform 1 0 10028 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _292_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 10028 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1636915332
transform 1 0 9568 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1636915332
transform 1 0 9568 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1636915332
transform 1 0 10028 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_101
timestamp 1636915332
transform 1 0 9292 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_105
timestamp 1636915332
transform 1 0 9660 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100
timestamp 1636915332
transform 1 0 9200 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _407_
timestamp 1636915332
transform 1 0 10304 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1636915332
transform 1 0 10764 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_121
timestamp 1636915332
transform 1 0 11132 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116
timestamp 1636915332
transform 1 0 10672 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__RESET_B
timestamp 1636915332
transform -1 0 11592 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_118
timestamp 1636915332
transform 1 0 10856 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131
timestamp 1636915332
transform 1 0 12052 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_140
timestamp 1636915332
transform 1 0 12880 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_144
timestamp 1636915332
transform 1 0 13248 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1636915332
transform 1 0 11960 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1636915332
transform 1 0 13156 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1636915332
transform 1 0 11960 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _294_
timestamp 1636915332
transform 1 0 11592 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _295_
timestamp 1636915332
transform 1 0 12144 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _457_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 12052 0 -1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_0_157
timestamp 1636915332
transform 1 0 14444 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_165
timestamp 1636915332
transform 1 0 15180 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_170
timestamp 1636915332
transform 1 0 15640 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1636915332
transform 1 0 14352 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1636915332
transform 1 0 15548 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1636915332
transform 1 0 14352 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _332_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 15180 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _364_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 13984 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _449_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 16560 0 -1 1088
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_0_183
timestamp 1636915332
transform 1 0 16836 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_193
timestamp 1636915332
transform 1 0 17756 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_180
timestamp 1636915332
transform 1 0 16560 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1636915332
transform 1 0 16744 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1636915332
transform 1 0 17940 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1636915332
transform 1 0 16744 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _326_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 17204 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _327_
timestamp 1636915332
transform 1 0 18032 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _420_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 16836 0 -1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1636915332
transform -1 0 18860 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1636915332
transform -1 0 18860 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 18308 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1636915332
transform 1 0 1012 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1636915332
transform 1 0 276 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1636915332
transform 1 0 0 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1636915332
transform 1 0 1196 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtn_1  _448_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1288 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__RESET_B
timestamp 1636915332
transform 1 0 3956 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_34
timestamp 1636915332
transform 1 0 3128 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_45
timestamp 1636915332
transform 1 0 4140 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1636915332
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1636915332
transform -1 0 3956 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _315_
timestamp 1636915332
transform 1 0 3220 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_57
timestamp 1636915332
transform 1 0 5244 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1636915332
transform 1 0 5980 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _363_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5336 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _413_
timestamp 1636915332
transform 1 0 6072 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_2_75
timestamp 1636915332
transform 1 0 6900 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1636915332
transform 1 0 8004 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1636915332
transform 1 0 8372 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _291_
timestamp 1636915332
transform -1 0 9200 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_100
timestamp 1636915332
transform 1 0 9200 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_114
timestamp 1636915332
transform 1 0 10488 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1636915332
transform 1 0 10764 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1636915332
transform 1 0 11224 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _279_
timestamp 1636915332
transform 1 0 10856 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _366_
timestamp 1636915332
transform 1 0 10212 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1636915332
transform 1 0 9384 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_125
timestamp 1636915332
transform 1 0 11500 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_133
timestamp 1636915332
transform 1 0 12236 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1636915332
transform 1 0 13156 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _410_
timestamp 1636915332
transform 1 0 13248 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _411_
timestamp 1636915332
transform 1 0 12328 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__RESET_B
timestamp 1636915332
transform 1 0 15640 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__RESET_B
timestamp 1636915332
transform 1 0 14260 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_153
timestamp 1636915332
transform 1 0 14076 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_157
timestamp 1636915332
transform 1 0 14444 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_166
timestamp 1636915332
transform 1 0 15272 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1636915332
transform 1 0 15548 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _330_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 15272 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _433_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 15824 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1636915332
transform 1 0 17940 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _328_
timestamp 1636915332
transform -1 0 18400 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1636915332
transform -1 0 17940 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1636915332
transform -1 0 18584 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1636915332
transform -1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1636915332
transform 1 0 276 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1636915332
transform 1 0 0 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _446_
timestamp 1636915332
transform 1 0 552 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__RESET_B
timestamp 1636915332
transform 1 0 2484 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_29
timestamp 1636915332
transform 1 0 2668 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_43
timestamp 1636915332
transform 1 0 3956 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1636915332
transform 1 0 2392 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _335_
timestamp 1636915332
transform -1 0 3680 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _336_
timestamp 1636915332
transform -1 0 3128 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _337__6
timestamp 1636915332
transform -1 0 3404 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1636915332
transform -1 0 3956 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_51
timestamp 1636915332
transform 1 0 4692 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1636915332
transform 1 0 5704 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1636915332
transform 1 0 4784 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _392_
timestamp 1636915332
transform 1 0 4876 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1636915332
transform -1 0 6900 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__459__RESET_B
timestamp 1636915332
transform 1 0 6992 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_75
timestamp 1636915332
transform 1 0 6900 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1636915332
transform 1 0 7176 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _290_
timestamp 1636915332
transform -1 0 9476 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _459_
timestamp 1636915332
transform 1 0 7268 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_3_103
timestamp 1636915332
transform 1 0 9476 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_124
timestamp 1636915332
transform 1 0 11408 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1636915332
transform 1 0 9568 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1636915332
transform 1 0 11132 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _367_
timestamp 1636915332
transform 1 0 9660 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp 1636915332
transform -1 0 11132 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_131
timestamp 1636915332
transform 1 0 12052 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_135
timestamp 1636915332
transform 1 0 12420 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_142
timestamp 1636915332
transform 1 0 13064 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1636915332
transform 1 0 11960 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1636915332
transform 1 0 12512 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1636915332
transform -1 0 13064 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_150
timestamp 1636915332
transform 1 0 13800 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1636915332
transform 1 0 14352 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _281_
timestamp 1636915332
transform 1 0 14720 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _329_
timestamp 1636915332
transform -1 0 14720 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _331_
timestamp 1636915332
transform -1 0 14352 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _421_
timestamp 1636915332
transform 1 0 15272 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_3_183
timestamp 1636915332
transform 1 0 16836 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_195
timestamp 1636915332
transform 1 0 17940 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1636915332
transform 1 0 16744 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_201
timestamp 1636915332
transform 1 0 18492 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1636915332
transform -1 0 18860 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_11
timestamp 1636915332
transform 1 0 1012 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_14
timestamp 1636915332
transform 1 0 1288 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1636915332
transform 1 0 276 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1636915332
transform 1 0 0 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1636915332
transform 1 0 1196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_26
timestamp 1636915332
transform 1 0 2392 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_32
timestamp 1636915332
transform 1 0 2944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_37
timestamp 1636915332
transform 1 0 3404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1636915332
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _334_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3680 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _342_
timestamp 1636915332
transform -1 0 3404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_59
timestamp 1636915332
transform 1 0 5428 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1636915332
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1636915332
transform 1 0 5980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _289_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 7268 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _318_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 6808 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _391_
timestamp 1636915332
transform -1 0 5428 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__SET_B
timestamp 1636915332
transform 1 0 7912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_83
timestamp 1636915332
transform 1 0 7636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1636915332
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _308__5
timestamp 1636915332
transform 1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _312_
timestamp 1636915332
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _453_
timestamp 1636915332
transform 1 0 8464 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_4_113
timestamp 1636915332
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1636915332
transform 1 0 10764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _405_
timestamp 1636915332
transform 1 0 10856 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_4_127
timestamp 1636915332
transform 1 0 11684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1636915332
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _282_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 12236 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _287_
timestamp 1636915332
transform 1 0 13248 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _288_
timestamp 1636915332
transform -1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__SET_B
timestamp 1636915332
transform 1 0 15272 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__RESET_B
timestamp 1636915332
transform 1 0 15640 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_168
timestamp 1636915332
transform 1 0 15456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1636915332
transform 1 0 15548 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _422_
timestamp 1636915332
transform 1 0 13800 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _436_
timestamp 1636915332
transform -1 0 17940 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1636915332
transform -1 0 18308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_196
timestamp 1636915332
transform 1 0 18032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1636915332
transform 1 0 17940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1636915332
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1636915332
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__RESET_B
timestamp 1636915332
transform 1 0 2116 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1636915332
transform 1 0 0 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _454_
timestamp 1636915332
transform 1 0 276 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1636915332
transform -1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1636915332
transform 1 0 2392 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_25
timestamp 1636915332
transform 1 0 2300 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _296_
timestamp 1636915332
transform -1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_30
timestamp 1636915332
transform 1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_36
timestamp 1636915332
transform 1 0 3312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _341_
timestamp 1636915332
transform -1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_43
timestamp 1636915332
transform 1 0 3956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _333_
timestamp 1636915332
transform 1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1636915332
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_51
timestamp 1636915332
transform 1 0 4692 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_53
timestamp 1636915332
transform 1 0 4876 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1636915332
transform 1 0 4784 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _403_
timestamp 1636915332
transform 1 0 5428 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer4 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 6256 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_5_75
timestamp 1636915332
transform 1 0 6900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_87
timestamp 1636915332
transform 1 0 8004 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_92
timestamp 1636915332
transform 1 0 8464 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1636915332
transform 1 0 7176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _284_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _286_
timestamp 1636915332
transform 1 0 8096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _319_
timestamp 1636915332
transform -1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__SET_B
timestamp 1636915332
transform 1 0 9384 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_100
timestamp 1636915332
transform 1 0 9200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_105
timestamp 1636915332
transform 1 0 9660 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1636915332
transform 1 0 9568 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1636915332
transform -1 0 10028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _460_
timestamp 1636915332
transform 1 0 10028 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_5_131
timestamp 1636915332
transform 1 0 12052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_140
timestamp 1636915332
transform 1 0 12880 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_146
timestamp 1636915332
transform 1 0 13432 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1636915332
transform 1 0 11960 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _355_
timestamp 1636915332
transform 1 0 12236 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_2  _357_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 14352 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_157
timestamp 1636915332
transform 1 0 14444 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1636915332
transform 1 0 14352 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _354_
timestamp 1636915332
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _434_
timestamp 1636915332
transform -1 0 16744 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_5_183
timestamp 1636915332
transform 1 0 16836 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_195
timestamp 1636915332
transform 1 0 17940 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1636915332
transform 1 0 16744 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_201
timestamp 1636915332
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1636915332
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1636915332
transform 1 0 1012 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_14
timestamp 1636915332
transform 1 0 1288 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1636915332
transform 1 0 276 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1636915332
transform 1 0 276 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1636915332
transform 1 0 0 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1636915332
transform 1 0 0 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1636915332
transform 1 0 1196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _307_
timestamp 1636915332
transform -1 0 2300 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_1  _455_
timestamp 1636915332
transform 1 0 460 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__o21ai_1  _306_
timestamp 1636915332
transform -1 0 2852 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _305_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2300 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1636915332
transform -1 0 3128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _298_
timestamp 1636915332
transform 1 0 2852 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1636915332
transform 1 0 2392 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2ai_1  _303_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3220 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _299_
timestamp 1636915332
transform -1 0 4232 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1636915332
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_34
timestamp 1636915332
transform 1 0 3128 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp 1636915332
transform 1 0 3404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  rebuffer3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 4600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _302_
timestamp 1636915332
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1636915332
transform 1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_48
timestamp 1636915332
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _316_
timestamp 1636915332
transform 1 0 4968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _309_
timestamp 1636915332
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1636915332
transform 1 0 4784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_57
timestamp 1636915332
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_53
timestamp 1636915332
transform 1 0 4876 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_pll_clk
timestamp 1636915332
transform -1 0 7176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _325_
timestamp 1636915332
transform 1 0 6256 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _317_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 6624 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1636915332
transform 1 0 5980 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_71
timestamp 1636915332
transform 1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_65
timestamp 1636915332
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_72
timestamp 1636915332
transform 1 0 6624 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_50
timestamp 1636915332
transform 1 0 4600 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__RESET_B
timestamp 1636915332
transform 1 0 8464 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_94
timestamp 1636915332
transform 1 0 8648 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1636915332
transform 1 0 7176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1636915332
transform 1 0 8372 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _285_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8372 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _323_
timestamp 1636915332
transform 1 0 8924 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _324_
timestamp 1636915332
transform 1 0 7268 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1636915332
transform 1 0 8096 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _369_
timestamp 1636915332
transform 1 0 9568 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _322_
timestamp 1636915332
transform 1 0 9660 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1636915332
transform 1 0 9568 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_100
timestamp 1636915332
transform 1 0 9200 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_111
timestamp 1636915332
transform 1 0 10212 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_102
timestamp 1636915332
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _409_
timestamp 1636915332
transform 1 0 10488 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_1  _344_
timestamp 1636915332
transform 1 0 11408 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1636915332
transform 1 0 10764 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_123
timestamp 1636915332
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_118
timestamp 1636915332
transform 1 0 10856 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _370_
timestamp 1636915332
transform 1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _345_
timestamp 1636915332
transform 1 0 12420 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1636915332
transform 1 0 11960 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_134
timestamp 1636915332
transform 1 0 12328 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_130
timestamp 1636915332
transform 1 0 11960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__SET_B
timestamp 1636915332
transform 1 0 12236 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1636915332
transform 1 0 13156 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_144
timestamp 1636915332
transform 1 0 13248 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_142
timestamp 1636915332
transform 1 0 13064 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _445_
timestamp 1636915332
transform 1 0 12420 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _417_
timestamp 1636915332
transform 1 0 14536 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _356_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 13892 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1636915332
transform 1 0 14352 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_157
timestamp 1636915332
transform 1 0 14444 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_150
timestamp 1636915332
transform 1 0 13800 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__RESET_B
timestamp 1636915332
transform 1 0 14536 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1636915332
transform 1 0 15548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_170
timestamp 1636915332
transform 1 0 15640 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__SET_B
timestamp 1636915332
transform 1 0 15364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_4  _437_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 15732 0 1 3264
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_1  _430_
timestamp 1636915332
transform -1 0 16560 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1636915332
transform -1 0 18308 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_180
timestamp 1636915332
transform 1 0 16560 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_183
timestamp 1636915332
transform 1 0 16836 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_195
timestamp 1636915332
transform 1 0 17940 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1636915332
transform 1 0 16744 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1636915332
transform 1 0 17940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  split2
timestamp 1636915332
transform -1 0 18400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_200
timestamp 1636915332
transform 1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1636915332
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1636915332
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1636915332
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_14
timestamp 1636915332
transform 1 0 1288 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1636915332
transform 1 0 276 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_9
timestamp 1636915332
transform 1 0 828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1636915332
transform 1 0 0 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1636915332
transform 1 0 1196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _304__4
timestamp 1636915332
transform -1 0 828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__SET_B
timestamp 1636915332
transform 1 0 2392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__456__RESET_B
timestamp 1636915332
transform 1 0 3404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_28
timestamp 1636915332
transform 1 0 2576 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_36
timestamp 1636915332
transform 1 0 3312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1636915332
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtn_1  _456_
timestamp 1636915332
transform 1 0 3680 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__SET_B
timestamp 1636915332
transform 1 0 5796 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_60
timestamp 1636915332
transform 1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1636915332
transform 1 0 5980 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_2  _450_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 6072 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1636915332
transform 1 0 8372 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _368_
timestamp 1636915332
transform 1 0 8004 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _451_
timestamp 1636915332
transform 1 0 8464 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_8_112
timestamp 1636915332
transform 1 0 10304 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_116
timestamp 1636915332
transform 1 0 10672 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_118
timestamp 1636915332
transform 1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1636915332
transform 1 0 10764 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _321_
timestamp 1636915332
transform -1 0 11776 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__RESET_B
timestamp 1636915332
transform 1 0 13524 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_135
timestamp 1636915332
transform 1 0 12420 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_144
timestamp 1636915332
transform 1 0 13248 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1636915332
transform 1 0 13156 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_1  _320_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 11776 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _343_
timestamp 1636915332
transform 1 0 12144 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _476_
timestamp 1636915332
transform -1 0 15548 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__RESET_B
timestamp 1636915332
transform 1 0 15640 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1636915332
transform 1 0 15548 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _438_
timestamp 1636915332
transform -1 0 17940 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_6  FILLER_8_196
timestamp 1636915332
transform 1 0 18032 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1636915332
transform 1 0 17940 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1636915332
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1636915332
transform 1 0 276 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1636915332
transform 1 0 0 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _463_
timestamp 1636915332
transform 1 0 460 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__463__SET_B
timestamp 1636915332
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_29
timestamp 1636915332
transform 1 0 2668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_41
timestamp 1636915332
transform 1 0 3772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_49
timestamp 1636915332
transform 1 0 4508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1636915332
transform 1 0 2392 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _371_
timestamp 1636915332
transform 1 0 3864 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_9_53
timestamp 1636915332
transform 1 0 4876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_65
timestamp 1636915332
transform 1 0 5980 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1636915332
transform 1 0 4784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_77
timestamp 1636915332
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_79
timestamp 1636915332
transform 1 0 7268 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_97
timestamp 1636915332
transform 1 0 8924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1636915332
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _213_
timestamp 1636915332
transform -1 0 9384 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _423_
timestamp 1636915332
transform 1 0 7452 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__RESET_B
timestamp 1636915332
transform 1 0 9660 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_102
timestamp 1636915332
transform 1 0 9384 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1636915332
transform 1 0 9568 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _452_
timestamp 1636915332
transform 1 0 9844 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_9_127
timestamp 1636915332
transform 1 0 11684 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_131
timestamp 1636915332
transform 1 0 12052 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_143
timestamp 1636915332
transform 1 0 13156 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1636915332
transform 1 0 11960 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _383_
timestamp 1636915332
transform 1 0 13248 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__RESET_B
timestamp 1636915332
transform 1 0 14720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_151
timestamp 1636915332
transform 1 0 13892 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_155
timestamp 1636915332
transform 1 0 14260 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_157
timestamp 1636915332
transform 1 0 14444 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1636915332
transform 1 0 14352 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _435_
timestamp 1636915332
transform 1 0 14904 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_9_183
timestamp 1636915332
transform 1 0 16836 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_188
timestamp 1636915332
transform 1 0 17296 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1636915332
transform 1 0 16744 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _378_
timestamp 1636915332
transform 1 0 16928 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_200
timestamp 1636915332
transform 1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1636915332
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_14
timestamp 1636915332
transform 1 0 1288 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_22
timestamp 1636915332
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1636915332
transform 1 0 276 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_9
timestamp 1636915332
transform 1 0 828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1636915332
transform 1 0 0 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1636915332
transform 1 0 1196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _265__3
timestamp 1636915332
transform -1 0 828 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_28
timestamp 1636915332
transform 1 0 2576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1636915332
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_2  _252_
timestamp 1636915332
transform 1 0 3680 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1636915332
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _372_
timestamp 1636915332
transform 1 0 3312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _373_
timestamp 1636915332
transform 1 0 2668 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_10_50
timestamp 1636915332
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_62
timestamp 1636915332
transform 1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1636915332
transform 1 0 5980 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _414_
timestamp 1636915332
transform -1 0 5704 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _424_
timestamp 1636915332
transform 1 0 6072 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_10_88
timestamp 1636915332
transform 1 0 8096 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_92
timestamp 1636915332
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1636915332
transform 1 0 8372 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _211_
timestamp 1636915332
transform 1 0 7544 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 10488 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk_A
timestamp 1636915332
transform 1 0 10488 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_116
timestamp 1636915332
transform 1 0 10672 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_122
timestamp 1636915332
transform 1 0 11224 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1636915332
transform 1 0 10764 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_pll_clk
timestamp 1636915332
transform 1 0 10856 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_131
timestamp 1636915332
transform 1 0 12052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_142
timestamp 1636915332
transform 1 0 13064 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_144
timestamp 1636915332
transform 1 0 13248 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1636915332
transform 1 0 13156 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _207_
timestamp 1636915332
transform 1 0 12236 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _208_
timestamp 1636915332
transform -1 0 12052 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _382_
timestamp 1636915332
transform -1 0 13892 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__SET_B
timestamp 1636915332
transform 1 0 15824 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_151
timestamp 1636915332
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_168
timestamp 1636915332
transform 1 0 15456 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_170
timestamp 1636915332
transform 1 0 15640 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1636915332
transform 1 0 15548 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _379_
timestamp 1636915332
transform 1 0 13984 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _416_
timestamp 1636915332
transform 1 0 14628 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1636915332
transform -1 0 18308 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_196
timestamp 1636915332
transform 1 0 18032 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1636915332
transform 1 0 17940 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _474_
timestamp 1636915332
transform 1 0 16008 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1636915332
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1636915332
transform 1 0 18308 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1636915332
transform 1 0 0 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _266_
timestamp 1636915332
transform -1 0 2392 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _464_
timestamp 1636915332
transform 1 0 276 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__RESET_B
timestamp 1636915332
transform 1 0 2852 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_33
timestamp 1636915332
transform 1 0 3036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_41
timestamp 1636915332
transform 1 0 3772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1636915332
transform 1 0 2392 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _267_
timestamp 1636915332
transform -1 0 2852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _401_
timestamp 1636915332
transform 1 0 3864 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_51
timestamp 1636915332
transform 1 0 4692 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1636915332
transform 1 0 5704 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_74
timestamp 1636915332
transform 1 0 6808 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1636915332
transform 1 0 4784 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _415_
timestamp 1636915332
transform 1 0 4876 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_79
timestamp 1636915332
transform 1 0 7268 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_87
timestamp 1636915332
transform 1 0 8004 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1636915332
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _212_
timestamp 1636915332
transform 1 0 8464 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _215_
timestamp 1636915332
transform -1 0 9476 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _217_
timestamp 1636915332
transform 1 0 8096 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_103
timestamp 1636915332
transform 1 0 9476 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1636915332
transform 1 0 9568 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _473_
timestamp 1636915332
transform 1 0 9660 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__RESET_B
timestamp 1636915332
transform 1 0 11776 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1636915332
transform 1 0 11960 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _475_
timestamp 1636915332
transform 1 0 12052 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__RESET_B
timestamp 1636915332
transform 1 0 14444 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_151
timestamp 1636915332
transform 1 0 13892 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_155
timestamp 1636915332
transform 1 0 14260 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1636915332
transform 1 0 14352 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1636915332
transform 1 0 14628 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _439_
timestamp 1636915332
transform 1 0 14904 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1636915332
transform 1 0 16744 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _209_
timestamp 1636915332
transform 1 0 16836 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _393_
timestamp 1636915332
transform 1 0 17664 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_201
timestamp 1636915332
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1636915332
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1636915332
transform 1 0 1012 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_14
timestamp 1636915332
transform 1 0 1288 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_20
timestamp 1636915332
transform 1 0 1840 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1636915332
transform 1 0 276 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1636915332
transform 1 0 0 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1636915332
transform 1 0 1196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _264_
timestamp 1636915332
transform -1 0 2300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_35
timestamp 1636915332
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_49
timestamp 1636915332
transform 1 0 4508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1636915332
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1636915332
transform -1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _256_
timestamp 1636915332
transform 1 0 2300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _263_
timestamp 1636915332
transform -1 0 3220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1636915332
transform 1 0 3680 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_61
timestamp 1636915332
transform 1 0 5612 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_66
timestamp 1636915332
transform 1 0 6072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_70
timestamp 1636915332
transform 1 0 6440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1636915332
transform 1 0 5980 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _425_
timestamp 1636915332
transform 1 0 6532 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_87
timestamp 1636915332
transform 1 0 8004 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_92
timestamp 1636915332
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_96
timestamp 1636915332
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1636915332
transform 1 0 8372 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _214_
timestamp 1636915332
transform 1 0 8096 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk90
timestamp 1636915332
transform -1 0 10764 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_12_124
timestamp 1636915332
transform 1 0 11408 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1636915332
transform 1 0 10764 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _216_
timestamp 1636915332
transform 1 0 10856 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__SET_B
timestamp 1636915332
transform 1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk90_A
timestamp 1636915332
transform 1 0 11776 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_130
timestamp 1636915332
transform 1 0 11960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_142
timestamp 1636915332
transform 1 0 13064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_144
timestamp 1636915332
transform 1 0 13248 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1636915332
transform 1 0 13156 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1636915332
transform -1 0 11776 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__RESET_B
timestamp 1636915332
transform 1 0 15640 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_168
timestamp 1636915332
transform 1 0 15456 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1636915332
transform 1 0 15548 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_1  _271_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 13800 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1636915332
transform -1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _419_
timestamp 1636915332
transform 1 0 14352 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _442_
timestamp 1636915332
transform 1 0 15824 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1636915332
transform -1 0 18308 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_196
timestamp 1636915332
transform 1 0 18032 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1636915332
transform 1 0 17940 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1636915332
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1636915332
transform 1 0 18308 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1636915332
transform 1 0 0 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1636915332
transform 1 0 0 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1636915332
transform 1 0 276 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1636915332
transform 1 0 1012 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _270_
timestamp 1636915332
transform -1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _269_
timestamp 1636915332
transform -1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1636915332
transform -1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1636915332
transform 1 0 1196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_23
timestamp 1636915332
transform 1 0 2116 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_18
timestamp 1636915332
transform 1 0 1656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_14
timestamp 1636915332
transform 1 0 1288 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtn_1  _462_
timestamp 1636915332
transform 1 0 276 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__462__RESET_B
timestamp 1636915332
transform 1 0 2484 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_38
timestamp 1636915332
transform 1 0 3496 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_37
timestamp 1636915332
transform 1 0 3404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1636915332
transform 1 0 2392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1636915332
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o21bai_1  _259_
timestamp 1636915332
transform -1 0 5060 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _262_
timestamp 1636915332
transform 1 0 2484 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _389_
timestamp 1636915332
transform 1 0 3680 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _390_
timestamp 1636915332
transform 1 0 2668 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_1  _260_
timestamp 1636915332
transform -1 0 5796 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _253_
timestamp 1636915332
transform -1 0 5428 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1636915332
transform 1 0 4784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_53
timestamp 1636915332
transform 1 0 4876 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_50
timestamp 1636915332
transform 1 0 4600 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__SET_B
timestamp 1636915332
transform 1 0 4968 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_pll_clk90
timestamp 1636915332
transform -1 0 7176 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _249__2
timestamp 1636915332
transform -1 0 6348 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1636915332
transform 1 0 5980 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_73
timestamp 1636915332
transform 1 0 6716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_69
timestamp 1636915332
transform 1 0 6348 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_63
timestamp 1636915332
transform 1 0 5796 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_1  _465_
timestamp 1636915332
transform 1 0 5152 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _386_
timestamp 1636915332
transform 1 0 7268 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1636915332
transform -1 0 7544 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1636915332
transform 1 0 7176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_78
timestamp 1636915332
transform 1 0 7176 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_82
timestamp 1636915332
transform 1 0 7544 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_77
timestamp 1636915332
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _221_
timestamp 1636915332
transform -1 0 9016 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1636915332
transform 1 0 8372 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_92
timestamp 1636915332
transform 1 0 8464 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_88
timestamp 1636915332
transform 1 0 8096 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_90
timestamp 1636915332
transform 1 0 8280 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_98
timestamp 1636915332
transform 1 0 9016 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _229_
timestamp 1636915332
transform -1 0 10396 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _226_
timestamp 1636915332
transform 1 0 9292 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1636915332
transform 1 0 9568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_100
timestamp 1636915332
transform 1 0 9200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__RESET_B
timestamp 1636915332
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__SET_B
timestamp 1636915332
transform 1 0 9844 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_pll_clk90
timestamp 1636915332
transform 1 0 11224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _230_
timestamp 1636915332
transform -1 0 10764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1636915332
transform 1 0 10764 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_118
timestamp 1636915332
transform 1 0 10856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _472_
timestamp 1636915332
transform 1 0 10028 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _359_
timestamp 1636915332
transform 1 0 12052 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1636915332
transform 1 0 11960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _276_
timestamp 1636915332
transform 1 0 13156 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _275_
timestamp 1636915332
transform -1 0 13800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1636915332
transform 1 0 12880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1636915332
transform 1 0 13156 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_142
timestamp 1636915332
transform 1 0 13064 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_138
timestamp 1636915332
transform 1 0 12696 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_138
timestamp 1636915332
transform 1 0 12696 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__o2bb2ai_2  _360_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 14352 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_126
timestamp 1636915332
transform 1 0 11592 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__SET_B
timestamp 1636915332
transform 1 0 15364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_165
timestamp 1636915332
transform 1 0 15180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_170
timestamp 1636915332
transform 1 0 15640 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1636915332
transform 1 0 14352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1636915332
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_1  _274_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 13800 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _399_
timestamp 1636915332
transform -1 0 15180 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_4  _443_
timestamp 1636915332
transform 1 0 15732 0 1 7616
box -38 -48 2246 592
use sky130_fd_sc_hd__dfstp_1  _461_
timestamp 1636915332
transform 1 0 14444 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1636915332
transform 1 0 16376 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_186
timestamp 1636915332
transform 1 0 17112 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_198
timestamp 1636915332
transform 1 0 18216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_196
timestamp 1636915332
transform 1 0 18032 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1636915332
transform 1 0 16744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1636915332
transform 1 0 17940 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 1636915332
transform 1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1636915332
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1636915332
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__SET_B
timestamp 1636915332
transform 1 0 2208 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1636915332
transform 1 0 0 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _467_
timestamp 1636915332
transform 1 0 276 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1636915332
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_34
timestamp 1636915332
transform 1 0 3128 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_40
timestamp 1636915332
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_47
timestamp 1636915332
transform 1 0 4324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1636915332
transform 1 0 2392 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o211ai_1  _258_
timestamp 1636915332
transform -1 0 4324 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _261_
timestamp 1636915332
transform 1 0 2852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_51
timestamp 1636915332
transform 1 0 4692 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_61
timestamp 1636915332
transform 1 0 5612 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_69
timestamp 1636915332
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1636915332
transform 1 0 4784 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _218_
timestamp 1636915332
transform -1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _227_
timestamp 1636915332
transform 1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _236_
timestamp 1636915332
transform -1 0 7176 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_83
timestamp 1636915332
transform 1 0 7636 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_98
timestamp 1636915332
transform 1 0 9016 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1636915332
transform 1 0 7176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _235_
timestamp 1636915332
transform -1 0 7636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _374_
timestamp 1636915332
transform -1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _385_
timestamp 1636915332
transform 1 0 7820 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_115
timestamp 1636915332
transform 1 0 10580 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1636915332
transform 1 0 9568 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1636915332
transform -1 0 10304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _224_
timestamp 1636915332
transform -1 0 10028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1636915332
transform 1 0 10304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1636915332
transform 1 0 10672 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__RESET_B
timestamp 1636915332
transform 1 0 12328 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1636915332
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_129
timestamp 1636915332
transform 1 0 11868 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_131
timestamp 1636915332
transform 1 0 12052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1636915332
transform 1 0 11960 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _441_
timestamp 1636915332
transform 1 0 12512 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_15_160
timestamp 1636915332
transform 1 0 14720 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1636915332
transform 1 0 14352 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _358_
timestamp 1636915332
transform -1 0 14720 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _440_
timestamp 1636915332
transform 1 0 14812 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1636915332
transform -1 0 18308 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_183
timestamp 1636915332
transform 1 0 16836 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_195
timestamp 1636915332
transform 1 0 17940 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1636915332
transform 1 0 16744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1636915332
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1636915332
transform 1 0 18308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_14
timestamp 1636915332
transform 1 0 1288 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_18
timestamp 1636915332
transform 1 0 1656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1636915332
transform 1 0 276 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_7
timestamp 1636915332
transform 1 0 644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1636915332
transform 1 0 0 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1636915332
transform 1 0 1196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _245__1
timestamp 1636915332
transform -1 0 644 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _246_
timestamp 1636915332
transform 1 0 1748 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_32
timestamp 1636915332
transform 1 0 2944 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_40
timestamp 1636915332
transform 1 0 3680 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_48
timestamp 1636915332
transform 1 0 4416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1636915332
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1636915332
transform 1 0 3036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1636915332
transform 1 0 2668 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _247_
timestamp 1636915332
transform -1 0 2668 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _250_
timestamp 1636915332
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _257_
timestamp 1636915332
transform 1 0 3312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_57
timestamp 1636915332
transform 1 0 5244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_66
timestamp 1636915332
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1636915332
transform 1 0 5980 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _220_
timestamp 1636915332
transform -1 0 5244 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _228_
timestamp 1636915332
transform 1 0 5612 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _232_
timestamp 1636915332
transform -1 0 6992 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_80
timestamp 1636915332
transform 1 0 7360 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_88
timestamp 1636915332
transform 1 0 8096 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_92
timestamp 1636915332
transform 1 0 8464 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1636915332
transform 1 0 8372 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1636915332
transform 1 0 8740 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _231_
timestamp 1636915332
transform -1 0 7360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _234_
timestamp 1636915332
transform -1 0 9752 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_118
timestamp 1636915332
transform 1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1636915332
transform 1 0 10764 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _233_
timestamp 1636915332
transform -1 0 10120 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _375_
timestamp 1636915332
transform 1 0 10120 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _397_
timestamp 1636915332
transform 1 0 11132 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__RESET_B
timestamp 1636915332
transform 1 0 12144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_130
timestamp 1636915332
transform 1 0 11960 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1636915332
transform 1 0 13156 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1636915332
transform 1 0 12328 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _431_
timestamp 1636915332
transform -1 0 15088 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__SET_B
timestamp 1636915332
transform 1 0 15088 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__RESET_B
timestamp 1636915332
transform 1 0 15640 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_166
timestamp 1636915332
transform 1 0 15272 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1636915332
transform 1 0 15548 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _444_
timestamp 1636915332
transform 1 0 15824 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_6  FILLER_16_196
timestamp 1636915332
transform 1 0 18032 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1636915332
transform 1 0 17940 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1636915332
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1636915332
transform 1 0 0 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _237_
timestamp 1636915332
transform -1 0 2392 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _466_
timestamp 1636915332
transform 1 0 276 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__RESET_B
timestamp 1636915332
transform 1 0 3036 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__RESET_B
timestamp 1636915332
transform 1 0 3496 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_35
timestamp 1636915332
transform 1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1636915332
transform 1 0 2392 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__o21bai_1  _239_
timestamp 1636915332
transform 1 0 2484 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _243_
timestamp 1636915332
transform 1 0 3680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _396_
timestamp 1636915332
transform 1 0 3956 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__RESET_B
timestamp 1636915332
transform 1 0 5152 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1636915332
transform 1 0 4784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1636915332
transform -1 0 5152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _471_
timestamp 1636915332
transform 1 0 5336 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_17_88
timestamp 1636915332
transform 1 0 8096 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_98
timestamp 1636915332
transform 1 0 9016 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1636915332
transform 1 0 7176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _394_
timestamp 1636915332
transform 1 0 8188 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _395_
timestamp 1636915332
transform 1 0 7268 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_112
timestamp 1636915332
transform 1 0 10304 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1636915332
transform 1 0 9568 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _376_
timestamp 1636915332
transform 1 0 9292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _377_
timestamp 1636915332
transform -1 0 10304 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _426_
timestamp 1636915332
transform 1 0 10396 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_ext_clk_A
timestamp 1636915332
transform -1 0 12512 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp 1636915332
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_131
timestamp 1636915332
transform 1 0 12052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1636915332
transform 1 0 11960 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ext_clk
timestamp 1636915332
transform 1 0 12512 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__SET_B
timestamp 1636915332
transform 1 0 14628 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_157
timestamp 1636915332
transform 1 0 14444 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1636915332
transform 1 0 14352 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _428_
timestamp 1636915332
transform 1 0 14812 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_17_183
timestamp 1636915332
transform 1 0 16836 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_195
timestamp 1636915332
transform 1 0 17940 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1636915332
transform 1 0 16744 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_201
timestamp 1636915332
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1636915332
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1636915332
transform -1 0 1472 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_11
timestamp 1636915332
transform 1 0 1012 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1636915332
transform 1 0 276 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1636915332
transform 1 0 0 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1636915332
transform 1 0 1196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_12  input3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1472 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1636915332
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2ai_1  _244_
timestamp 1636915332
transform -1 0 3588 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtn_1  _468_
timestamp 1636915332
transform 1 0 3680 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__RESET_B
timestamp 1636915332
transform 1 0 5796 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_60
timestamp 1636915332
transform 1 0 5520 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1636915332
transform 1 0 5980 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _469_
timestamp 1636915332
transform 1 0 6072 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__SET_B
timestamp 1636915332
transform 1 0 8188 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_87
timestamp 1636915332
transform 1 0 8004 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1636915332
transform 1 0 8372 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _470_
timestamp 1636915332
transform 1 0 8464 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__S
timestamp 1636915332
transform 1 0 11132 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__RESET_B
timestamp 1636915332
transform 1 0 10580 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_113
timestamp 1636915332
transform 1 0 10396 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1636915332
transform 1 0 10764 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _350_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 11132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _432_
timestamp 1636915332
transform 1 0 11316 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1636915332
transform 1 0 13156 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _346__9
timestamp 1636915332
transform 1 0 13248 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _429_
timestamp 1636915332
transform 1 0 13524 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_18_168
timestamp 1636915332
transform 1 0 15456 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_170
timestamp 1636915332
transform 1 0 15640 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1636915332
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _348__7
timestamp 1636915332
transform 1 0 15732 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1636915332
transform -1 0 18308 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_196
timestamp 1636915332
transform 1 0 18032 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1636915332
transform 1 0 17940 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _427_
timestamp 1636915332
transform 1 0 16008 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1636915332
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1636915332
transform 1 0 18308 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1636915332
transform 1 0 1012 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_14
timestamp 1636915332
transform 1 0 1288 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1636915332
transform 1 0 276 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1636915332
transform 1 0 0 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1636915332
transform 1 0 1196 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1636915332
transform -1 0 2392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _248_
timestamp 1636915332
transform -1 0 2116 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_33
timestamp 1636915332
transform 1 0 3036 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_40
timestamp 1636915332
transform 1 0 3680 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1636915332
transform 1 0 2392 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1636915332
transform 1 0 3588 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _240_
timestamp 1636915332
transform 1 0 2484 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_53
timestamp 1636915332
transform 1 0 4876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_66
timestamp 1636915332
transform 1 0 6072 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1636915332
transform 1 0 4784 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1636915332
transform 1 0 5980 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_82
timestamp 1636915332
transform 1 0 7544 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_90
timestamp 1636915332
transform 1 0 8280 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_92
timestamp 1636915332
transform 1 0 8464 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1636915332
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1636915332
transform 1 0 8372 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  output10
timestamp 1636915332
transform 1 0 7268 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_105
timestamp 1636915332
transform 1 0 9660 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_116
timestamp 1636915332
transform 1 0 10672 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_118
timestamp 1636915332
transform 1 0 10856 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1636915332
transform 1 0 9568 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1636915332
transform 1 0 10764 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _349_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10948 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_ext_clk
timestamp 1636915332
transform 1 0 10028 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output12
timestamp 1636915332
transform 1 0 10396 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1636915332
transform 1 0 11776 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1636915332
transform 1 0 11960 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1636915332
transform 1 0 13156 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _418_
timestamp 1636915332
transform -1 0 14076 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 12052 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1636915332
transform -1 0 13156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__SET_B
timestamp 1636915332
transform 1 0 14076 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _384__13 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 14720 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1636915332
transform 1 0 14352 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_155
timestamp 1636915332
transform 1 0 14260 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _347__8
timestamp 1636915332
transform -1 0 15180 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1636915332
transform 1 0 14720 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_ext_clk
timestamp 1636915332
transform -1 0 15548 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1636915332
transform 1 0 15548 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_170
timestamp 1636915332
transform 1 0 15640 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__SET_B
timestamp 1636915332
transform 1 0 15824 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1636915332
transform -1 0 17940 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_174
timestamp 1636915332
transform 1 0 16008 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_183
timestamp 1636915332
transform 1 0 16836 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_191
timestamp 1636915332
transform 1 0 17572 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1636915332
transform 1 0 16744 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1636915332
transform 1 0 17940 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _381_
timestamp 1636915332
transform 1 0 18032 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1636915332
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1636915332
transform 1 0 18308 0 -1 10880
box -38 -48 314 592
<< labels >>
rlabel metal5 s 0 4812 18860 5132 6 VGND
port 0 nsew ground input
rlabel metal5 s 0 8192 18860 8512 6 VGND
port 0 nsew ground input
rlabel metal4 s 4654 -48 4974 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 7754 -48 8074 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 10854 -48 11174 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 13954 -48 14274 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 17054 -48 17374 10928 6 VGND
port 0 nsew ground input
rlabel metal5 s 0 3122 18860 3442 6 VPWR
port 1 nsew power input
rlabel metal5 s 0 6502 18860 6822 6 VPWR
port 1 nsew power input
rlabel metal5 s 0 9882 18860 10202 6 VPWR
port 1 nsew power input
rlabel metal4 s 3104 -48 3424 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 6204 -48 6524 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 9304 -48 9624 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 12404 -48 12724 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 15504 -48 15824 10928 6 VPWR
port 1 nsew power input
rlabel metal2 s 7102 11200 7158 12000 6 core_clk
port 2 nsew signal tristate
rlabel metal2 s 4250 11200 4306 12000 6 ext_clk
port 3 nsew signal input
rlabel metal3 s 19200 688 20000 808 6 ext_clk_sel
port 4 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 ext_reset
port 5 nsew signal input
rlabel metal2 s 15658 11200 15714 12000 6 pll_clk
port 6 nsew signal input
rlabel metal2 s 18510 11200 18566 12000 6 pll_clk90
port 7 nsew signal input
rlabel metal2 s 1398 11200 1454 12000 6 resetb
port 8 nsew signal input
rlabel metal2 s 12806 11200 12862 12000 6 resetb_sync
port 9 nsew signal tristate
rlabel metal3 s 19200 6672 20000 6792 6 sel2[0]
port 10 nsew signal input
rlabel metal3 s 19200 8168 20000 8288 6 sel2[1]
port 11 nsew signal input
rlabel metal3 s 19200 9664 20000 9784 6 sel2[2]
port 12 nsew signal input
rlabel metal3 s 19200 2184 20000 2304 6 sel[0]
port 13 nsew signal input
rlabel metal3 s 19200 3680 20000 3800 6 sel[1]
port 14 nsew signal input
rlabel metal3 s 19200 5176 20000 5296 6 sel[2]
port 15 nsew signal input
rlabel metal2 s 9954 11200 10010 12000 6 user_clk
port 16 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 12000
<< end >>
