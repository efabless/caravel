magic
tech sky130A
timestamp 0
<< properties >>
string FIXED_BBOX 0 0 0 0
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 264461246
string GDS_FILE /home/hosni/caravan/caravel/openlane/caravan_core/runs/23_05_29_20_16/results/signoff/caravan_core.magic.gds
string GDS_START 62452652
<< end >>

