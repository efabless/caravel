* NGSPICE file created from mgmt_protect.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=5.36e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VNB VPB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VNB VPB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_2 Y A VPWR VGND VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_2 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__einvp_8 A Z TE VPWR VGND VNB VPB
X0 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X1 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X4 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X8 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X9 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X21 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X26 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X30 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X32 VPWR TE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VGND TE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_4 Y A B VGND VPWR VNB VPB
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_1 Y B A VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_12 A Y VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A X VGND VPWR VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_12 A X VGND VPWR VNB VPB
X0 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND A X VNB VPB
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 X A VGND VPWR VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_8 A Y VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_8 Y A VGND VPWR VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_8 A X VGND VPWR VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VNB VPB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_6 Y A VPWR VGND VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_4 Y A VPWR VGND VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_2 Y A B VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_8 A B Y VGND VPWR VNB VPB
X0 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2b_2 VPWR VGND X B A_N VNB VPB
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_16 Y A VGND VPWR VNB VPB
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt mprj2_logic_high HI vccd2 vssd2
XFILLER_0_57 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_209 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_69 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_81 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_181 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_29 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_193 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_95 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XPHY_0 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_1 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_85 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_1_41 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_53 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_2 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_3 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_141 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_197 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_153 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_165 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_209 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_113 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_69 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_169 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_125 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_15 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_181 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_137 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_193 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_29 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_107 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_197 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_153 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_165 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_113 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_3 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_169 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_125 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_137 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_81 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
Xinst inst/LO HI vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__conb_1
XFILLER_0_85 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_41 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_109 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_97 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_53 vccd2 vssd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
.ends

.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295] HI[296]
+ HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304] HI[305]
+ HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314] HI[315]
+ HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324] HI[325]
+ HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334] HI[335]
+ HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344] HI[345]
+ HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354] HI[355]
+ HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364] HI[365]
+ HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374] HI[375]
+ HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384] HI[385]
+ HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394] HI[395]
+ HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403] HI[404]
+ HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413] HI[414]
+ HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423] HI[424]
+ HI[425] HI[426] HI[427] HI[428] HI[42] HI[430] HI[431] HI[432] HI[433] HI[434] HI[435]
+ HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443] HI[444] HI[445]
+ HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453] HI[454] HI[455]
+ HI[456] HI[457] HI[458] HI[459] HI[45] HI[460] HI[461] HI[462] HI[46] HI[47] HI[48]
+ HI[49] HI[4] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57] HI[58] HI[59]
+ HI[5] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68] HI[69] HI[6]
+ HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79] HI[7] HI[80]
+ HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8] HI[90] HI[91]
+ HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1 HI[287] HI[429]
+ vssd1
Xinsts\[210\] insts\[210\]/LO HI[210] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[308\] insts\[308\]/LO HI[308] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[425\] insts\[425\]/LO HI[425] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[160\] insts\[160\]/LO HI[160] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_357 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_302 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[258\] insts\[258\]/LO HI[258] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[40\] insts\[40\]/LO HI[40] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[375\] insts\[375\]/LO HI[375] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[88\] insts\[88\]/LO HI[88] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_165 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[123\] insts\[123\]/LO HI[123] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_0_669 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[338\] insts\[338\]/LO HI[338] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[240\] insts\[240\]/LO HI[240] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[9\] insts\[9\]/LO HI[9] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[455\] insts\[455\]/LO HI[455] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[288\] insts\[288\]/LO HI[288] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[190\] insts\[190\]/LO HI[190] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[70\] insts\[70\]/LO HI[70] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[203\] insts\[203\]/LO HI[203] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_561 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[418\] insts\[418\]/LO HI[418] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[153\] insts\[153\]/LO HI[153] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[320\] insts\[320\]/LO HI[320] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[33\] insts\[33\]/LO HI[33] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[368\] insts\[368\]/LO HI[368] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[270\] insts\[270\]/LO HI[270] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_177 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_486 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[116\] insts\[116\]/LO HI[116] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[400\] insts\[400\]/LO HI[400] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[233\] insts\[233\]/LO HI[233] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[183\] insts\[183\]/LO HI[183] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[350\] insts\[350\]/LO HI[350] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[448\] insts\[448\]/LO HI[448] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_721 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[63\] insts\[63\]/LO HI[63] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[398\] insts\[398\]/LO HI[398] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_573 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[146\] insts\[146\]/LO HI[146] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[313\] insts\[313\]/LO HI[313] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[26\] insts\[26\]/LO HI[26] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_3_3 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[430\] insts\[430\]/LO HI[430] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_189 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[263\] insts\[263\]/LO HI[263] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[380\] insts\[380\]/LO HI[380] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[109\] insts\[109\]/LO HI[109] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[93\] insts\[93\]/LO HI[93] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_3_498 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_80 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[226\] insts\[226\]/LO HI[226] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[343\] insts\[343\]/LO HI[343] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[176\] insts\[176\]/LO HI[176] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[56\] insts\[56\]/LO HI[56] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[460\] insts\[460\]/LO HI[460] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[293\] insts\[293\]/LO HI[293] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_541 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_585 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[139\] insts\[139\]/LO HI[139] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[306\] insts\[306\]/LO HI[306] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[19\] insts\[19\]/LO HI[19] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_393 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[423\] insts\[423\]/LO HI[423] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[256\] insts\[256\]/LO HI[256] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[373\] insts\[373\]/LO HI[373] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_0_617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[86\] insts\[86\]/LO HI[86] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[121\] insts\[121\]/LO HI[121] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[219\] insts\[219\]/LO HI[219] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[336\] insts\[336\]/LO HI[336] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[169\] insts\[169\]/LO HI[169] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[49\] insts\[49\]/LO HI[49] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[286\] insts\[286\]/LO HI[286] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[7\] insts\[7\]/LO HI[7] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[453\] insts\[453\]/LO HI[453] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_597 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[201\] insts\[201\]/LO HI[201] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[416\] insts\[416\]/LO HI[416] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[249\] insts\[249\]/LO HI[249] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[151\] insts\[151\]/LO HI[151] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_681 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[31\] insts\[31\]/LO HI[31] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_0_629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[366\] insts\[366\]/LO HI[366] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[199\] insts\[199\]/LO HI[199] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[79\] insts\[79\]/LO HI[79] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[114\] insts\[114\]/LO HI[114] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[329\] insts\[329\]/LO HI[329] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[231\] insts\[231\]/LO HI[231] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[446\] insts\[446\]/LO HI[446] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[181\] insts\[181\]/LO HI[181] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[279\] insts\[279\]/LO HI[279] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[61\] insts\[61\]/LO HI[61] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[396\] insts\[396\]/LO HI[396] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[144\] insts\[144\]/LO HI[144] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[409\] insts\[409\]/LO HI[409] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[311\] insts\[311\]/LO HI[311] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[24\] insts\[24\]/LO HI[24] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[359\] insts\[359\]/LO HI[359] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[261\] insts\[261\]/LO HI[261] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[107\] insts\[107\]/LO HI[107] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[91\] insts\[91\]/LO HI[91] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[224\] insts\[224\]/LO HI[224] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XPHY_0 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[439\] insts\[439\]/LO HI[439] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[174\] insts\[174\]/LO HI[174] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[341\] insts\[341\]/LO HI[341] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[54\] insts\[54\]/LO HI[54] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[389\] insts\[389\]/LO HI[389] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[291\] insts\[291\]/LO HI[291] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[137\] insts\[137\]/LO HI[137] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[304\] insts\[304\]/LO HI[304] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[17\] insts\[17\]/LO HI[17] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[421\] insts\[421\]/LO HI[421] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[254\] insts\[254\]/LO HI[254] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[371\] insts\[371\]/LO HI[371] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[84\] insts\[84\]/LO HI[84] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[217\] insts\[217\]/LO HI[217] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XPHY_1 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[334\] insts\[334\]/LO HI[334] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[167\] insts\[167\]/LO HI[167] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[47\] insts\[47\]/LO HI[47] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_309 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[5\] insts\[5\]/LO HI[5] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[451\] insts\[451\]/LO HI[451] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[284\] insts\[284\]/LO HI[284] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_331 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_172 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[247\] insts\[247\]/LO HI[247] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[414\] insts\[414\]/LO HI[414] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_470 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_96 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[364\] insts\[364\]/LO HI[364] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[197\] insts\[197\]/LO HI[197] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[77\] insts\[77\]/LO HI[77] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[112\] insts\[112\]/LO HI[112] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XPHY_2 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[327\] insts\[327\]/LO HI[327] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_557 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[444\] insts\[444\]/LO HI[444] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[277\] insts\[277\]/LO HI[277] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_343 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[394\] insts\[394\]/LO HI[394] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_118 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_184 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[407\] insts\[407\]/LO HI[407] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[142\] insts\[142\]/LO HI[142] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[22\] insts\[22\]/LO HI[22] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[357\] insts\[357\]/LO HI[357] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[105\] insts\[105\]/LO HI[105] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XPHY_3 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[222\] insts\[222\]/LO HI[222] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[437\] insts\[437\]/LO HI[437] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[172\] insts\[172\]/LO HI[172] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_355 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[52\] insts\[52\]/LO HI[52] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[387\] insts\[387\]/LO HI[387] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_196 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[135\] insts\[135\]/LO HI[135] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[302\] insts\[302\]/LO HI[302] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[15\] insts\[15\]/LO HI[15] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[252\] insts\[252\]/LO HI[252] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[82\] insts\[82\]/LO HI[82] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XPHY_4 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[215\] insts\[215\]/LO HI[215] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[165\] insts\[165\]/LO HI[165] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[332\] insts\[332\]/LO HI[332] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_301 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_367 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[45\] insts\[45\]/LO HI[45] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_109 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[3\] insts\[3\]/LO HI[3] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_142 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[282\] insts\[282\]/LO HI[282] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[128\] insts\[128\]/LO HI[128] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[412\] insts\[412\]/LO HI[412] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[245\] insts\[245\]/LO HI[245] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[362\] insts\[362\]/LO HI[362] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[195\] insts\[195\]/LO HI[195] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[75\] insts\[75\]/LO HI[75] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XPHY_5 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[110\] insts\[110\]/LO HI[110] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[208\] insts\[208\]/LO HI[208] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_505 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[158\] insts\[158\]/LO HI[158] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[325\] insts\[325\]/LO HI[325] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_379 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[38\] insts\[38\]/LO HI[38] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[442\] insts\[442\]/LO HI[442] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[275\] insts\[275\]/LO HI[275] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_154 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_121 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[392\] insts\[392\]/LO HI[392] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[405\] insts\[405\]/LO HI[405] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[140\] insts\[140\]/LO HI[140] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[238\] insts\[238\]/LO HI[238] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[20\] insts\[20\]/LO HI[20] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[355\] insts\[355\]/LO HI[355] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[188\] insts\[188\]/LO HI[188] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_709 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[68\] insts\[68\]/LO HI[68] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_517 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[103\] insts\[103\]/LO HI[103] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[318\] insts\[318\]/LO HI[318] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[220\] insts\[220\]/LO HI[220] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[170\] insts\[170\]/LO HI[170] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[435\] insts\[435\]/LO HI[435] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_689 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_133 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[268\] insts\[268\]/LO HI[268] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[50\] insts\[50\]/LO HI[50] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[385\] insts\[385\]/LO HI[385] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[98\] insts\[98\]/LO HI[98] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_442 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_68 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[133\] insts\[133\]/LO HI[133] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[300\] insts\[300\]/LO HI[300] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[13\] insts\[13\]/LO HI[13] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XPHY_7 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[348\] insts\[348\]/LO HI[348] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[250\] insts\[250\]/LO HI[250] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[298\] insts\[298\]/LO HI[298] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_529 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[80\] insts\[80\]/LO HI[80] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[213\] insts\[213\]/LO HI[213] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_337 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[428\] insts\[428\]/LO HI[428] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[330\] insts\[330\]/LO HI[330] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[163\] insts\[163\]/LO HI[163] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[43\] insts\[43\]/LO HI[43] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[378\] insts\[378\]/LO HI[378] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[280\] insts\[280\]/LO HI[280] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[1\] insts\[1\]/LO HI[1] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_454 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_421 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_410 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[126\] insts\[126\]/LO HI[126] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[410\] insts\[410\]/LO HI[410] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[243\] insts\[243\]/LO HI[243] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[458\] insts\[458\]/LO HI[458] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[360\] insts\[360\]/LO HI[360] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[193\] insts\[193\]/LO HI[193] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[73\] insts\[73\]/LO HI[73] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[206\] insts\[206\]/LO HI[206] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_625 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_113 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[156\] insts\[156\]/LO HI[156] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[323\] insts\[323\]/LO HI[323] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[36\] insts\[36\]/LO HI[36] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[273\] insts\[273\]/LO HI[273] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[440\] insts\[440\]/LO HI[440] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_433 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[390\] insts\[390\]/LO HI[390] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[119\] insts\[119\]/LO HI[119] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[403\] insts\[403\]/LO HI[403] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[236\] insts\[236\]/LO HI[236] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_0_701 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[353\] insts\[353\]/LO HI[353] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[186\] insts\[186\]/LO HI[186] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[66\] insts\[66\]/LO HI[66] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[101\] insts\[101\]/LO HI[101] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[149\] insts\[149\]/LO HI[149] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_637 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[316\] insts\[316\]/LO HI[316] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[29\] insts\[29\]/LO HI[29] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[433\] insts\[433\]/LO HI[433] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[266\] insts\[266\]/LO HI[266] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[383\] insts\[383\]/LO HI[383] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[96\] insts\[96\]/LO HI[96] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_253 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[131\] insts\[131\]/LO HI[131] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[229\] insts\[229\]/LO HI[229] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_0_713 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[11\] insts\[11\]/LO HI[11] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[346\] insts\[346\]/LO HI[346] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[179\] insts\[179\]/LO HI[179] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[59\] insts\[59\]/LO HI[59] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_307 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[296\] insts\[296\]/LO HI[296] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[309\] insts\[309\]/LO HI[309] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[211\] insts\[211\]/LO HI[211] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[426\] insts\[426\]/LO HI[426] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[161\] insts\[161\]/LO HI[161] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[259\] insts\[259\]/LO HI[259] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[41\] insts\[41\]/LO HI[41] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_490 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_722 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[376\] insts\[376\]/LO HI[376] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_265 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[89\] insts\[89\]/LO HI[89] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_60 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[124\] insts\[124\]/LO HI[124] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_0_725 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[241\] insts\[241\]/LO HI[241] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[339\] insts\[339\]/LO HI[339] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_319 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[456\] insts\[456\]/LO HI[456] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[289\] insts\[289\]/LO HI[289] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[191\] insts\[191\]/LO HI[191] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[71\] insts\[71\]/LO HI[71] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[204\] insts\[204\]/LO HI[204] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[419\] insts\[419\]/LO HI[419] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[154\] insts\[154\]/LO HI[154] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[321\] insts\[321\]/LO HI[321] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[34\] insts\[34\]/LO HI[34] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[369\] insts\[369\]/LO HI[369] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_277 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_233 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[271\] insts\[271\]/LO HI[271] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_72 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[117\] insts\[117\]/LO HI[117] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[234\] insts\[234\]/LO HI[234] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[401\] insts\[401\]/LO HI[401] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[351\] insts\[351\]/LO HI[351] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[449\] insts\[449\]/LO HI[449] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[184\] insts\[184\]/LO HI[184] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[64\] insts\[64\]/LO HI[64] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[399\] insts\[399\]/LO HI[399] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[147\] insts\[147\]/LO HI[147] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[314\] insts\[314\]/LO HI[314] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[27\] insts\[27\]/LO HI[27] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[431\] insts\[431\]/LO HI[431] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_289 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_245 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[264\] insts\[264\]/LO HI[264] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[381\] insts\[381\]/LO HI[381] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[94\] insts\[94\]/LO HI[94] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[227\] insts\[227\]/LO HI[227] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[344\] insts\[344\]/LO HI[344] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[177\] insts\[177\]/LO HI[177] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[57\] insts\[57\]/LO HI[57] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[461\] insts\[461\]/LO HI[461] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[294\] insts\[294\]/LO HI[294] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[307\] insts\[307\]/LO HI[307] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_471 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[424\] insts\[424\]/LO HI[424] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[257\] insts\[257\]/LO HI[257] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_85 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_511 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[374\] insts\[374\]/LO HI[374] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[87\] insts\[87\]/LO HI[87] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[122\] insts\[122\]/LO HI[122] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[337\] insts\[337\]/LO HI[337] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_108 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[8\] insts\[8\]/LO HI[8] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[454\] insts\[454\]/LO HI[454] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[287\] insts\[287\]/LO HI[287] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_653 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[202\] insts\[202\]/LO HI[202] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_461 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[417\] insts\[417\]/LO HI[417] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[152\] insts\[152\]/LO HI[152] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_97 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[32\] insts\[32\]/LO HI[32] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[367\] insts\[367\]/LO HI[367] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[115\] insts\[115\]/LO HI[115] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[232\] insts\[232\]/LO HI[232] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[447\] insts\[447\]/LO HI[447] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[182\] insts\[182\]/LO HI[182] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[62\] insts\[62\]/LO HI[62] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_665 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[397\] insts\[397\]/LO HI[397] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_484 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[145\] insts\[145\]/LO HI[145] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[312\] insts\[312\]/LO HI[312] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[25\] insts\[25\]/LO HI[25] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_281 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[262\] insts\[262\]/LO HI[262] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_3 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[108\] insts\[108\]/LO HI[108] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[92\] insts\[92\]/LO HI[92] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[225\] insts\[225\]/LO HI[225] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[342\] insts\[342\]/LO HI[342] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[175\] insts\[175\]/LO HI[175] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[55\] insts\[55\]/LO HI[55] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[292\] insts\[292\]/LO HI[292] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_441 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[138\] insts\[138\]/LO HI[138] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[305\] insts\[305\]/LO HI[305] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[18\] insts\[18\]/LO HI[18] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_293 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[422\] insts\[422\]/LO HI[422] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[255\] insts\[255\]/LO HI[255] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[372\] insts\[372\]/LO HI[372] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[85\] insts\[85\]/LO HI[85] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[120\] insts\[120\]/LO HI[120] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[218\] insts\[218\]/LO HI[218] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[335\] insts\[335\]/LO HI[335] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[168\] insts\[168\]/LO HI[168] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[48\] insts\[48\]/LO HI[48] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[6\] insts\[6\]/LO HI[6] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[452\] insts\[452\]/LO HI[452] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[285\] insts\[285\]/LO HI[285] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[200\] insts\[200\]/LO HI[200] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_261 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[415\] insts\[415\]/LO HI[415] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[150\] insts\[150\]/LO HI[150] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[248\] insts\[248\]/LO HI[248] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_581 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[30\] insts\[30\]/LO HI[30] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[365\] insts\[365\]/LO HI[365] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[198\] insts\[198\]/LO HI[198] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[78\] insts\[78\]/LO HI[78] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[113\] insts\[113\]/LO HI[113] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[230\] insts\[230\]/LO HI[230] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[328\] insts\[328\]/LO HI[328] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[445\] insts\[445\]/LO HI[445] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[278\] insts\[278\]/LO HI[278] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[180\] insts\[180\]/LO HI[180] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[60\] insts\[60\]/LO HI[60] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[395\] insts\[395\]/LO HI[395] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_273 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[408\] insts\[408\]/LO HI[408] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[143\] insts\[143\]/LO HI[143] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[310\] insts\[310\]/LO HI[310] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[23\] insts\[23\]/LO HI[23] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[358\] insts\[358\]/LO HI[358] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[260\] insts\[260\]/LO HI[260] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[106\] insts\[106\]/LO HI[106] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[90\] insts\[90\]/LO HI[90] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[223\] insts\[223\]/LO HI[223] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[438\] insts\[438\]/LO HI[438] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[340\] insts\[340\]/LO HI[340] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[173\] insts\[173\]/LO HI[173] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[53\] insts\[53\]/LO HI[53] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[388\] insts\[388\]/LO HI[388] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[290\] insts\[290\]/LO HI[290] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_230 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[136\] insts\[136\]/LO HI[136] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[303\] insts\[303\]/LO HI[303] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[16\] insts\[16\]/LO HI[16] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[420\] insts\[420\]/LO HI[420] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[253\] insts\[253\]/LO HI[253] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[370\] insts\[370\]/LO HI[370] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[83\] insts\[83\]/LO HI[83] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[216\] insts\[216\]/LO HI[216] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[166\] insts\[166\]/LO HI[166] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[333\] insts\[333\]/LO HI[333] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[46\] insts\[46\]/LO HI[46] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[450\] insts\[450\]/LO HI[450] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[283\] insts\[283\]/LO HI[283] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[4\] insts\[4\]/LO HI[4] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_710 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_242 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[129\] insts\[129\]/LO HI[129] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[413\] insts\[413\]/LO HI[413] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[246\] insts\[246\]/LO HI[246] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[196\] insts\[196\]/LO HI[196] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[363\] insts\[363\]/LO HI[363] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[76\] insts\[76\]/LO HI[76] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[209\] insts\[209\]/LO HI[209] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[111\] insts\[111\]/LO HI[111] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[159\] insts\[159\]/LO HI[159] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[326\] insts\[326\]/LO HI[326] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[39\] insts\[39\]/LO HI[39] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_722 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[443\] insts\[443\]/LO HI[443] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_221 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_254 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[276\] insts\[276\]/LO HI[276] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[393\] insts\[393\]/LO HI[393] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[406\] insts\[406\]/LO HI[406] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[141\] insts\[141\]/LO HI[141] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[239\] insts\[239\]/LO HI[239] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[21\] insts\[21\]/LO HI[21] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[356\] insts\[356\]/LO HI[356] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[189\] insts\[189\]/LO HI[189] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[69\] insts\[69\]/LO HI[69] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[104\] insts\[104\]/LO HI[104] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[221\] insts\[221\]/LO HI[221] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[319\] insts\[319\]/LO HI[319] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[436\] insts\[436\]/LO HI[436] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[171\] insts\[171\]/LO HI[171] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[269\] insts\[269\]/LO HI[269] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[51\] insts\[51\]/LO HI[51] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[386\] insts\[386\]/LO HI[386] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[99\] insts\[99\]/LO HI[99] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[134\] insts\[134\]/LO HI[134] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[301\] insts\[301\]/LO HI[301] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[14\] insts\[14\]/LO HI[14] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[349\] insts\[349\]/LO HI[349] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[251\] insts\[251\]/LO HI[251] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[299\] insts\[299\]/LO HI[299] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[81\] insts\[81\]/LO HI[81] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[214\] insts\[214\]/LO HI[214] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[429\] insts\[429\]/LO HI[429] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[164\] insts\[164\]/LO HI[164] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[331\] insts\[331\]/LO HI[331] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[44\] insts\[44\]/LO HI[44] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[379\] insts\[379\]/LO HI[379] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[2\] insts\[2\]/LO HI[2] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[281\] insts\[281\]/LO HI[281] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[127\] insts\[127\]/LO HI[127] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[411\] insts\[411\]/LO HI[411] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[244\] insts\[244\]/LO HI[244] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[459\] insts\[459\]/LO HI[459] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[361\] insts\[361\]/LO HI[361] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[194\] insts\[194\]/LO HI[194] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_0_641 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[74\] insts\[74\]/LO HI[74] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_405 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_449 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[207\] insts\[207\]/LO HI[207] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[157\] insts\[157\]/LO HI[157] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[324\] insts\[324\]/LO HI[324] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[37\] insts\[37\]/LO HI[37] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[441\] insts\[441\]/LO HI[441] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_533 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[274\] insts\[274\]/LO HI[274] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[391\] insts\[391\]/LO HI[391] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[404\] insts\[404\]/LO HI[404] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[237\] insts\[237\]/LO HI[237] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_609 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[354\] insts\[354\]/LO HI[354] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[187\] insts\[187\]/LO HI[187] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[67\] insts\[67\]/LO HI[67] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_0_697 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[102\] insts\[102\]/LO HI[102] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_417 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[317\] insts\[317\]/LO HI[317] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[434\] insts\[434\]/LO HI[434] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_545 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[267\] insts\[267\]/LO HI[267] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_589 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[384\] insts\[384\]/LO HI[384] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_386 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[97\] insts\[97\]/LO HI[97] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[132\] insts\[132\]/LO HI[132] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[12\] insts\[12\]/LO HI[12] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[347\] insts\[347\]/LO HI[347] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_1_429 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[297\] insts\[297\]/LO HI[297] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[212\] insts\[212\]/LO HI[212] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[162\] insts\[162\]/LO HI[162] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[427\] insts\[427\]/LO HI[427] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_502 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[42\] insts\[42\]/LO HI[42] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[377\] insts\[377\]/LO HI[377] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_398 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_365 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_321 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[0\] insts\[0\]/LO HI[0] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[125\] insts\[125\]/LO HI[125] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[242\] insts\[242\]/LO HI[242] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[457\] insts\[457\]/LO HI[457] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[192\] insts\[192\]/LO HI[192] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[72\] insts\[72\]/LO HI[72] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[205\] insts\[205\]/LO HI[205] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_569 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_514 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[155\] insts\[155\]/LO HI[155] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[322\] insts\[322\]/LO HI[322] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[35\] insts\[35\]/LO HI[35] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[272\] insts\[272\]/LO HI[272] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_377 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_333 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[118\] insts\[118\]/LO HI[118] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_141 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_130 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[402\] insts\[402\]/LO HI[402] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[235\] insts\[235\]/LO HI[235] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_0_601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[352\] insts\[352\]/LO HI[352] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[185\] insts\[185\]/LO HI[185] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[65\] insts\[65\]/LO HI[65] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[100\] insts\[100\]/LO HI[100] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[148\] insts\[148\]/LO HI[148] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_526 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[315\] insts\[315\]/LO HI[315] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[28\] insts\[28\]/LO HI[28] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[265\] insts\[265\]/LO HI[265] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[432\] insts\[432\]/LO HI[432] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_345 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[382\] insts\[382\]/LO HI[382] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_2_197 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_153 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[95\] insts\[95\]/LO HI[95] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[130\] insts\[130\]/LO HI[130] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[228\] insts\[228\]/LO HI[228] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
XFILLER_0_613 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[10\] insts\[10\]/LO HI[10] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[178\] insts\[178\]/LO HI[178] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[345\] insts\[345\]/LO HI[345] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[58\] insts\[58\]/LO HI[58] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[462\] insts\[462\]/LO HI[462] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xinsts\[295\] insts\[295\]/LO HI[295] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
.ends

.subckt sky130_fd_sc_hd__inv_16 Y A VGND VPWR VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hvl__conb_1 VGND VNB VPWR VPB LO HI
R0 VGND LO sky130_fd_pr__res_generic_po w=510000u l=45000u
R1 HI VPWR sky130_fd_pr__res_generic_po w=510000u l=45000u
.ends

.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 X A VPWR VGND VNB VPB LVPWR
X0 a_30_1337# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X1 VGND a_30_1337# a_30_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X2 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X5 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X6 VGND A a_30_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X7 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X8 a_389_141# a_30_207# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X9 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X10 LVPWR a_389_141# X LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 VGND a_389_141# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X12 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X13 LVPWR a_389_1337# a_389_141# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 a_30_207# a_30_1337# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X15 a_389_1337# a_389_141# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt mgmt_protect_hv mprj2_vdd_logic1 mprj_vdd_logic1 vccd vssd vdda1 vdda2 dw_6116_1496#
+ vssa1 dw_13698_1476# vssa2
Xmprj2_logic_high_hvl vssa2 vssa2 vdda2 vdda2 mprj2_logic_high_hvl/LO mprj2_logic_high_lv/A
+ sky130_fd_sc_hvl__conb_1
Xmprj_logic_high_hvl vssa1 vssa1 vdda1 vdda1 mprj_logic_high_hvl/LO mprj_logic_high_lv/A
+ sky130_fd_sc_hvl__conb_1
Xmprj_logic_high_lv mprj_vdd_logic1 mprj_logic_high_lv/A vdda1 vssd vssd vdda1 vccd
+ sky130_fd_sc_hvl__lsbufhv2lv_1
Xmprj2_logic_high_lv mprj2_vdd_logic1 mprj2_logic_high_lv/A vdda2 vssd vssd vdda2
+ vccd sky130_fd_sc_hvl__lsbufhv2lv_1
.ends

.subckt sky130_fd_sc_hd__and2_4 X B A VGND VPWR VNB VPB
X0 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND B a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 X A VGND VPWR VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 X A VGND VPWR VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102]
+ la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107]
+ la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[10] la_iena_mprj[110] la_iena_mprj[111]
+ la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116]
+ la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[11] la_iena_mprj[120]
+ la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125]
+ la_iena_mprj[126] la_iena_mprj[127] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14]
+ la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19]
+ la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23]
+ la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28]
+ la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32]
+ la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37]
+ la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3] la_iena_mprj[40] la_iena_mprj[41]
+ la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46]
+ la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[4] la_iena_mprj[50]
+ la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55]
+ la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[5]
+ la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64]
+ la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69]
+ la_iena_mprj[6] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73]
+ la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78]
+ la_iena_mprj[79] la_iena_mprj[7] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82]
+ la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87]
+ la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[8] la_iena_mprj[90] la_iena_mprj[91]
+ la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96]
+ la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[9] la_oenb_core[0]
+ la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104]
+ la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109]
+ la_oenb_core[10] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113]
+ la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118]
+ la_oenb_core[119] la_oenb_core[11] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122]
+ la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127]
+ la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16]
+ la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[1] la_oenb_core[20]
+ la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25]
+ la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[2]
+ la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34]
+ la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39]
+ la_oenb_core[3] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43]
+ la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48]
+ la_oenb_core[49] la_oenb_core[4] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52]
+ la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57]
+ la_oenb_core[58] la_oenb_core[59] la_oenb_core[5] la_oenb_core[60] la_oenb_core[61]
+ la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66]
+ la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[6] la_oenb_core[70]
+ la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75]
+ la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[7]
+ la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84]
+ la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89]
+ la_oenb_core[8] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93]
+ la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98]
+ la_oenb_core[99] la_oenb_core[9] la_oenb_mprj[0] la_oenb_mprj[100] la_oenb_mprj[101]
+ la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106]
+ la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[10] la_oenb_mprj[110]
+ la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115]
+ la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[11]
+ la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124]
+ la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] la_oenb_mprj[12] la_oenb_mprj[13]
+ la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18]
+ la_oenb_mprj[19] la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22]
+ la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27]
+ la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31]
+ la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36]
+ la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40]
+ la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45]
+ la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4]
+ la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54]
+ la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59]
+ la_oenb_mprj[5] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63]
+ la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68]
+ la_oenb_mprj[69] la_oenb_mprj[6] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72]
+ la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77]
+ la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[7] la_oenb_mprj[80] la_oenb_mprj[81]
+ la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86]
+ la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[8] la_oenb_mprj[90]
+ la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95]
+ la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[9]
+ mprj_ack_i_core mprj_ack_i_user mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11]
+ mprj_adr_o_core[12] mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15]
+ mprj_adr_o_core[16] mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19]
+ mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23]
+ mprj_adr_o_core[24] mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27]
+ mprj_adr_o_core[28] mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31]
+ mprj_adr_o_core[3] mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7]
+ mprj_adr_o_core[8] mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11]
+ mprj_adr_o_user[12] mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15]
+ mprj_adr_o_user[16] mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19]
+ mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23]
+ mprj_adr_o_user[24] mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27]
+ mprj_adr_o_user[28] mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31]
+ mprj_adr_o_user[3] mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7]
+ mprj_adr_o_user[8] mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0]
+ mprj_dat_i_core[10] mprj_dat_i_core[11] mprj_dat_i_core[12] mprj_dat_i_core[13]
+ mprj_dat_i_core[14] mprj_dat_i_core[15] mprj_dat_i_core[16] mprj_dat_i_core[17]
+ mprj_dat_i_core[18] mprj_dat_i_core[19] mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21]
+ mprj_dat_i_core[22] mprj_dat_i_core[23] mprj_dat_i_core[24] mprj_dat_i_core[25]
+ mprj_dat_i_core[26] mprj_dat_i_core[27] mprj_dat_i_core[28] mprj_dat_i_core[29]
+ mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31] mprj_dat_i_core[3] mprj_dat_i_core[4]
+ mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7] mprj_dat_i_core[8] mprj_dat_i_core[9]
+ mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11] mprj_dat_i_user[12] mprj_dat_i_user[13]
+ mprj_dat_i_user[14] mprj_dat_i_user[15] mprj_dat_i_user[16] mprj_dat_i_user[17]
+ mprj_dat_i_user[18] mprj_dat_i_user[19] mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21]
+ mprj_dat_i_user[22] mprj_dat_i_user[23] mprj_dat_i_user[24] mprj_dat_i_user[25]
+ mprj_dat_i_user[26] mprj_dat_i_user[27] mprj_dat_i_user[28] mprj_dat_i_user[29]
+ mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31] mprj_dat_i_user[3] mprj_dat_i_user[4]
+ mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7] mprj_dat_i_user[8] mprj_dat_i_user[9]
+ mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13]
+ mprj_dat_o_core[14] mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17]
+ mprj_dat_o_core[18] mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21]
+ mprj_dat_o_core[22] mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25]
+ mprj_dat_o_core[26] mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29]
+ mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4]
+ mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9]
+ mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13]
+ mprj_dat_o_user[14] mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17]
+ mprj_dat_o_user[18] mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21]
+ mprj_dat_o_user[22] mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25]
+ mprj_dat_o_user[26] mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29]
+ mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4]
+ mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9]
+ mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2] mprj_sel_o_core[3]
+ mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3] mprj_stb_o_core
+ mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood user1_vdd_powergood
+ user2_vcc_powergood user2_vdd_powergood user_clock user_clock2 user_irq[0] user_irq[1]
+ user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2] user_irq_ena[0] user_irq_ena[1]
+ user_irq_ena[2] user_reset vccd vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd vssd1 vssd2
XFILLER_45_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_973 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_133 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[34\]_A input59/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_516 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[72\] vccd vssd user_to_mprj_in_gates\[72\]/B mprj_logic_high_inst/HI[402]
+ input357/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_8_1644 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input127_A la_data_out_core[96] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_439 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[50\] la_buf\[50\]/TE _642_/A la_buf_enable\[50\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_26_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_501_ _501_/Y _501_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_37_1808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_432_ _432_/Y _432_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_2_1276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2233 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_363_ _363_/A _363_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_input496_A la_oenb_mprj[82] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input92_A la_data_out_core[64] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_497 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2288 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1565 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[36\] _500_/Y la_data_in_core[36] la_buf\[36\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[108\] vccd vssd user_to_mprj_in_gates\[108\]/B mprj_logic_high_inst/HI[438]
+ input269/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_10_851 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[8\] user_wb_dat_gates\[8\]/Y input580/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_10_895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[25\]_A input49/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1419 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_553 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_715 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_217 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2008 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_910 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[25\] user_to_mprj_in_gates\[25\]/Y user_to_mprj_in_gates\[25\]/B
+ input49/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_53_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1763 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1985 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[16\]_A input39/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[100\]_A input5/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1469 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1197 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_129 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[76\] _339_/Y la_oenb_core[76] mprj_logic_high_inst/HI[278]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[98\] la_buf\[98\]/TE _361_/A la_buf_enable\[98\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[24\] _456_/Y mprj_dat_o_user[24] mprj_dat_buf\[24\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input244_A la_data_out_mprj[86] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2039 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[104\]_TE mprj_logic_high_inst/HI[306] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input411_A la_oenb_mprj[120] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input509_A la_oenb_mprj[94] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1062 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2041 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
X_415_ _415_/A _415_/Y vssd vccd vssd vccd sky130_fd_sc_hd__inv_12
XFILLER_41_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_346_ _346_/Y _346_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_35_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2063 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output728_A output728/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output630_A output630/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1177 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[122\]_A input285/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2174 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1137 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1560 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[4\] la_buf\[4\]/TE _596_/A la_buf_enable\[4\]/B vssd vccd vssd vccd
+ sky130_fd_sc_hd__and2b_1
XFILLER_31_1771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1211 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1807 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[127\]_TE mprj_logic_high_inst/HI[329] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_501 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2050 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_707 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[113\]_A input275/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[35\] vccd vssd user_to_mprj_in_gates\[35\]/B mprj_logic_high_inst/HI[365]
+ input316/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_30_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[13\] la_buf\[13\]/TE _605_/A la_buf_enable\[13\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_7_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_86 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input194_A la_data_out_mprj[40] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input361_A la_iena_mprj[76] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[41\]_TE la_buf\[41\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2007 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input459_A la_oenb_mprj[49] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input55_A la_data_out_core[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input626_A user_irq_ena[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[26\]_TE mprj_logic_high_inst/HI[228] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[92\]_A_N _355_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_501 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[104\]_A input265/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_581 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[30\]_A_N _622_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1891 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1711 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output678_A output678/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_329_ _329_/A _329_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_30_798 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1755 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1619 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[45\]_A_N _637_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[92\] user_to_mprj_in_gates\[92\]/Y user_to_mprj_in_gates\[92\]/B
+ input123/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_48_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1575 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1035 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_898 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_356 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1991 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_253 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[64\]_TE la_buf\[64\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_297 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[49\]_TE mprj_logic_high_inst/HI[251] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput504 vccd vssd _600_/A la_oenb_mprj[8] vssd vccd sky130_fd_sc_hd__buf_2
Xinput515 la_oenb_mprj[9] _601_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput526 vccd vssd _418_/A mprj_adr_o_core[18] vssd vccd sky130_fd_sc_hd__buf_2
Xinput537 vccd vssd _428_/A mprj_adr_o_core[28] vssd vccd sky130_fd_sc_hd__buf_2
Xinput559 mprj_dat_i_user[18] input559/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
Xuser_to_mprj_oen_buffers\[109\] _372_/Y la_oenb_core[109] mprj_logic_high_inst/HI[311]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_29_821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput548 mprj_adr_o_core[9] _409_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_ena_buf\[93\]_A input380/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[39\] _631_/Y la_oenb_core[39] mprj_logic_high_inst/HI[241]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_16_515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input207_A la_data_out_mprj[52] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input576_A mprj_dat_i_user[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_246 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[13\]_TE mprj_dat_buf\[13\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_441 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1895 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__402__A _402_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2173 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[84\]_A input370/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_662 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[62\] user_to_mprj_in_gates\[62\]/Y output713/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_50_805 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1221 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[87\]_TE la_buf\[87\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[20\] user_wb_dat_gates\[20\]/Y input562/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_50_1421 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1427 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[75\]_A input360/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_161 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_120 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1029 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_304 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_540 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1983 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1169 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[80\] la_buf\[80\]/TE _343_/A la_buf_enable\[80\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xinput301 vssd vccd input301/X la_iena_mprj[21] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput312 vccd vssd la_iena_mprj[31] input312/X vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input157_A la_data_out_mprj[122] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_949 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput334 vssd vccd input334/X la_iena_mprj[51] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput323 vssd vccd input323/X la_iena_mprj[41] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput345 vssd vccd input345/X la_iena_mprj[61] vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_input324_A la_iena_mprj[42] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput356 vssd vccd input356/X la_iena_mprj[71] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput367 vssd vccd input367/X la_iena_mprj[81] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput378 vssd vccd input378/X la_iena_mprj[91] vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_in_ena_buf\[66\]_A input350/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input18_A la_data_out_core[112] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1645 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput389 _363_/A la_oenb_mprj[100] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[66\] _530_/Y la_data_in_core[66] la_buf\[66\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_45_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_594_ _594_/A _594_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_38_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1785 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1173 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[122\] _586_/Y la_data_in_core[122] la_buf\[122\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_8_599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[70\]_B user_to_mprj_in_gates\[70\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1681 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1578 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output710_A output710/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[57\]_A input340/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1876 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[55\] user_to_mprj_in_gates\[55\]/Y user_to_mprj_in_gates\[55\]/B
+ input82/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_48_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1694 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1814 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[61\]_B user_to_mprj_in_gates\[61\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1309 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1776 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[48\]_A input330/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_495 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2150 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_189 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input274_A la_iena_mprj[112] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[52\]_B user_to_mprj_in_gates\[52\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1791 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input441_A la_oenb_mprj[32] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input539_A mprj_adr_o_core[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput120 vccd vssd input120/X la_data_out_core[8] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_1_764 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput131 vccd vssd input131/X la_data_out_core[9] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_ena_buf\[39\]_A input320/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_797 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput142 _573_/A la_data_out_mprj[109] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput153 la_data_out_mprj[119] _583_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_48_245 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xinput164 la_data_out_mprj[13] _477_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput175 la_data_out_mprj[23] _487_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput186 la_data_out_mprj[33] _497_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_48_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_481 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput197 la_data_out_mprj[43] _507_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
X_646_ _646_/A _646_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_577_ _577_/A _577_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[6\]_A _438_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1869 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1257 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[25\] user_to_mprj_in_gates\[25\]/Y output672/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_16_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output660_A output660/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_886 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1593 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output758_A output758/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput627 vccd vssd la_data_in_mprj[0] output627/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_gates\[43\]_B user_to_mprj_in_gates\[43\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xoutput638 vccd vssd la_data_in_mprj[10] output638/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput649 vccd vssd la_data_in_mprj[11] output649/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_45_2065 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[112\]_TE la_buf\[112\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1397 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[27\]_TE mprj_adr_buf\[27\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_473 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_19 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2069 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[34\]_B user_to_mprj_in_gates\[34\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[95\]_A user_to_mprj_in_gates\[95\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[65\] vccd vssd user_to_mprj_in_gates\[65\]/B mprj_logic_high_inst/HI[395]
+ input349/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_6_2070 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__500__A _500_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_749 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_500_ _500_/Y _500_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_45_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[21\] _613_/Y la_oenb_core[21] mprj_logic_high_inst/HI[223]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[3\] _595_/Y la_oenb_core[3] mprj_logic_high_inst/HI[205]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[43\] la_buf\[43\]/TE _635_/A la_buf_enable\[43\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_26_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_431_ _431_/A _431_/Y vssd vccd vssd vccd sky130_fd_sc_hd__inv_8
XFILLER_26_97 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_362_ _362_/A _362_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_42_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input489_A la_oenb_mprj[76] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input391_A la_oenb_mprj[102] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input85_A la_data_out_core[58] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1820 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_863 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[122\]_A _586_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[29\] _493_/Y la_data_in_core[29] la_buf\[29\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_13_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[25\]_B user_to_mprj_in_gates\[25\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[86\]_A user_to_mprj_in_gates\[86\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1337 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_68 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__410__A _410_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_204 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1929 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_922 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_629_ _629_/A _629_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_in_buffers\[10\]_A user_to_mprj_in_gates\[10\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_32_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_410 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[18\] user_to_mprj_in_gates\[18\]/Y user_to_mprj_in_gates\[18\]/B
+ input41/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_buffers\[124\]_A user_to_mprj_in_gates\[124\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[113\]_A _577_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1953 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[16\]_B user_to_mprj_in_gates\[16\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[77\]_A user_to_mprj_in_gates\[77\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[28\] output776/A user_wb_dat_gates\[28\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_la_buf\[50\]_A _514_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[100\]_B user_to_mprj_in_gates\[100\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[82\]_TE mprj_logic_high_inst/HI[284] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1987 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2287 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[115\]_A user_to_mprj_in_gates\[115\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[104\]_A _568_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[68\]_A user_to_mprj_in_gates\[68\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[41\]_A _505_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_314 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[69\] _332_/Y la_oenb_core[69] mprj_logic_high_inst/HI[271]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_47_1993 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xmprj_dat_buf\[17\] _449_/Y mprj_dat_o_user[17] mprj_dat_buf\[17\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input237_A la_data_out_mprj[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1497 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input404_A la_oenb_mprj[114] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_218 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1074 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_414_ _414_/Y _414_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkinv_8
X_345_ _345_/Y _345_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_41_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_936 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[120\] vccd vssd user_to_mprj_in_gates\[120\]/B mprj_logic_high_inst/HI[450]
+ input283/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_buffers\[106\]_A user_to_mprj_in_gates\[106\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__405__A _405_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[59\]_A user_to_mprj_in_gates\[59\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_52_7 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[32\]_A _496_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[12\] _412_/Y mprj_adr_o_user[12] mprj_adr_buf\[12\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_48_1757 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[50\]_B la_buf_enable\[50\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[126\] user_to_mprj_in_gates\[126\]/Y output656/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
Xuser_to_mprj_in_buffers\[92\] user_to_mprj_in_gates\[92\]/Y output746/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_2_892 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1239 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1908 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_557 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[122\]_B mprj_logic_high_inst/HI[452] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[99\]_A _563_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[2\] output778/A user_wb_dat_gates\[2\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_33_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_785 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1572 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1783 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[23\]_A _487_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1223 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[41\]_B la_buf_enable\[41\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1109 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[113\]_B mprj_logic_high_inst/HI[443] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_719 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[28\] vccd vssd user_to_mprj_in_gates\[28\]/B mprj_logic_high_inst/HI[358]
+ input308/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_23_273 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_98 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input187_A la_data_out_mprj[34] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[14\]_A _478_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2019 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[32\]_B la_buf_enable\[32\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input354_A la_iena_mprj[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input48_A la_data_out_core[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[1\]_A input299/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input521_A mprj_adr_o_core[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input619_A mprj_stb_o_core vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[111\] la_buf\[111\]/TE _374_/A la_buf_enable\[111\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xla_buf\[96\] _560_/Y la_data_in_core[96] la_buf\[96\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[1\] vccd vssd user_to_mprj_in_gates\[1\]/B mprj_logic_high_inst/HI[331]
+ input299/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_8_1272 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[104\]_B mprj_logic_high_inst/HI[434] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_34_549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[99\]_B la_buf_enable\[99\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1171 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1767 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_991 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output740_A output740/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1003 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1587 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[23\]_B la_buf_enable\[23\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1047 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[85\] user_to_mprj_in_gates\[85\]/Y user_to_mprj_in_gates\[85\]/B
+ input115/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_6_1913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[92\]_A _355_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2328 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[14\]_B la_buf_enable\[14\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput516 mprj_ack_i_user input516/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
Xinput505 _353_/A la_oenb_mprj[90] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput527 _419_/A mprj_adr_o_core[19] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput549 vccd vssd mprj_cyc_o_core _393_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_2146 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput538 vccd vssd _429_/A mprj_adr_o_core[29] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_29_833 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[93\]_B mprj_logic_high_inst/HI[423] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_365 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1701 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input102_A la_data_out_core[73] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_869 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[83\]_A _346_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1907 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input471_A la_oenb_mprj[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input569_A mprj_dat_i_user[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[7\] _471_/Y la_data_in_core[7] la_buf\[7\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf\[11\] _475_/Y la_data_in_core[11] la_buf\[11\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_10_1675 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_497 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_118 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_107 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[4\] _404_/Y mprj_adr_o_user[4] mprj_adr_buf\[4\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_19_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[84\]_B mprj_logic_high_inst/HI[414] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1091 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1854 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_357 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[55\] user_to_mprj_in_gates\[55\]/Y output705/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_37_1233 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output690_A output690/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output788_A output788/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[117\]_TE mprj_logic_high_inst/HI[319] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1266 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[74\]_A _337_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1299 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[13\] user_wb_dat_gates\[13\]/Y input554/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_50_1477 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_781 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_wb_dat_buffers\[10\] output757/A user_wb_dat_gates\[10\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_48_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[1\]_A input561/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2350 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[111\] user_to_mprj_in_gates\[111\]/Y user_to_mprj_in_gates\[111\]/B
+ input17/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[75\]_B mprj_logic_high_inst/HI[405] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_633 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_132 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_677 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_165 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[31\]_TE la_buf\[31\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[1\]_A input43/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[65\]_A _657_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[16\]_TE mprj_logic_high_inst/HI[218] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[91\]_A_N _354_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_552 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__503__A _503_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[95\] vccd vssd user_to_mprj_in_gates\[95\]/B mprj_logic_high_inst/HI[425]
+ input382/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_27_2103 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_77 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[121\] _384_/Y la_oenb_core[121] mprj_logic_high_inst/HI[323]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_7_2208 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xmprj_sel_buf\[2\] _398_/Y mprj_sel_o_user[2] mprj_sel_buf\[2\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xinput302 vssd vccd input302/X la_iena_mprj[22] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput335 vssd vccd input335/X la_iena_mprj[52] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput324 vssd vccd input324/X la_iena_mprj[42] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput313 vssd vccd input313/X la_iena_mprj[32] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xuser_to_mprj_oen_buffers\[51\] _643_/Y la_oenb_core[51] mprj_logic_high_inst/HI[253]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[73\] la_buf\[73\]/TE _336_/A la_buf_enable\[73\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xinput346 vssd vccd input346/X la_iena_mprj[62] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput357 vssd vccd input357/X la_iena_mprj[72] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput368 vssd vccd input368/X la_iena_mprj[82] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput379 vssd vccd input379/X la_iena_mprj[92] vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_in_ena_buf\[66\]_B mprj_logic_high_inst/HI[396] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input317_A la_iena_mprj[36] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[44\]_A_N _636_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_593_ _593_/A _593_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_16_335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1520 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[59\] _523_/Y la_data_in_core[59] la_buf\[59\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_31_305 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[56\]_A _648_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[59\]_A_N _651_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1851 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[115\] _579_/Y la_data_in_core[115] la_buf\[115\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__413__A _413_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1546 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1513 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_405 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output703_A output703/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[57\]_B mprj_logic_high_inst/HI[387] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_48_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[54\]_TE la_buf\[54\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_2029 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[39\]_TE mprj_logic_high_inst/HI[241] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[48\] user_to_mprj_in_gates\[48\]/Y user_to_mprj_in_gates\[48\]/B
+ input74/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_1_1651 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_165 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[47\]_A _639_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1203 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1012 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1733 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2191 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[48\]_B mprj_logic_high_inst/HI[378] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1404 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2127 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_600 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[10\] vccd vssd user_to_mprj_in_gates\[10\]/B mprj_logic_high_inst/HI[340]
+ input271/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[38\]_A _630_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2162 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[99\] _362_/Y la_oenb_core[99] mprj_logic_high_inst/HI[301]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_31_87 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input267_A la_iena_mprj[106] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj2_vdd_pwrgood vccd vssd output791/A mprj2_vdd_pwrgood/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput110 vccd vssd input110/X la_data_out_core[80] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_46_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[77\]_TE la_buf\[77\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input434_A la_oenb_mprj[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input30_A la_data_out_core[123] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput121 vccd vssd input121/X la_data_out_core[90] vssd vccd sky130_fd_sc_hd__buf_4
Xinput132 la_data_out_mprj[0] _464_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput143 la_data_out_mprj[10] _474_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput154 la_data_out_mprj[11] _475_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_ena_buf\[39\]_B mprj_logic_high_inst/HI[369] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput165 vccd vssd la_data_out_mprj[14] _478_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput176 la_data_out_mprj[24] _488_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput187 la_data_out_mprj[34] _498_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_input601_A mprj_dat_o_core[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_622 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput198 vccd vssd la_data_out_mprj[44] _508_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_645_ _645_/Y _645_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_17_655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_576_ _576_/A _576_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__408__A _408_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[29\]_A _621_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[18\] user_to_mprj_in_gates\[18\]/Y output664/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_9_898 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output653_A output653/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput628 vccd vssd la_data_in_mprj[100] output628/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput639 vccd vssd la_data_in_mprj[110] output639/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_45_1321 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_581 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[25\]_A _425_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[26\]_TE mprj_dat_buf\[26\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_945 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1169 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[5\]_TE mprj_logic_high_inst/HI[207] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_50_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[2\]_A _594_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1099 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[16\]_A _416_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2082 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[58\] vccd vssd user_to_mprj_in_gates\[58\]/B mprj_logic_high_inst/HI[388]
+ input341/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_45_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_430_ _430_/Y _430_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkinv_8
XFILLER_26_65 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[14\] _606_/Y la_oenb_core[14] mprj_logic_high_inst/HI[216]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_361_ _361_/A _361_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
Xla_buf_enable\[36\] la_buf\[36\]/TE _628_/A la_buf_enable\[36\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_39_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input384_A la_iena_mprj[97] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_813 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input78_A la_data_out_core[51] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input551_A mprj_dat_i_user[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1009 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1145 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1251 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_216 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[0\]_TE mprj_sel_buf\[0\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1295 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_628_ _628_/A _628_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_33_934 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2335 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_559_ _559_/A _559_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output770_A output770/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1449 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__601__A _601_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1911 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1999 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2211 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_205 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_326 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__511__A _511_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_525 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input132_A la_data_out_mprj[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1487 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1031 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1593 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2010 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_413_ _413_/Y _413_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_6
XFILLER_53_41 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input599_A mprj_dat_o_core[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_344_ _344_/A _344_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_35_2054 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[41\] _505_/Y la_data_in_core[41] la_buf\[41\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[102\]_TE la_buf\[102\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[113\] vccd vssd user_to_mprj_in_gates\[113\]/B mprj_logic_high_inst/HI[443]
+ input275/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_mprj_adr_buf\[17\]_TE mprj_adr_buf\[17\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1695 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_153 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[1\]_TE mprj_adr_buf\[1\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__421__A _421_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[119\] user_to_mprj_in_gates\[119\]/Y output648/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_42_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[29\]_A _461_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[85\] user_to_mprj_in_gates\[85\]/Y output738/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_49_385 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[30\] user_to_mprj_in_gates\[30\]/Y user_to_mprj_in_gates\[30\]/B
+ input55/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_33_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_775 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[1\]_A _401_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__331__A _331_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[5\]_TE mprj_dat_buf\[5\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1763 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[27\]_A user_wb_dat_gates\[27\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_25_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2030 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1599 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[125\]_TE la_buf\[125\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_ack_gate_A input516/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2205 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__506__A _506_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1971 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[81\] _344_/Y la_oenb_core[81] mprj_logic_high_inst/HI[283]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_2_101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_3 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2345 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input347_A la_iena_mprj[63] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[1\]_B mprj_logic_high_inst/HI[331] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1666 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1104 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input514_A la_oenb_mprj[99] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[18\]_A user_wb_dat_gates\[18\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_46_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[89\] _553_/Y la_data_in_core[89] la_buf\[89\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[104\] la_buf\[104\]/TE _367_/A la_buf_enable\[104\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_46_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[72\]_TE mprj_logic_high_inst/HI[274] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_701 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1871 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__416__A _416_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output733_A output733/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1015 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[78\] user_to_mprj_in_gates\[78\]/Y user_to_mprj_in_gates\[78\]/B
+ input107/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_42_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1925 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_333 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[122\]_B la_buf_enable\[122\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2269 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[91\]_A input122/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj2_pwrgood_A mprj2_pwrgood/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput506 _354_/A la_oenb_mprj[91] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput517 mprj_adr_o_core[0] _400_/A vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
Xinput528 vccd vssd _401_/A mprj_adr_o_core[1] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_40_1806 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1413 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xinput539 mprj_adr_o_core[2] _402_/A vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
XFILLER_5_2158 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_333 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[113\]_B la_buf_enable\[113\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[40\] vccd vssd user_to_mprj_in_gates\[40\]/B mprj_logic_high_inst/HI[370]
+ input322/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[95\]_TE mprj_logic_high_inst/HI[297] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_561 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_65 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input297_A la_iena_mprj[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[4\]_A user_wb_dat_gates\[4\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[82\]_A input112/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input60_A la_data_out_core[35] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input464_A la_oenb_mprj[53] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[104\]_B la_buf_enable\[104\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[7\]_A _471_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_333 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[48\] user_to_mprj_in_gates\[48\]/Y output697/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_15_572 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2113 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output683_A output683/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1289 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[73\]_A input102/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[1\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1227 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1683 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2191 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[104\] user_to_mprj_in_gates\[104\]/Y user_to_mprj_in_gates\[104\]/B
+ input9/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_34_881 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[1\]_B user_to_mprj_in_gates\[1\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_40_328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[64\]_A input92/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2148 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[88\] vccd vssd user_to_mprj_in_gates\[88\]/B mprj_logic_high_inst/HI[418]
+ input374/X vssd vccd sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[114\] _377_/Y la_oenb_core[114] mprj_logic_high_inst/HI[316]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xinput303 vssd vccd input303/X la_iena_mprj[23] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput336 vssd vccd input336/X la_iena_mprj[53] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput325 vccd vssd la_iena_mprj[43] input325/X vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput314 vccd vssd la_iena_mprj[33] input314/X vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput347 vssd vccd input347/X la_iena_mprj[63] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput358 vssd vccd input358/X la_iena_mprj[73] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput369 vssd vccd input369/X la_iena_mprj[83] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xla_buf_enable\[66\] la_buf\[66\]/TE _329_/A la_buf_enable\[66\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[44\] _636_/Y la_oenb_core[44] mprj_logic_high_inst/HI[246]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_1_1107 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_irq_buffers\[2\] user_irq_gates\[2\]/Y output794/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
X_592_ _592_/Y _592_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_29_697 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input212_A la_data_out_mprj[57] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1532 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2119 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input581_A mprj_dat_i_user[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1142 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[55\]_A input82/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[108\] _572_/Y la_data_in_core[108] la_buf\[108\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_45_1558 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1569 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[101\] user_to_mprj_in_gates\[101\]/Y output629/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_48_973 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[5\]_A user_to_mprj_in_gates\[5\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_50_637 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1253 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__604__A _604_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[46\]_A input72/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1215 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1024 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[0\] _432_/Y mprj_dat_o_user[0] mprj_dat_buf\[0\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_6_2231 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1839 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1057 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_612 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1841 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2174 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__514__A _514_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[121\]_A input28/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[37\]_A input62/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_99 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1509 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input162_A la_data_out_mprj[127] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput111 vccd vssd input111/X la_data_out_core[81] vssd vccd sky130_fd_sc_hd__buf_4
Xinput100 vccd vssd input100/X la_data_out_core[71] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_42_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput122 vccd vssd input122/X la_data_out_core[91] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_44_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[107\]_TE mprj_logic_high_inst/HI[309] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input427_A la_oenb_mprj[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput133 _564_/A la_data_out_mprj[100] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput144 _574_/A la_data_out_mprj[110] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_input23_A la_data_out_core[117] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput166 vccd vssd la_data_out_mprj[15] _479_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput177 la_data_out_mprj[25] _489_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput155 vccd vssd _584_/A la_data_out_mprj[120] vssd vccd sky130_fd_sc_hd__buf_2
X_644_ _644_/A _644_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput199 vccd vssd la_data_out_mprj[45] _509_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput188 vccd vssd la_data_out_mprj[35] _499_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1477 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[71\] _535_/Y la_data_in_core[71] la_buf\[71\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_575_ _575_/Y _575_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_17_667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1827 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_800 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[28\]_A input52/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__424__A _424_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_383 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[112\]_A input18/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput629 vccd vssd la_data_in_mprj[101] output629/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_output646_A output646/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[21\]_TE la_buf\[21\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_247 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[90\]_A_N _353_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[60\] user_to_mprj_in_gates\[60\]/Y user_to_mprj_in_gates\[60\]/B
+ input88/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_48_781 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[19\]_A input42/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1061 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__334__A _334_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_A input8/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[43\]_A_N _635_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2265 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2107 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[58\]_A_N _650_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2094 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_217 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_902 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__509__A _509_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_360_ _360_/A _360_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_14_615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[29\] la_buf\[29\]/TE _621_/A la_buf_enable\[29\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_42_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1281 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1855 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_887 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[44\]_TE la_buf\[44\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input377_A la_iena_mprj[90] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2321 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[29\]_TE mprj_logic_high_inst/HI[231] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input544_A mprj_adr_o_core[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_707 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_228 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_627_ _627_/A _627_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA__419__A _419_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_946 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_475 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1791 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_558_ _558_/A _558_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_445 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_489_ _489_/Y _489_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_20_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[30\] user_to_mprj_in_gates\[30\]/Y output678/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_31_1900 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output763_A output763/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1392 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1381 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[1\]_B la_buf_enable\[1\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1923 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2223 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[125\]_A input288/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__329__A _329_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_721 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[67\]_TE la_buf\[67\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_305 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[70\] vccd vssd user_to_mprj_in_gates\[70\]/B mprj_logic_high_inst/HI[400]
+ input355/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_47_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[116\]_A input278/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input125_A la_data_out_core[94] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1561 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1054 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1087 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_412_ _412_/A _412_/Y vssd vccd vssd vccd sky130_fd_sc_hd__inv_12
XFILLER_53_75 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
X_343_ _343_/Y _343_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input494_A la_oenb_mprj[80] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input90_A la_data_out_core[62] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[34\] _498_/Y la_data_in_core[34] la_buf\[34\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_13_1630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[106\] vccd vssd user_to_mprj_in_gates\[106\]/B mprj_logic_high_inst/HI[436]
+ input267/X vssd vccd sky130_fd_sc_hd__and2_1
Xuser_wb_dat_gates\[6\] user_wb_dat_gates\[6\]/Y input578/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_13_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[16\]_TE mprj_dat_buf\[16\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_861 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2037 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1169 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[107\]_A input268/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[78\] user_to_mprj_in_gates\[78\]/Y output730/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_40_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_721 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_765 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[23\] user_to_mprj_in_gates\[23\]/Y user_to_mprj_in_gates\[23\]/B
+ input47/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_9_471 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__612__A _612_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1720 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2042 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1589 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1330 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_ack_gate_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_459 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1803 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__522__A _522_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1273 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1847 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[74\] _337_/Y la_oenb_core[74] mprj_logic_high_inst/HI[276]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[96\] la_buf\[96\]/TE _359_/A la_buf_enable\[96\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xoutput790 vccd vssd user2_vcc_powergood output790/A vssd vccd sky130_fd_sc_hd__buf_2
Xmprj_dat_buf\[22\] _454_/Y mprj_dat_o_user[22] mprj_dat_buf\[22\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input242_A la_data_out_mprj[84] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[96\]_A input383/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_301 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1932 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1296 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input507_A la_oenb_mprj[92] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_529 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1449 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_724 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[20\]_A input300/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__432__A _432_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_485 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output726_A output726/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1027 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[87\]_A input373/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_161 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__607__A _607_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1972 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1961 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[11\]_A input282/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[2\] la_buf\[2\]/TE _594_/A la_buf_enable\[2\]/B vssd vccd vssd vccd
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_gates\[91\]_B user_to_mprj_in_gates\[91\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA__342__A _342_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput507 _355_/A la_oenb_mprj[92] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput518 vccd vssd mprj_adr_o_core[10] _410_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_user_to_mprj_in_ena_buf\[78\]_A input363/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput529 mprj_adr_o_core[20] _420_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_29_857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_827 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[33\] vccd vssd user_to_mprj_in_gates\[33\]/B mprj_logic_high_inst/HI[363]
+ input314/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_3_1171 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__517__A _517_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_99 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[11\] la_buf\[11\]/TE _603_/A la_buf_enable\[11\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_32_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_739 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input192_A la_data_out_mprj[39] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[82\]_B user_to_mprj_in_gates\[82\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1810 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input457_A la_oenb_mprj[47] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input53_A la_data_out_core[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input624_A user_irq_ena[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1729 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[69\]_A input353/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1442 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_389 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1834 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1845 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__427__A _427_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_595 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output676_A output676/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[73\]_B user_to_mprj_in_gates\[73\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[115\]_TE la_buf\[115\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[90\] user_to_mprj_in_gates\[90\]/Y user_to_mprj_in_gates\[90\]/B
+ input121/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_48_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1239 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1701 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__337__A _337_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[64\]_B user_to_mprj_in_gates\[64\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[62\]_TE mprj_logic_high_inst/HI[264] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xinput326 vssd vccd input326/X la_iena_mprj[44] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput304 vssd vccd input304/X la_iena_mprj[24] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput315 vssd vccd input315/X la_iena_mprj[34] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xuser_to_mprj_oen_buffers\[107\] _370_/Y la_oenb_core[107] mprj_logic_high_inst/HI[309]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_40_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput337 vssd vccd input337/X la_iena_mprj[54] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput348 vssd vccd input348/X la_iena_mprj[64] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput359 vssd vccd input359/X la_iena_mprj[74] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_591_ _591_/Y _591_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[59\] la_buf\[59\]/TE _651_/A la_buf_enable\[59\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_16_315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[37\] _629_/Y la_oenb_core[37] mprj_logic_high_inst/HI[239]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input205_A la_data_out_mprj[50] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1290 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input574_A mprj_dat_i_user[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1739 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[55\]_B user_to_mprj_in_gates\[55\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1463 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1673 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1835 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2009 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[40\]_A user_to_mprj_in_gates\[40\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[60\] user_to_mprj_in_gates\[60\]/Y output711/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output793_A output793/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[9\]_A _441_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1065 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_863 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[46\]_B user_to_mprj_in_gates\[46\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[80\]_A _544_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[85\]_TE mprj_logic_high_inst/HI[287] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__620__A _620_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2243 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[31\]_A user_to_mprj_in_gates\[31\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_624 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1897 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_373 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[37\]_B user_to_mprj_in_gates\[37\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[98\]_A user_to_mprj_in_gates\[98\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[71\]_A _535_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[121\]_B user_to_mprj_in_gates\[121\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_5_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1813 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__530__A _530_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput101 vccd vssd input101/X la_data_out_core[72] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_46_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input155_A la_data_out_mprj[120] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput123 vccd vssd input123/X la_data_out_core[92] vssd vccd sky130_fd_sc_hd__buf_4
Xinput112 vccd vssd input112/X la_data_out_core[82] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_44_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput134 _565_/A la_data_out_mprj[101] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput145 vccd vssd _575_/A la_data_out_mprj[111] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_40_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input322_A la_iena_mprj[40] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput167 la_data_out_mprj[16] _480_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput178 vccd vssd la_data_out_mprj[26] _490_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput156 la_data_out_mprj[121] _585_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_input16_A la_data_out_core[110] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_643_ _643_/A _643_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_29_473 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[22\]_A user_to_mprj_in_gates\[22\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_17_613 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput189 vssd vccd _500_/A la_data_out_mprj[36] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_45_933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[30\]_A input573/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_574_ _574_/A _574_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
Xla_buf\[64\] _528_/Y la_data_in_core[64] la_buf\[64\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_17_679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1984 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1904 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1249 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[125\]_A _589_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_823 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[28\]_B user_to_mprj_in_gates\[28\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1650 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[89\]_A user_to_mprj_in_gates\[89\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[62\]_A _526_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[112\]_B user_to_mprj_in_gates\[112\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xla_buf\[120\] _584_/Y la_data_in_core[120] la_buf\[120\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xmprj_adr_buf\[28\] _428_/Y mprj_adr_o_user[28] mprj_adr_buf\[28\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[80\]_B la_buf_enable\[80\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__440__A _440_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output639_A output639/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1873 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[13\]_A user_to_mprj_in_gates\[13\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[53\] user_to_mprj_in_gates\[53\]/Y user_to_mprj_in_gates\[53\]/B
+ input80/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_3_1737 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[21\]_A input563/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_413 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[127\]_A user_to_mprj_in_gates\[127\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2028 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__615__A _615_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[116\]_A _580_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[19\]_B user_to_mprj_in_gates\[19\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[53\]_A _517_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_B user_to_mprj_in_gates\[103\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[71\]_B la_buf_enable\[71\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__350__A _350_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input8_A la_data_out_core[103] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1565 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_410 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[12\]_A input553/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_914 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_78 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[118\]_A user_to_mprj_in_gates\[118\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[107\]_A _571_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__525__A _525_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_77 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[44\]_A _508_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2008 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1867 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[62\]_B la_buf_enable\[62\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input272_A la_iena_mprj[110] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1591 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_16 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input537_A mprj_adr_o_core[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[127\] la_buf\[127\]/TE _390_/A la_buf_enable\[127\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_29_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_626_ _626_/A _626_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_487 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_557_ _557_/Y _557_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_buffers\[109\]_A user_to_mprj_in_gates\[109\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_488_ _488_/A _488_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA__435__A _435_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_620 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2050 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[35\]_A _499_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[23\] user_to_mprj_in_gates\[23\]/Y output670/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output756_A output756/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[53\]_B la_buf_enable\[53\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[120\]_A _383_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1131 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1979 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1039 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[125\]_B mprj_logic_high_inst/HI[455] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_3_2235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_218 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_774 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1812 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_777 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__345__A _345_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_608 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[26\]_A _490_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[44\]_B la_buf_enable\[44\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2041 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1985 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1805 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[111\]_A _374_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[63\] vccd vssd user_to_mprj_in_gates\[63\]/B mprj_logic_high_inst/HI[393]
+ input347/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_8_1467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1309 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[116\]_B mprj_logic_high_inst/HI[446] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input118_A la_data_out_core[88] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[41\] la_buf\[41\]/TE _633_/A la_buf_enable\[41\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[1\] _593_/Y la_oenb_core[1] mprj_logic_high_inst/HI[203]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_411_ _411_/Y _411_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_4
X_342_ _342_/Y _342_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf\[11\]_TE la_buf\[11\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input83_A la_data_out_core[56] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input487_A la_oenb_mprj[74] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[17\]_A _481_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[27\] _491_/Y la_data_in_core[27] la_buf\[27\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_13_1642 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_656 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[35\]_B la_buf_enable\[35\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[4\]_A input332/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[102\]_A _365_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_549 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1771 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[107\]_B mprj_logic_high_inst/HI[437] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1061 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_609_ _609_/A _609_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_la_buf_enable\[42\]_A_N _634_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1668 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_210 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[29\] user_wb_dat_gates\[29\]/Y input571/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_2
Xuser_to_mprj_in_gates\[16\] user_to_mprj_in_gates\[16\]/Y user_to_mprj_in_gates\[16\]/B
+ input39/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_53_1477 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[57\]_A_N _649_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[26\] output774/A user_wb_dat_gates\[26\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_la_buf_enable\[26\]_B la_buf_enable\[26\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1732 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[127\] user_to_mprj_in_gates\[127\]/Y user_to_mprj_in_gates\[127\]/B
+ input34/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_5_1629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2098 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[34\]_TE la_buf\[34\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1397 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[19\]_TE mprj_logic_high_inst/HI[221] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_221 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[95\]_A _358_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_57 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1951 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[17\]_B la_buf_enable\[17\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput780 vccd vssd mprj_dat_i_core[31] output780/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[67\] _330_/Y la_oenb_core[67] mprj_logic_high_inst/HI[269]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xoutput791 vccd vssd user2_vdd_powergood output791/A vssd vccd sky130_fd_sc_hd__buf_2
Xla_buf_enable\[89\] la_buf\[89\]/TE _352_/A la_buf_enable\[89\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_ena_buf\[96\]_B mprj_logic_high_inst/HI[426] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1231 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[15\] _447_/Y mprj_dat_o_user[15] mprj_dat_buf\[15\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_19_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input235_A la_data_out_mprj[78] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_357 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input402_A la_oenb_mprj[112] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2129 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[86\]_A _349_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_714 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[2\]_TE la_buf\[2\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[20\]_B mprj_logic_high_inst/HI[350] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_7_921 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2225 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[10\] _410_/Y mprj_adr_o_user[10] mprj_adr_buf\[10\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[124\] user_to_mprj_in_gates\[124\]/Y output654/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_oen_buffers\[10\]_A _602_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_692 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output719_A output719/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[87\]_B mprj_logic_high_inst/HI[417] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[57\]_TE la_buf\[57\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[90\] user_to_mprj_in_gates\[90\]/Y output744/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_42_1145 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_571 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_buffers\[0\] output756/A user_wb_dat_gates\[0\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_user_to_mprj_oen_buffers\[77\]_A _340_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1940 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[11\]_B mprj_logic_high_inst/HI[341] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA__623__A _623_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[4\]_A input576/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput508 vccd vssd _356_/A la_oenb_mprj[93] vssd vccd sky130_fd_sc_hd__buf_2
Xinput519 vssd vccd _411_/A mprj_adr_o_core[11] vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_in_ena_buf\[78\]_B mprj_logic_high_inst/HI[408] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1551 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_817 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_305 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[4\]_A input76/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_327 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[26\] vccd vssd user_to_mprj_in_gates\[26\]/B mprj_logic_high_inst/HI[356]
+ input306/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_52_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[68\]_A _331_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_574 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__533__A _533_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1369 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_77 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input185_A la_data_out_mprj[32] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1822 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1866 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input352_A la_iena_mprj[68] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input46_A la_data_out_core[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[69\]_B mprj_logic_high_inst/HI[399] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xla_buf\[94\] _558_/Y la_data_in_core[94] la_buf\[94\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input617_A mprj_sel_o_core[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_305 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[59\]_A _651_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1578 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output669_A output669/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__443__A _443_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1365 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[83\] user_to_mprj_in_gates\[83\]/Y user_to_mprj_in_gates\[83\]/B
+ input113/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_26_1630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1757 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[29\]_TE mprj_dat_buf\[29\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__618__A _618_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1492 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_809 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_850 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[8\]_TE mprj_logic_high_inst/HI[210] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_33_393 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__353__A _353_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1391 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1987 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_909 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xinput327 vssd vccd input327/X la_iena_mprj[45] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput305 vssd vccd input305/X la_iena_mprj[25] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput316 vssd vccd input316/X la_iena_mprj[35] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_29_600 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_78 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput338 vssd vccd input338/X la_iena_mprj[55] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput349 vssd vccd input349/X la_iena_mprj[65] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_590_ _590_/A _590_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_5_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__528__A _528_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_327 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input100_A la_data_out_core[71] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input567_A mprj_dat_i_user[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[5\] _469_/Y la_data_in_core[5] la_buf\[5\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_6_49 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_pwrgood_A mprj_pwrgood/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1505 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[3\]_TE mprj_sel_buf\[3\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[2\] _402_/Y mprj_adr_o_user[2] mprj_adr_buf\[2\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_441 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_165 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__438__A _438_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[53\] user_to_mprj_in_gates\[53\]/Y output703/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output786_A output786/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[10\]_A _442_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_875 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[11\] user_wb_dat_gates\[11\]/Y input552/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_34_1965 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[28\]_A _428_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2255 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1418 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__348__A _348_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[5\]_A _597_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2121 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[93\] vccd vssd user_to_mprj_in_gates\[93\]/B mprj_logic_high_inst/HI[423]
+ input380/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_mprj_adr_buf\[19\]_A _419_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput102 vccd vssd input102/X la_data_out_core[73] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_44_2261 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1869 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xmprj_sel_buf\[0\] _396_/Y mprj_sel_o_user[0] mprj_sel_buf\[0\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xinput124 vccd vssd input124/X la_data_out_core[93] vssd vccd sky130_fd_sc_hd__buf_4
Xinput113 vccd vssd input113/X la_data_out_core[83] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_40_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput135 la_data_out_mprj[102] _566_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_input148_A la_data_out_mprj[114] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2169 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[71\] la_buf\[71\]/TE _334_/A la_buf_enable\[71\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xinput168 la_data_out_mprj[17] _481_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput146 _576_/A la_data_out_mprj[112] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput157 _586_/A la_data_out_mprj[122] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
X_642_ _642_/A _642_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_29_441 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xinput179 vccd vssd la_data_out_mprj[27] _491_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_945 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input315_A la_iena_mprj[34] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[30\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_573_ _573_/A _573_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_44_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[57\] _521_/Y la_data_in_core[57] la_buf\[57\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[105\]_TE la_buf\[105\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_130 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1927 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_835 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1662 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_buffers\[2\]_A user_irq_gates\[2\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[113\] _577_/Y la_data_in_core[113] la_buf\[113\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_adr_buf\[4\]_TE mprj_adr_buf\[4\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1313 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output701_A output701/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[21\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[46\] user_to_mprj_in_gates\[46\]/Y input72/X user_to_mprj_in_gates\[46\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_23_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_469 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[52\]_TE mprj_logic_high_inst/HI[254] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2349 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1003 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__631__A _631_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[8\]_TE mprj_dat_buf\[8\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[8\] user_to_mprj_in_gates\[8\]/Y input120/X user_to_mprj_in_gates\[8\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_28_1533 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1340 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1373 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[12\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_639 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1851 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_89 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[97\] _360_/Y la_oenb_core[97] mprj_logic_high_inst/HI[299]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_13_1879 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__541__A _541_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input265_A la_iena_mprj[104] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_28 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input432_A la_oenb_mprj[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[90\]_TE la_buf\[90\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_411 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_625_ _625_/A _625_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_29_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[75\]_TE mprj_logic_high_inst/HI[277] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
X_556_ _556_/A _556_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_499 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_487_ _487_/Y _487_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_51_2073 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2062 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_632 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[16\] user_to_mprj_in_gates\[16\]/Y output662/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_47_2109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__451__A _451_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output749_A output749/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output651_A output651/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1706 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1728 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_786 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__626__A _626_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[4\]_A _404_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__361__A _361_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1478 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1953 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2097 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1341 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1479 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[56\] vccd vssd user_to_mprj_in_gates\[56\]/B mprj_logic_high_inst/HI[386]
+ input339/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_41_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[98\]_TE mprj_logic_high_inst/HI[300] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_410_ _410_/A _410_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_14_403 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_341_ _341_/Y _341_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA__536__A _536_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[12\] _604_/Y la_oenb_core[12] mprj_logic_high_inst/HI[214]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[34\] la_buf\[34\]/TE _626_/A la_buf_enable\[34\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_14_447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[8\] user_to_mprj_in_gates\[8\]/Y output743/A vccd vssd vssd
+ vccd sky130_fd_sc_hd__clkinv_4
XFILLER_35_1345 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_620 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input382_A la_iena_mprj[95] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1654 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input76_A la_data_out_core[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_668 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_830 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[4\]_B mprj_logic_high_inst/HI[334] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xmprj_stb_buf _394_/Y mprj_stb_o_user mprj_stb_buf/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_46_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_517 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_608_ _608_/A _608_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_2_2291 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__446__A _446_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_222 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output699_A output699/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_539_ _539_/A _539_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_417 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_wb_dat_buffers\[19\] output766/A user_wb_dat_gates\[19\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_5_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1744 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[125\]_B la_buf_enable\[125\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_517 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__356__A _356_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_553 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1665 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1643 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[94\]_A input125/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1253 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1963 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput781 vccd vssd mprj_dat_i_core[3] output781/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput770 vccd vssd mprj_dat_i_core[22] output770/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_43_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput792 vccd vssd user_irq[0] output792/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_8_1243 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[116\]_B la_buf_enable\[116\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input130_A la_data_out_core[99] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_77 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1118 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1287 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input228_A la_data_out_mprj[71] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_594 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_723 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_buffers\[7\]_A user_wb_dat_gates\[7\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input597_A mprj_dat_o_core[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[111\] vccd vssd user_to_mprj_in_gates\[111\]/B mprj_logic_high_inst/HI[441]
+ input273/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[85\]_A input115/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_clk_buf_A _391_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_977 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2259 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[30\]_TE mprj_adr_buf\[30\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[117\] user_to_mprj_in_gates\[117\]/Y output646/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf_enable\[107\]_B la_buf_enable\[107\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_837 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[83\] user_to_mprj_in_gates\[83\]/Y output736/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_18_583 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_542 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1952 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_A input105/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[4\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1923 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2045 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xinput509 vccd vssd _357_/A la_oenb_mprj[94] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_44_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[4\]_B user_to_mprj_in_gates\[4\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_24_520 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[19\] vccd vssd user_to_mprj_in_gates\[19\]/B mprj_logic_high_inst/HI[349]
+ input298/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_51_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[67\]_A input95/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1834 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input178_A la_data_out_mprj[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_936 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[41\]_A_N _633_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input345_A la_iena_mprj[61] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input39_A la_data_out_core[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[56\]_A_N _648_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input512_A la_oenb_mprj[97] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_133 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[87\] _551_/Y la_data_in_core[87] la_buf\[87\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_5_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[102\] la_buf\[102\]/TE _365_/A la_buf_enable\[102\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_46_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_545 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[58\]_A input85/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1860 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_785 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[24\]_TE la_buf\[24\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1929 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output731_A output731/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[76\] user_to_mprj_in_gates\[76\]/Y user_to_mprj_in_gates\[76\]/B
+ input105/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_38_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[8\]_A user_to_mprj_in_gates\[8\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1313 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_862 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__634__A _634_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[49\]_A input75/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1955 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1999 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xinput317 vssd vccd input317/X la_iena_mprj[36] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput306 vssd vccd input306/X la_iena_mprj[26] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_29_57 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xinput339 vssd vccd input339/X la_iena_mprj[56] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput328 vccd vssd la_iena_mprj[46] input328/X vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__544__A _544_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_865 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[124\]_A input31/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input295_A la_iena_mprj[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[47\]_TE la_buf\[47\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input462_A la_oenb_mprj[51] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_irq_ena_buf\[2\] vccd vssd user_irq_gates\[2\]/B user_irq_ena_buf\[2\]/B input626/X
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_4_799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1285 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1995 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_497 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1001 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[46\] user_to_mprj_in_gates\[46\]/Y output695/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_output681_A output681/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__454__A _454_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[115\]_A input21/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output779_A output779/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1049 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2195 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_943 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_965 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__629__A _629_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[102\] user_to_mprj_in_gates\[102\]/Y user_to_mprj_in_gates\[102\]/B
+ input7/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_53_445 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__364__A _364_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_A input11/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_386 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1763 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[86\] vccd vssd user_to_mprj_in_gates\[86\]/B mprj_logic_high_inst/HI[416]
+ input372/X vssd vccd sky130_fd_sc_hd__and2_1
Xinput125 input125/X la_data_out_core[94] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput114 vccd vssd input114/X la_data_out_core[84] vssd vccd sky130_fd_sc_hd__buf_4
Xinput103 vccd vssd input103/X la_data_out_core[74] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_49_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[112\] _375_/Y la_oenb_core[112] mprj_logic_high_inst/HI[314]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xinput136 la_data_out_mprj[103] _567_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_40_2137 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xinput169 la_data_out_mprj[18] _482_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput147 _577_/A la_data_out_mprj[113] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput158 vccd vssd _587_/A la_data_out_mprj[123] vssd vccd sky130_fd_sc_hd__buf_2
Xuser_to_mprj_oen_buffers\[42\] _634_/Y la_oenb_core[42] mprj_logic_high_inst/HI[244]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__539__A _539_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[64\] la_buf\[64\]/TE _656_/A la_buf_enable\[64\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
X_641_ _641_/Y _641_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_5_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_buffers\[0\] user_irq_gates\[0\]/Y output792/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_44_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2011 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input210_A la_data_out_mprj[55] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1942 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
X_572_ _572_/A _572_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_44_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input308_A la_iena_mprj[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_131 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_120 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2233 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1543 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[19\]_TE mprj_dat_buf\[19\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1674 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[106\] _570_/Y la_data_in_core[106] la_buf\[106\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__449__A _449_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2164 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_445 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[39\] user_to_mprj_in_gates\[39\]/Y user_to_mprj_in_gates\[39\]/B
+ input64/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_23_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_0 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1605 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_880 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[4\]_B la_buf_enable\[4\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__359__A _359_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_640 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input160_A la_data_out_mprj[125] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input258_A la_data_out_mprj[99] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1645 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1509 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[119\]_A input281/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input425_A la_oenb_mprj[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1149 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input21_A la_data_out_core[115] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_721 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[120\]_TE mprj_logic_high_inst/HI[322] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
X_624_ _624_/A _624_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_45_765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_467 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_555_ _555_/A _555_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
X_486_ _486_/Y _486_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_18_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_we_buf _395_/Y mprj_we_o_user mprj_we_buf/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[50\]_A input333/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_611 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2096 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_872 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output644_A output644/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xmprj_pwrgood vccd vssd output788/A mprj_pwrgood/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_29_1865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1019 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2290 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1525 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_798 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_245 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[41\]_A input323/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2261 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1869 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__642__A _642_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1397 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1447 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[49\] vccd vssd user_to_mprj_in_gates\[49\]/B mprj_logic_high_inst/HI[379]
+ input331/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_42_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_23 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_340_ _340_/Y _340_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_14_415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[32\]_A input313/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1493 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[27\] la_buf\[27\]/TE _619_/A la_buf_enable\[27\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA__552__A _552_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input375_A la_iena_mprj[89] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input69_A la_data_out_core[43] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1117 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[99\]_A input386/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input542_A mprj_adr_o_core[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[42\]_TE mprj_logic_high_inst/HI[244] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1751 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_607_ _607_/A _607_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_17_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_538_ _538_/Y _538_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_234 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[23\]_A input303/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1435 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_469_ _469_/A _469_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_289 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__462__A _462_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output761_A output761/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[118\]_TE la_buf\[118\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1756 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2181 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__637__A _637_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[14\]_A input293/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1699 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[94\]_B user_to_mprj_in_gates\[94\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA__372__A _372_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[80\]_TE la_buf\[80\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[65\]_TE mprj_logic_high_inst/HI[267] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput760 vccd vssd mprj_dat_i_core[13] output760/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput771 vccd vssd mprj_dat_i_core[23] output771/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput793 vccd vssd user_irq[1] output793/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_28_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1211 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput782 vccd vssd mprj_dat_i_core[4] output782/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_43_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2040 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_529 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input123_A la_data_out_core[92] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__547__A _547_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_540 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[1\]_A input625/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1831 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_we_buf_A _395_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input492_A la_oenb_mprj[79] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[85\]_B user_to_mprj_in_gates\[85\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xla_buf\[32\] _496_/Y la_data_in_core[32] la_buf\[32\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[104\] vccd vssd user_to_mprj_in_gates\[104\]/B mprj_logic_high_inst/HI[434]
+ input265/X vssd vccd sky130_fd_sc_hd__and2_1
Xuser_wb_dat_gates\[4\] user_wb_dat_gates\[4\]/Y input576/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_48_2205 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_484 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_477 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_989 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[70\]_A user_to_mprj_in_gates\[70\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_37_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[76\] user_to_mprj_in_gates\[76\]/Y output728/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_4_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__457__A _457_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_551 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_882 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_370 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_554 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[21\] user_to_mprj_in_gates\[21\]/Y user_to_mprj_in_gates\[21\]/B
+ input45/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_33_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_B user_to_mprj_in_gates\[76\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[88\]_TE mprj_logic_high_inst/HI[290] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1552 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[31\] output780/A user_wb_dat_gates\[31\]/Y vccd vssd vssd vccd
+ sky130_fd_sc_hd__inv_6
XFILLER_47_1025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[9\] _441_/Y mprj_dat_o_user[9] mprj_dat_buf\[9\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_5_2107 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1531 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[61\]_A user_to_mprj_in_gates\[61\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA__367__A _367_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2131 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_373 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[67\]_B user_to_mprj_in_gates\[67\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[72\] _335_/Y la_oenb_core[72] mprj_logic_high_inst/HI[274]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[94\] la_buf\[94\]/TE _357_/A la_buf_enable\[94\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_43_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[20\] _452_/Y mprj_dat_o_user[20] mprj_dat_buf\[20\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input338_A la_iena_mprj[55] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input240_A la_data_out_mprj[82] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[52\]_A user_to_mprj_in_gates\[52\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_19_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1732 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input505_A la_oenb_mprj[90] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_189 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_893 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_510 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_543 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_587 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[58\]_B user_to_mprj_in_gates\[58\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[92\]_A _556_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1872 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_753 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output724_A output724/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_992 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[43\]_A user_to_mprj_in_gates\[43\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[69\] user_to_mprj_in_gates\[69\]/Y user_to_mprj_in_gates\[69\]/B
+ input97/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_38_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_307 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_329 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_370 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[49\]_B user_to_mprj_in_gates\[49\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[83\]_A _547_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[0\] la_buf\[0\]/TE _592_/A la_buf_enable\[0\]/B vssd vccd vssd vccd
+ sky130_fd_sc_hd__and2b_1
XANTENNA__650__A _650_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput318 vssd vccd input318/X la_iena_mprj[37] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput307 vssd vccd input307/X la_iena_mprj[27] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[34\]_A user_to_mprj_in_gates\[34\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput329 vssd vccd input329/X la_iena_mprj[47] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1225 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[31\] vccd vssd user_to_mprj_in_gates\[31\]/B mprj_logic_high_inst/HI[361]
+ input312/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_45_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[20\]_TE mprj_adr_buf\[20\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_693 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_855 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[74\]_A _538_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[124\]_B user_to_mprj_in_gates\[124\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_8_539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input190_A la_data_out_mprj[37] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[92\]_B la_buf_enable\[92\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input288_A la_iena_mprj[125] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__560__A _560_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1621 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input455_A la_oenb_mprj[45] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1455 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input51_A la_data_out_core[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input622_A user_irq_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[25\]_A user_to_mprj_in_gates\[25\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1827 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1562 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[65\]_A _529_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[115\]_B user_to_mprj_in_gates\[115\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[39\] user_to_mprj_in_gates\[39\]/Y output687/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_30_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output674_A output674/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[83\]_B la_buf_enable\[83\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__470__A _470_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1705 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1197 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[16\]_A user_to_mprj_in_gates\[16\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1916 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[24\]_A input566/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1409 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[119\]_A _583_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[40\]_A_N _632_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__645__A _645_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[56\]_A _520_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_B user_to_mprj_in_gates\[106\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_31_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[74\]_B la_buf_enable\[74\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[55\]_A_N _647_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__380__A _380_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1731 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[79\] vccd vssd user_to_mprj_in_gates\[79\]/B mprj_logic_high_inst/HI[409]
+ input364/X vssd vccd sky130_fd_sc_hd__and2_1
Xinput126 input126/X la_data_out_core[95] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput115 vccd vssd input115/X la_data_out_core[85] vssd vccd sky130_fd_sc_hd__buf_4
Xinput104 vccd vssd input104/X la_data_out_core[75] vssd vccd sky130_fd_sc_hd__buf_4
Xuser_to_mprj_oen_buffers\[105\] _368_/Y la_oenb_core[105] mprj_logic_high_inst/HI[307]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xinput137 la_data_out_mprj[104] _568_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput148 vssd vccd _578_/A la_data_out_mprj[114] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput159 _588_/A la_data_out_mprj[124] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1180 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[15\]_A input556/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_640_ _640_/A _640_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_5_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_571_ _571_/A _571_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_44_413 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[57\] la_buf\[57\]/TE _649_/A la_buf_enable\[57\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[35\] _627_/Y la_oenb_core[35] mprj_logic_high_inst/HI[237]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_22_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1077 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2023 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1311 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[14\]_TE la_buf\[14\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input203_A la_data_out_mprj[49] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__555__A _555_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_132 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_121 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_110 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2289 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input99_A la_data_out_core[70] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[47\]_A _511_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input572_A mprj_dat_i_user[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[65\]_B la_buf_enable\[65\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1686 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_81 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1061 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_273 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output791_A output791/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1464 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_1 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__465__A _465_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_641 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[38\]_A _502_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[56\]_B la_buf_enable\[56\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[123\]_A _386_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[37\]_TE la_buf\[37\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_785 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_608 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__375__A _375_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_980 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[29\]_A _493_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_818 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[47\]_B la_buf_enable\[47\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[114\]_A _377_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1583 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_523 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1117 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input153_A la_data_out_mprj[119] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2093 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[119\]_B mprj_logic_high_inst/HI[449] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input320_A la_iena_mprj[39] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_623_ _623_/A _623_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_29_240 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input418_A la_oenb_mprj[127] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input14_A la_data_out_core[109] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[62\] _526_/Y la_data_in_core[62] la_buf\[62\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_45_777 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_554_ _554_/A _554_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
X_485_ _485_/Y _485_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_18_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[5\]_TE la_buf\[5\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[50\]_B mprj_logic_high_inst/HI[380] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[38\]_B la_buf_enable\[38\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[26\] _426_/Y mprj_adr_o_user[26] mprj_adr_buf\[26\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[7\]_A input365/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_884 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[40\]_A _632_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[105\]_A _368_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output637_A output637/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1281 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1167 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1719 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput490 _340_/A la_oenb_mprj[77] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xuser_to_mprj_in_gates\[51\] user_to_mprj_in_gates\[51\]/Y user_to_mprj_in_gates\[51\]/B
+ input78/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_35_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_427 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[41\]_B mprj_logic_high_inst/HI[371] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_31_471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1425 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[29\]_B la_buf_enable\[29\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_309 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[31\]_A _623_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input6_A la_data_out_core[101] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2233 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[98\]_A _361_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_427 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_769 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[32\]_B mprj_logic_high_inst/HI[362] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_637 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input368_A la_iena_mprj[82] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input270_A la_iena_mprj[109] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2144 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[22\]_A _614_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[99\]_B mprj_logic_high_inst/HI[429] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1421 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_876 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input535_A mprj_adr_o_core[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[125\] la_buf\[125\]/TE _388_/A la_buf_enable\[125\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_1_397 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1763 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1627 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[89\]_A _352_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_606_ _606_/A _606_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
X_537_ _537_/A _537_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_246 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[23\]_B mprj_logic_high_inst/HI[353] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
X_468_ _468_/Y _468_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_41_780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_399_ _399_/Y _399_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
Xuser_to_mprj_in_buffers\[21\] user_to_mprj_in_gates\[21\]/Y output668/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_9_475 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output754_A output754/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2320 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[13\]_A _605_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[99\] user_to_mprj_in_gates\[99\]/Y user_to_mprj_in_gates\[99\]/B
+ input130/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_29_1685 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2013 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1481 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_725 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[14\]_B mprj_logic_high_inst/HI[344] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_23_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__653__A _653_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_791 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[7\]_A input579/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[110\]_TE mprj_logic_high_inst/HI[312] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput750 vccd vssd la_data_in_mprj[96] output750/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput761 vccd vssd mprj_dat_i_core[14] output761/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput772 vccd vssd mprj_dat_i_core[24] output772/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1785 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput794 vccd vssd user_irq[2] output794/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_8_1223 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput783 vccd vssd mprj_dat_i_core[5] output783/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_43_1649 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1173 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[61\] vccd vssd user_to_mprj_in_gates\[61\]/B mprj_logic_high_inst/HI[391]
+ input345/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_41_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2052 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[7\]_A input109/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input116_A la_data_out_core[86] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_ena_buf\[1\]_B user_irq_ena_buf\[1\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1111 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__563__A _563_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input81_A la_data_out_core[54] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input485_A la_oenb_mprj[72] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_913 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[25\] _489_/Y la_data_in_core[25] la_buf\[25\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_6_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_496 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_809 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_861 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[69\] user_to_mprj_in_gates\[69\]/Y output720/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_382 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[27\] user_wb_dat_gates\[27\]/Y input569/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_33_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__473__A _473_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[14\] user_to_mprj_in_gates\[14\]/Y input37/X user_to_mprj_in_gates\[14\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_31_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1564 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_buffers\[24\] output772/A user_wb_dat_gates\[24\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_47_1037 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[125\] user_to_mprj_in_gates\[125\]/Y user_to_mprj_in_gates\[125\]/B
+ input32/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA__648__A _648_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_809 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[31\]_A _463_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_544 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_385 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__383__A _383_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_739 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[32\]_TE mprj_logic_high_inst/HI[234] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1615 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1085 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2125 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[65\] _657_/Y la_oenb_core[65] mprj_logic_high_inst/HI[267]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[87\] la_buf\[87\]/TE _350_/A la_buf_enable\[87\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_8_1031 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[13\] _445_/Y mprj_dat_o_user[13] mprj_dat_buf\[13\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_19_305 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input233_A la_data_out_mprj[76] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__558__A _558_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[108\]_TE la_buf\[108\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input400_A la_oenb_mprj[110] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[22\]_A _454_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_522 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_555 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_525 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_81 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[7\]_TE mprj_adr_buf\[7\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[122\] user_to_mprj_in_gates\[122\]/Y output652/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_3_971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output717_A output717/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__468__A _468_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[70\]_TE la_buf\[70\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[13\]_A _445_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_382 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_buffers\[20\]_A user_wb_dat_gates\[20\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[55\]_TE mprj_logic_high_inst/HI[257] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_385 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1085 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput308 vssd vccd input308/X la_iena_mprj[28] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput319 vssd vccd input319/X la_iena_mprj[38] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1351 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__378__A _378_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1395 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_105 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2205 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[8\]_A _600_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[11\]_A user_wb_dat_gates\[11\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_38_1537 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_503 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[24\] vccd vssd user_to_mprj_in_gates\[24\]/B mprj_logic_high_inst/HI[354]
+ input304/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_51_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2345 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input183_A la_data_out_mprj[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_256 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input448_A la_oenb_mprj[39] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input350_A la_iena_mprj[66] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input44_A la_data_out_core[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[92\] _556_/Y la_data_in_core[92] la_buf\[92\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[93\]_TE la_buf\[93\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input615_A mprj_sel_o_core[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_81 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1602 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[78\]_TE mprj_logic_high_inst/HI[280] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_vdd_pwrgood vccd vssd output789/A mprj_vdd_pwrgood/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_1574 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1957 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output667_A output667/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[81\] user_to_mprj_in_gates\[81\]/Y user_to_mprj_in_gates\[81\]/B
+ input111/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_6_1502 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1568 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[24\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_105 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_322 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_27 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1754 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1787 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput127 input127/X la_data_out_core[96] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput116 input116/X la_data_out_core[86] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput105 vccd vssd input105/X la_data_out_core[76] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_49_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput138 vssd vccd _569_/A la_data_out_mprj[105] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput149 _579_/A la_data_out_mprj[115] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1192 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[9\]_A_N _601_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1900 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[15\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_570_ _570_/Y _570_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_2_1933 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2035 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_469 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[28\] _620_/Y la_oenb_core[28] mprj_logic_high_inst/HI[230]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XPHY_100 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_650 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_133 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_122 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_111 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[0\]_A _464_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_193 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_697 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input398_A la_oenb_mprj[109] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__571__A _571_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input565_A mprj_dat_i_user[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[3\] _467_/Y la_data_in_core[3] la_buf\[3\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_49_2164 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1231 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_gates\[0\]_A input621/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_753 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[0\] _400_/Y mprj_adr_o_user[0] mprj_adr_buf\[0\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_7_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_2 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[51\] user_to_mprj_in_gates\[51\]/Y output701/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_44_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output784_A output784/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__481__A _481_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1618 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1039 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2237 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[10\]_TE mprj_adr_buf\[10\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__656__A _656_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[7\]_A _407_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_992 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1507 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__391__A _391_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_329 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[91\] vccd vssd user_to_mprj_in_gates\[91\]/B mprj_logic_high_inst/HI[421]
+ input378/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_46_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input146_A la_data_out_mprj[112] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_622_ _622_/A _622_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_29_252 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1989 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1967 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input313_A la_iena_mprj[32] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__566__A _566_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_553_ _553_/A _553_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_53_2319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[55\] _519_/Y la_data_in_core[55] la_buf\[55\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_484_ _484_/A _484_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_53_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[127\] vccd vssd user_to_mprj_in_gates\[127\]/B mprj_logic_high_inst/HI[457]
+ input290/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_18_1727 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1197 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_81 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_841 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[7\]_B mprj_logic_high_inst/HI[337] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[19\] _419_/Y mprj_adr_o_user[19] mprj_adr_buf\[19\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xla_buf\[111\] _575_/Y la_data_in_core[111] la_buf\[111\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_29_1845 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[99\] user_to_mprj_in_gates\[99\]/Y output753/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_7_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1641 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput480 la_oenb_mprj[68] _331_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput491 _341_/A la_oenb_mprj[78] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_la_buf_enable\[54\]_A_N _646_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__476__A _476_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[9\] output787/A user_wb_dat_gates\[9\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
Xuser_to_mprj_in_gates\[44\] user_to_mprj_in_gates\[44\]/Y user_to_mprj_in_gates\[44\]/B
+ input70/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_35_277 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[69\]_A_N _332_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2149 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[6\] user_to_mprj_in_gates\[6\]/Y input98/X user_to_mprj_in_gates\[6\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[30\]_A input55/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2289 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_550 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_561 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__386__A _386_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_2141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2049 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_439 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[97\]_A input128/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1337 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_601 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1640 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_634 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[95\] _358_/Y la_oenb_core[95] mprj_logic_high_inst/HI[297]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_48_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2123 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input263_A la_iena_mprj[102] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[21\]_A input45/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[119\]_B la_buf_enable\[119\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input430_A la_oenb_mprj[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input528_A mprj_adr_o_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[8\] vccd vssd user_to_mprj_in_gates\[8\]/B mprj_logic_high_inst/HI[338]
+ input376/X vssd vccd sky130_fd_sc_hd__and2_1
Xla_buf_enable\[118\] la_buf\[118\]/TE _381_/A la_buf_enable\[118\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_24_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_553 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1076 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_605_ _605_/Y _605_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_27_70 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_536_ _536_/Y _536_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_17_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[88\]_A input118/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_467_ _467_/Y _467_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_20_409 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1448 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
X_398_ _398_/Y _398_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_18_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1702 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[27\]_TE la_buf\[27\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[14\] user_to_mprj_in_gates\[14\]/Y output660/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_9_487 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output747_A output747/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[12\]_A input35/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1313 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2025 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[79\]_A input108/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[7\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_608 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput740 vccd vssd la_data_in_mprj[87] output740/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput751 vccd vssd la_data_in_mprj[97] output751/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput762 vccd vssd mprj_dat_i_core[15] output762/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput784 vccd vssd mprj_dat_i_core[6] output784/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput773 vccd vssd mprj_dat_i_core[25] output773/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_43_1617 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2064 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[7\]_B user_to_mprj_in_gates\[7\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[54\] vccd vssd user_to_mprj_in_gates\[54\]/B mprj_logic_high_inst/HI[384]
+ input337/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_41_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input109_A la_data_out_core[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_523 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[10\] _602_/Y la_oenb_core[10] mprj_logic_high_inst/HI[212]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_19_1822 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[32\] la_buf\[32\]/TE _624_/A la_buf_enable\[32\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_in_buffers\[6\] user_to_mprj_in_gates\[6\]/Y output721/A vccd vssd vssd
+ vccd sky130_fd_sc_hd__clkinv_4
XFILLER_14_269 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_413 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input380_A la_iena_mprj[93] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input478_A la_oenb_mprj[66] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input74_A la_data_out_core[48] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[18\] _482_/Y la_data_in_core[18] la_buf\[18\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_6_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1790 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_173 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_195 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1791 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_309 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output697_A output697/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1201 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_519_ _519_/Y _519_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_21_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1289 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[17\] user_wb_dat_gates\[17\]/Y output764/A vccd vssd vssd vccd
+ sky130_fd_sc_hd__clkinv_4
Xuser_to_mprj_in_gates\[118\] user_to_mprj_in_gates\[118\]/Y user_to_mprj_in_gates\[118\]/B
+ input24/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_3_1132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_501 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_556 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_707 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1329 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_917 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1561 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1425 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[58\] _650_/Y la_oenb_core[58] mprj_logic_high_inst/HI[260]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_8_1043 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_637 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_851 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input226_A la_data_out_mprj[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1817 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_865 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__574__A _574_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1229 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[127\]_A input34/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_397 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[100\]_A input261/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input595_A mprj_dat_o_core[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_559 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_751 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_983 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[115\] user_to_mprj_in_gates\[115\]/Y output644/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_46_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_637 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[81\] user_to_mprj_in_gates\[81\]/Y output734/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_37_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2017 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[100\]_TE mprj_logic_high_inst/HI[302] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__484__A _484_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_A input24/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1974 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1903 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput309 vssd vccd input309/X la_iena_mprj[29] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2181 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__394__A _394_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[109\]_A input14/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_161 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_813 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[17\] vccd vssd user_to_mprj_in_gates\[17\]/B mprj_logic_high_inst/HI[347]
+ input296/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_16_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_725 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input176_A la_data_out_mprj[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_268 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_769 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input343_A la_iena_mprj[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input37_A la_data_out_core[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__569__A _569_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[123\]_TE mprj_logic_high_inst/HI[325] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[85\] _549_/Y la_data_in_core[85] la_buf\[85\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_19_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input510_A la_oenb_mprj[95] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input608_A mprj_dat_o_core[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[100\] la_buf\[100\]/TE _363_/A la_buf_enable\[100\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_35_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_607 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1586 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[80\]_A input366/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_835 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_301 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_375 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__479__A _479_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[74\] user_to_mprj_in_gates\[74\]/Y user_to_mprj_in_gates\[74\]/B
+ input103/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_6_1514 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_401 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[22\]_TE mprj_logic_high_inst/HI[224] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_489 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_467 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_437 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[71\]_A input356/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_161 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1593 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[7\]_B la_buf_enable\[7\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1782 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput117 vccd vssd input117/X la_data_out_core[87] vssd vccd sky130_fd_sc_hd__buf_4
Xinput106 vccd vssd input106/X la_data_out_core[77] vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA__389__A _389_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput128 vccd vssd input128/X la_data_out_core[97] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_44_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput139 vccd vssd _570_/A la_data_out_mprj[106] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_44_1597 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1057 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1851 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2069 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[62\]_A input346/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_134 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_123 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_101 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_112 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_327 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input293_A la_iena_mprj[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input558_A mprj_dat_i_user[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input460_A la_oenb_mprj[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1243 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2176 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[60\]_TE la_buf\[60\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_ena_buf\[0\] vccd vssd user_irq_gates\[0\]/B user_irq_ena_buf\[0\]/B input624/X
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[45\]_TE mprj_logic_high_inst/HI[247] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1845 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_gates\[0\]_B user_irq_gates\[0\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_437 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1433 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[53\]_A input336/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_3 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_662 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_654 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[44\] user_to_mprj_in_gates\[44\]/Y output693/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_34_1733 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output777_A output777/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1007 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[1\]_A _397_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[100\] user_to_mprj_in_gates\[100\]/Y input5/X user_to_mprj_in_gates\[100\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_39_2345 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[44\]_A input326/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_816 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[83\]_TE la_buf\[83\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_1964 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_809 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1590 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[68\]_TE mprj_logic_high_inst/HI[270] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1563 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[84\] vccd vssd user_to_mprj_in_gates\[84\]/B mprj_logic_high_inst/HI[414]
+ input370/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_49_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[110\] _373_/Y la_oenb_core[110] mprj_logic_high_inst/HI[312]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[40\] _632_/Y la_oenb_core[40] mprj_logic_high_inst/HI[242]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[62\] la_buf\[62\]/TE _654_/A la_buf_enable\[62\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
X_621_ _621_/A _621_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_29_264 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input139_A la_data_out_mprj[106] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_245 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_552_ _552_/Y _552_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_ena_buf\[35\]_A input316/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input306_A la_iena_mprj[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1775 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_483_ _483_/A _483_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_13_643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[48\] _512_/Y la_data_in_core[48] la_buf\[48\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_34_1029 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__582__A _582_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[2\]_A _434_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[104\] _568_/Y la_data_in_core[104] la_buf\[104\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_7_2321 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput470 la_oenb_mprj[59] _651_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput481 la_oenb_mprj[69] _332_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_36_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput492 _342_/A la_oenb_mprj[79] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_36_757 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[26\]_A input306/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[37\] user_to_mprj_in_gates\[37\]/Y user_to_mprj_in_gates\[37\]/B
+ input62/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_1_1296 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_462 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__492__A _492_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[8\]_A_N _600_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2013 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1345 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[91\]_A user_to_mprj_in_gates\[91\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[30\]_B user_to_mprj_in_gates\[30\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1389 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1141 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1163 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1016 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[17\]_A input296/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1049 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_15 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_749 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_B user_to_mprj_in_gates\[97\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_22_451 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_646 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2113 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[88\] _351_/Y la_oenb_core[88] mprj_logic_high_inst/HI[290]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_11_1371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2157 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[21\]_B user_to_mprj_in_gates\[21\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input256_A la_data_out_mprj[97] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[82\]_A user_to_mprj_in_gates\[82\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__577__A _577_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input423_A la_oenb_mprj[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_604_ _604_/A _604_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
X_535_ _535_/A _535_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_27_82 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[88\]_B user_to_mprj_in_gates\[88\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_466_ _466_/Y _466_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_43_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_397_ _397_/A _397_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_40_292 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1714 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[31\] _431_/Y mprj_adr_o_user[31] mprj_adr_buf\[31\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_9_499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[120\]_A user_to_mprj_in_gates\[120\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2344 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output642_A output642/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_2208 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[73\]_A user_to_mprj_in_gates\[73\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[12\]_B user_to_mprj_in_gates\[12\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_97 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__487__A _487_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_521 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[79\]_B user_to_mprj_in_gates\[79\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_34_2083 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[111\]_A user_to_mprj_in_gates\[111\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[100\]_A _564_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput730 vccd vssd la_data_in_mprj[78] output730/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput741 vccd vssd la_data_in_mprj[88] output741/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput752 vccd vssd la_data_in_mprj[98] output752/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput763 vccd vssd mprj_dat_i_core[16] output763/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_48_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[64\]_A user_to_mprj_in_gates\[64\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xoutput785 vccd vssd mprj_dat_i_core[7] output785/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput774 vccd vssd mprj_dat_i_core[26] output774/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA__397__A _397_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1916 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[47\] vccd vssd user_to_mprj_in_gates\[47\]/B mprj_logic_high_inst/HI[377]
+ input329/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_mprj_adr_buf\[23\]_TE mprj_adr_buf\[23\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[25\] la_buf\[25\]/TE _617_/A la_buf_enable\[25\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_7_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[53\]_A_N _645_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_469 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input373_A la_iena_mprj[87] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[102\]_A user_to_mprj_in_gates\[102\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input67_A la_data_out_core[41] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input540_A mprj_adr_o_core[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[55\]_A user_to_mprj_in_gates\[55\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[68\]_A_N _331_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2241 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1645 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_896 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_518_ _518_/A _518_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[95\]_A _559_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_708 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_449_ _449_/Y _449_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_4
XFILLER_31_2289 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[46\]_A user_to_mprj_in_gates\[46\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1578 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1100 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1144 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_863 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2101 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_373 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[86\]_A _550_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_719 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[37\]_A user_to_mprj_in_gates\[37\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[10\]_A _474_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1055 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input121_A la_data_out_core[90] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[17\]_TE la_buf\[17\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_863 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input219_A la_data_out_mprj[63] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[77\]_A _541_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[127\]_B user_to_mprj_in_gates\[127\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1631 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[100\]_B mprj_logic_high_inst/HI[430] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input490_A la_oenb_mprj[77] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[95\]_B la_buf_enable\[95\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input588_A mprj_dat_o_core[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[30\] _494_/Y la_data_in_core[30] la_buf\[30\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__590__A _590_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[102\] vccd vssd user_to_mprj_in_gates\[102\]/B mprj_logic_high_inst/HI[432]
+ input263/X vssd vccd sky130_fd_sc_hd__and2_1
Xuser_wb_dat_gates\[2\] input572/X user_wb_ack_gate/B user_wb_dat_gates\[2\]/Y vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_8
XFILLER_6_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2303 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[28\]_A user_to_mprj_in_gates\[28\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[108\] user_to_mprj_in_gates\[108\]/Y output636/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_37_104 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2071 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[74\] user_to_mprj_in_gates\[74\]/Y output726/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_46_693 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[118\]_B user_to_mprj_in_gates\[118\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[68\]_A _532_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1043 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[86\]_B la_buf_enable\[86\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2097 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1959 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[19\]_A user_to_mprj_in_gates\[19\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[7\] _439_/Y mprj_dat_o_user[7] mprj_dat_buf\[7\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_wb_dat_gates\[27\]_A input569/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1757 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_39 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[10\]_B la_buf_enable\[10\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1470 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[109\]_B user_to_mprj_in_gates\[109\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[59\]_A _523_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[77\]_B la_buf_enable\[77\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1613 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1447 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input169_A la_data_out_mprj[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[70\] _333_/Y la_oenb_core[70] mprj_logic_high_inst/HI[272]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[92\] la_buf\[92\]/TE _355_/A la_buf_enable\[92\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_43_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[18\]_A input559/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input336_A la_iena_mprj[53] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_137 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2338 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[78\] _542_/Y la_data_in_core[78] la_buf\[78\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input503_A la_oenb_mprj[89] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__585__A _585_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1598 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[8\]_TE la_buf\[8\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[80\]_B mprj_logic_high_inst/HI[410] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_15_343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1038 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[68\]_B la_buf_enable\[68\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_571 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[70\]_A _333_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output722_A output722/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2205 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1526 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[67\] user_to_mprj_in_gates\[67\]/Y user_to_mprj_in_gates\[67\]/B
+ input95/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_4_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__495__A _495_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[71\]_B mprj_logic_high_inst/HI[401] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[59\]_B la_buf_enable\[59\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[61\]_A _653_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[126\]_A _389_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput118 vccd vssd input118/X la_data_out_core[88] vssd vccd sky130_fd_sc_hd__buf_4
Xinput107 vccd vssd input107/X la_data_out_core[78] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_44_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput129 input129/X la_data_out_core[98] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_44_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1957 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[62\]_B mprj_logic_high_inst/HI[392] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XPHY_124 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_113 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_102 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_135 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1369 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1623 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input286_A la_iena_mprj[123] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[117\]_A _380_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[52\]_A _644_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input453_A la_oenb_mprj[43] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1741 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input620_A mprj_we_o_core vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_917 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1985 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1581 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[53\]_B mprj_logic_high_inst/HI[383] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XPHY_4 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1701 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_666 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[37\] user_to_mprj_in_gates\[37\]/Y output685/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_30_165 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output672_A output672/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[43\]_A _635_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[108\]_A _371_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1480 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1841 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1885 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1378 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1080 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[44\]_B mprj_logic_high_inst/HI[374] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1656 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_460 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_165 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_828 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[113\]_TE mprj_logic_high_inst/HI[315] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[34\]_A _626_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_clk_buf_TE mprj_clk_buf/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[77\] vccd vssd user_to_mprj_in_gates\[77\]/B mprj_logic_high_inst/HI[407]
+ input362/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_44_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[103\] _366_/Y la_oenb_core[103] mprj_logic_high_inst/HI[305]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_620_ _620_/Y _620_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
X_551_ _551_/A _551_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[33\] _625_/Y la_oenb_core[33] mprj_logic_high_inst/HI[235]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_adr_buf\[30\]_A _430_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[55\] la_buf\[55\]/TE _647_/A la_buf_enable\[55\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_ena_buf\[35\]_B mprj_logic_high_inst/HI[365] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_482_ _482_/Y _482_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input201_A la_data_out_mprj[47] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2012 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input97_A la_data_out_core[69] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input570_A mprj_dat_i_user[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[12\]_TE mprj_logic_high_inst/HI[214] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[25\]_A _617_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput482 la_oenb_mprj[6] _598_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput471 vccd vssd _597_/A la_oenb_mprj[5] vssd vccd sky130_fd_sc_hd__buf_2
Xinput460 vccd vssd _596_/A la_oenb_mprj[4] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_7_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[21\]_A _421_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput493 vccd vssd _599_/A la_oenb_mprj[7] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_ena_buf\[26\]_B mprj_logic_high_inst/HI[356] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1264 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_441 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_997 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj2_vdd_pwrgood_A mprj2_vdd_pwrgood/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[16\]_A _608_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1851 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2069 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1313 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_725 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[12\]_A _412_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1991 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[17\]_B mprj_logic_high_inst/HI[347] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_41_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[50\]_TE la_buf\[50\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2321 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[35\]_TE mprj_logic_high_inst/HI[237] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_658 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[109\]_A_N _372_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[29\] _461_/Y mprj_dat_o_user[29] mprj_dat_buf\[29\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input151_A la_data_out_mprj[117] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1479 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_389 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input249_A la_data_out_mprj[90] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_603_ _603_/A _603_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_24_1799 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input416_A la_oenb_mprj[125] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input12_A la_data_out_core[107] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_61 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[60\] _524_/Y la_data_in_core[60] la_buf\[60\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_534_ _534_/Y _534_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_205 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_94 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2129 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__593__A _593_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_465_ _465_/Y _465_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_41_761 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_396_ _396_/Y _396_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_9_423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1726 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[24\] _424_/Y mprj_adr_o_user[24] mprj_adr_buf\[24\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_5_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output635_A output635/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2091 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2196 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[73\]_TE la_buf\[73\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1495 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xinput290 vssd vccd input290/X la_iena_mprj[127] vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_oen_buffers\[58\]_TE mprj_logic_high_inst/HI[260] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2305 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2349 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_271 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2095 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[9\] la_buf\[9\]/TE _601_/A la_buf_enable\[9\]/B vssd vccd vssd vccd
+ sky130_fd_sc_hd__and2b_1
Xoutput720 vccd vssd la_data_in_mprj[69] output720/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_43_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput731 vccd vssd la_data_in_mprj[79] output731/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput742 vccd vssd la_data_in_mprj[89] output742/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput753 vccd vssd la_data_in_mprj[99] output753/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_28_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput786 vccd vssd mprj_dat_i_core[8] output786/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput764 vccd vssd mprj_dat_i_core[17] output764/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput775 vccd vssd mprj_dat_i_core[27] output775/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input4_A la_data_out_core[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1321 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[22\]_TE mprj_dat_buf\[22\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[18\] la_buf\[18\]/TE _610_/A la_buf_enable\[18\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_oen_buffers\[1\]_TE mprj_logic_high_inst/HI[203] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_17_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input199_A la_data_out_mprj[45] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_949 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input366_A la_iena_mprj[80] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_irq_gates\[1\] user_irq_gates\[1\]/Y user_irq_gates\[1\]/B input622/X vssd vccd
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_11_1191 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input533_A mprj_adr_o_core[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__588__A _588_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[96\]_TE la_buf\[96\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[123\] la_buf\[123\]/TE _386_/A la_buf_enable\[123\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_4_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[25\]_A _457_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[7\]_A_N _599_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_517_ _517_/Y _517_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_2_1381 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_448_ _448_/Y _448_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
X_379_ _379_/Y _379_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_35_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output752_A output752/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[97\] user_to_mprj_in_gates\[97\]/Y user_to_mprj_in_gates\[97\]/B
+ input128/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA__498__A _498_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1112 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[16\]_A _448_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[23\]_A user_wb_dat_gates\[23\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_37_875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1156 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_569 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_ack_buffer_A user_wb_ack_gate/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1309 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1743 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1798 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2117 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_buffers\[14\]_A user_wb_dat_gates\[14\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_21_1769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input114_A la_data_out_core[84] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_385 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1687 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_580 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1810 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input483_A la_oenb_mprj[70] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[23\] _487_/Y la_data_in_core[23] la_buf\[23\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_7_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_245 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2326 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_473 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2083 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1421 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_99 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[67\] user_to_mprj_in_gates\[67\]/Y output718/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_45_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[25\] user_wb_dat_gates\[25\]/Y input567/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_2
Xuser_to_mprj_in_gates\[12\] user_to_mprj_in_gates\[12\]/Y input35/X user_to_mprj_in_gates\[12\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_31_2021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1927 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_wb_dat_buffers\[22\] output770/A user_wb_dat_gates\[22\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_mprj_adr_buf\[13\]_TE mprj_adr_buf\[13\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[27\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_617 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[123\] user_to_mprj_in_gates\[123\]/Y user_to_mprj_in_gates\[123\]/B
+ input30/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_la_buf_enable\[52\]_A_N _644_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_333 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_804 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_377 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[67\]_A_N _330_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2290 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1729 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[0\]_A user_wb_dat_gates\[0\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_749 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[85\] la_buf\[85\]/TE _348_/A la_buf_enable\[85\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[63\] _655_/Y la_oenb_core[63] mprj_logic_high_inst/HI[265]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_27_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[18\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[11\] _443_/Y mprj_dat_o_user[11] mprj_dat_buf\[11\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_0_977 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input231_A la_data_out_mprj[74] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[1\]_TE mprj_dat_buf\[1\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input329_A la_iena_mprj[47] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1785 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[3\]_A _467_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[100\]_B la_buf_enable\[100\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_355 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[121\]_TE la_buf\[121\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_314 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[127\] _591_/Y la_data_in_core[127] la_buf\[127\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_28_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[120\] user_to_mprj_in_gates\[120\]/Y output650/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_26_2167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output715_A output715/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2138 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1735 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[60\]_A input88/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput108 vccd vssd input108/X la_data_out_core[79] vssd vccd sky130_fd_sc_hd__buf_4
Xinput119 vccd vssd input119/X la_data_out_core[89] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_44_1533 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_125 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_114 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_103 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_664 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[22\] vccd vssd user_to_mprj_in_gates\[22\]/B mprj_logic_high_inst/HI[352]
+ input302/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_12_303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_483 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_136 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_697 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1061 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1083 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input181_A la_data_out_mprj[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input279_A la_iena_mprj[117] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[51\]_A input78/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1267 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input446_A la_oenb_mprj[37] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input42_A la_data_out_core[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput620 mprj_we_o_core _395_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA__596__A _596_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[90\] _554_/Y la_data_in_core[90] la_buf\[90\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_0_796 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input613_A mprj_dat_o_core[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_789 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[91\]_TE mprj_logic_high_inst/HI[293] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_5 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[1\]_A user_to_mprj_in_gates\[1\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1746 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_188 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_10 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1069 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output665_A output665/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_391 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[42\]_A input68/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1313 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2058 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_269 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_601 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1668 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1911 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_678 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_645 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_807 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1999 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput90 vccd vssd input90/X la_data_out_core[62] vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_user_to_mprj_in_gates\[33\]_A input58/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1227 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_550_ _550_/A _550_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_22_1683 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[48\] la_buf\[48\]/TE _640_/A la_buf_enable\[48\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
X_481_ _481_/Y _481_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
Xuser_to_mprj_oen_buffers\[8\] _600_/Y la_oenb_core[8] mprj_logic_high_inst/HI[210]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[26\] _618_/Y la_oenb_core[26] mprj_logic_high_inst/HI[228]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_25_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input396_A la_oenb_mprj[107] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input563_A mprj_dat_i_user[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[1\] _465_/Y la_data_in_core[1] la_buf\[1\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_5_833 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[24\]_A input48/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1031 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1116 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput461 la_oenb_mprj[50] _642_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput450 vccd vssd _632_/A la_oenb_mprj[40] vssd vccd sky130_fd_sc_hd__buf_4
Xinput472 vccd vssd _652_/A la_oenb_mprj[60] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_7_1677 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput483 vccd vssd _333_/A la_oenb_mprj[70] vssd vccd sky130_fd_sc_hd__buf_2
Xinput494 _343_/A la_oenb_mprj[80] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1794 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_954 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output782_A output782/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_671 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[15\]_A input38/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_217 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2177 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1752 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2090 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1362 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1395 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input144_A la_data_out_mprj[110] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1193 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_602_ _602_/Y _602_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input311_A la_iena_mprj[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input409_A la_oenb_mprj[119] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_533_ _533_/Y _533_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_33_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_464_ _464_/A _464_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
Xla_buf\[53\] _517_/Y la_data_in_core[53] la_buf\[53\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[125\] vccd vssd user_to_mprj_in_gates\[125\]/B mprj_logic_high_inst/HI[455]
+ input288/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_13_431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1841 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_395_ _395_/Y _395_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_9_435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_475 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1885 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[17\] _417_/Y mprj_adr_o_user[17] mprj_adr_buf\[17\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_4_77 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1981 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[97\] user_to_mprj_in_gates\[97\]/Y output751/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output628_A output628/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2153 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2017 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1485 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xinput280 vssd vccd input280/X la_iena_mprj[118] vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_oen_buffers\[103\]_TE mprj_logic_high_inst/HI[305] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xinput291 input291/X la_iena_mprj[12] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_3_1349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[42\] user_to_mprj_in_gates\[42\]/Y user_to_mprj_in_gates\[42\]/B
+ input68/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_buffers\[7\] output785/A user_wb_dat_gates\[7\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_36_2317 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[121\]_A input284/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1985 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_991 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput721 vccd vssd la_data_in_mprj[6] output721/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput710 vccd vssd la_data_in_mprj[5] output710/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput754 vccd vssd la_data_in_mprj[9] output754/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput743 vccd vssd la_data_in_mprj[8] output743/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput732 vccd vssd la_data_in_mprj[7] output732/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_28_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput787 vccd vssd mprj_dat_i_core[9] output787/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput765 vccd vssd mprj_dat_i_core[18] output765/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput776 vccd vssd mprj_dat_i_core[28] output776/A vssd vccd sky130_fd_sc_hd__buf_2
Xuser_to_mprj_in_gates\[4\] user_to_mprj_in_gates\[4\]/Y input76/X user_to_mprj_in_gates\[4\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_45_2181 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1177 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[112\]_A input274/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1803 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1284 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_581 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_467 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[93\] _356_/Y la_oenb_core[93] mprj_logic_high_inst/HI[295]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_2_622 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input261_A la_iena_mprj[100] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input359_A la_iena_mprj[74] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[126\]_TE mprj_logic_high_inst/HI[328] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input526_A mprj_adr_o_core[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[6\] vccd vssd user_to_mprj_in_gates\[6\]/B mprj_logic_high_inst/HI[336]
+ input354/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_49_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[116\] la_buf\[116\]/TE _379_/A la_buf_enable\[116\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_24_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1614 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_516_ _516_/A _516_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[103\]_A input264/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_447_ _447_/A _447_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_20_209 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
X_378_ _378_/Y _378_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_35_1660 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[12\] output658/A user_to_mprj_in_gates\[12\]/Y vssd vccd
+ vssd vccd sky130_fd_sc_hd__clkinv_8
XANTENNA_output745_A output745/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[40\]_TE la_buf\[40\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2321 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2198 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1464 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[25\]_TE mprj_logic_high_inst/HI[227] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1951 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_887 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2147 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[108\]_A_N _371_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1402 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1479 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1782 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_629 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[52\] vccd vssd user_to_mprj_in_gates\[52\]/B mprj_logic_high_inst/HI[382]
+ input335/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_8_1079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[92\]_A input379/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_301 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input107_A la_data_out_core[78] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_389 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[30\] la_buf\[30\]/TE _622_/A la_buf_enable\[30\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_24_41 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[4\] user_to_mprj_in_gates\[4\]/Y output699/A vccd vssd vssd
+ vccd sky130_fd_sc_hd__clkinv_4
XFILLER_51_890 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_592 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_725 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input476_A la_oenb_mprj[64] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input72_A la_data_out_core[46] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[16\] _480_/Y la_data_in_core[16] la_buf\[16\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[63\]_TE la_buf\[63\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1877 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[48\]_TE mprj_logic_high_inst/HI[250] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_95 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__599__A _599_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2338 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1085 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[9\] _409_/Y mprj_adr_o_user[9] mprj_adr_buf\[9\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2095 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[83\]_A input369/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_109 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_161 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1190 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output695_A output695/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_890 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_529 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1056 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[18\] user_wb_dat_gates\[18\]/Y input559/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_50_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[15\] user_wb_dat_gates\[15\]/Y output762/A vccd vssd vssd vccd
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_mprj_dat_buf\[12\]_TE mprj_dat_buf\[12\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1261 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[116\] user_to_mprj_in_gates\[116\]/Y user_to_mprj_in_gates\[116\]/B
+ input22/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[74\]_A input359/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1508 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[86\]_TE la_buf\[86\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1129 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[6\]_A_N _598_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[126\] _389_/Y la_oenb_core[126] mprj_logic_high_inst/HI[328]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_47_1361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[56\] _648_/Y la_oenb_core[56] mprj_logic_high_inst/HI[258]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[78\] la_buf\[78\]/TE _341_/A la_buf_enable\[78\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_48_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input224_A la_data_out_mprj[68] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[65\]_A input349/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_665 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_827 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input593_A mprj_dat_o_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_61 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2102 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[113\] user_to_mprj_in_gates\[113\]/Y output642/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_26_2179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_293 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_415 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output708_A output708/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[56\]_A input339/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1449 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_860 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1703 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[60\]_B user_to_mprj_in_gates\[60\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput109 vccd vssd input109/X la_data_out_core[7] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_5_1005 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1589 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[47\]_A input329/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1915 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_985 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_462 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_115 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_104 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_137 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_126 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[15\] vccd vssd user_to_mprj_in_gates\[15\]/B mprj_logic_high_inst/HI[345]
+ input294/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_16_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1505 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_197 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input174_A la_data_out_mprj[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[51\]_B user_to_mprj_in_gates\[51\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_4_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input341_A la_iena_mprj[58] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput621 vssd vccd input621/X user_irq_core[0] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1033 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input439_A la_oenb_mprj[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput610 _438_/A mprj_dat_o_core[6] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_input35_A la_data_out_core[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[83\] _547_/Y la_data_in_core[83] la_buf\[83\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input606_A mprj_dat_o_core[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[38\]_A input319/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_6 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_613 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[5\]_A _437_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_22 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output658_A output658/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[51\]_A_N _643_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[42\]_B user_to_mprj_in_gates\[42\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1990 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1791 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2037 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[72\] user_to_mprj_in_gates\[72\]/Y user_to_mprj_in_gates\[72\]/B
+ input101/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_41_1729 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[66\]_A_N _329_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_245 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[29\]_A input309/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1060 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1625 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_977 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_657 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1382 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1522 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput91 vccd vssd input91/X la_data_out_core[63] vssd vccd sky130_fd_sc_hd__buf_4
Xinput80 vccd vssd input80/X la_data_out_core[53] vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_la_buf_enable\[19\]_A_N _611_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[33\]_B user_to_mprj_in_gates\[33\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_1_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[94\]_A user_to_mprj_in_gates\[94\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[111\]_TE la_buf\[111\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1239 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[26\]_TE mprj_adr_buf\[26\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1745 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1756 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_480_ _480_/Y _480_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_0_2181 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2003 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[19\] _611_/Y la_oenb_core[19] mprj_logic_high_inst/HI[221]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_13_635 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_63 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input291_A la_iena_mprj[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input389_A la_oenb_mprj[100] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[121\]_A _585_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input556_A mprj_dat_i_user[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1043 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[85\]_A user_to_mprj_in_gates\[85\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[24\]_B user_to_mprj_in_gates\[24\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_4_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2263 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__400__A _400_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput462 vccd vssd _643_/A la_oenb_mprj[51] vssd vccd sky130_fd_sc_hd__buf_2
Xinput451 la_oenb_mprj[41] _633_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput440 vccd vssd _623_/A la_oenb_mprj[31] vssd vccd sky130_fd_sc_hd__buf_2
Xinput473 vccd vssd _653_/A la_oenb_mprj[61] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_3_1509 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput484 la_oenb_mprj[71] _334_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput495 vccd vssd _344_/A la_oenb_mprj[81] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_36_749 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2201 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[42\] user_to_mprj_in_gates\[42\]/Y output691/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_16_495 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1522 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output775_A output775/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[123\]_A user_to_mprj_in_gates\[123\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[112\]_A _576_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_193 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[15\]_B user_to_mprj_in_gates\[15\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[76\]_A user_to_mprj_in_gates\[76\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1673 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1155 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_226 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_421 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1043 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1764 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[114\]_A user_to_mprj_in_gates\[114\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[103\]_A _567_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[67\]_A user_to_mprj_in_gates\[67\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[40\]_A _504_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[82\] vccd vssd user_to_mprj_in_gates\[82\]/B mprj_logic_high_inst/HI[412]
+ input368/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[81\]_TE mprj_logic_high_inst/HI[283] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_329 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[60\] la_buf\[60\]/TE _652_/A la_buf_enable\[60\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
X_601_ _601_/A _601_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_18_727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input137_A la_data_out_mprj[104] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2232 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_532_ _532_/Y _532_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input304_A la_iena_mprj[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_463_ _463_/A _463_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_53_1419 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[46\] _510_/Y la_data_in_core[46] la_buf\[46\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_41_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_394_ _394_/A _394_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_51_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[118\] vccd vssd user_to_mprj_in_gates\[118\]/B mprj_logic_high_inst/HI[448]
+ input280/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_buffers\[105\]_A user_to_mprj_in_gates\[105\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_487 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[58\]_A user_to_mprj_in_gates\[58\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[31\]_A _495_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[102\] _566_/Y la_data_in_core[102] la_buf\[102\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_42_1813 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1453 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput270 vssd vccd input270/X la_iena_mprj[109] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput281 vssd vccd input281/X la_iena_mprj[119] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput292 vssd vccd input292/X la_iena_mprj[13] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_51_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_579 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[98\]_A _562_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[121\]_B mprj_logic_high_inst/HI[451] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[35\] user_to_mprj_in_gates\[35\]/Y user_to_mprj_in_gates\[35\]/B
+ input60/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_32_730 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1915 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_970 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput700 vccd vssd la_data_in_mprj[50] output700/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_buffers\[49\]_A user_to_mprj_in_gates\[49\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xoutput711 vccd vssd la_data_in_mprj[60] output711/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_la_buf\[22\]_A _486_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput722 vccd vssd la_data_in_mprj[70] output722/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput733 vccd vssd la_data_in_mprj[80] output733/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput744 vccd vssd la_data_in_mprj[90] output744/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput755 vccd vssd mprj_ack_i_core output755/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput766 vccd vssd mprj_dat_i_core[19] output766/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput777 vccd vssd mprj_dat_i_core[29] output777/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput788 vccd vssd user1_vcc_powergood output788/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_48_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[40\]_B la_buf_enable\[40\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1145 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_557 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[89\]_A _553_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[112\]_B mprj_logic_high_inst/HI[442] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2175 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[86\] _349_/Y la_oenb_core[86] mprj_logic_high_inst/HI[288]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[13\]_A _477_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1223 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1201 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_645 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_122 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input254_A la_data_out_mprj[95] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[31\]_B la_buf_enable\[31\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_678 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_188 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[0\]_A input260/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input421_A la_oenb_mprj[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input519_A mprj_adr_o_core[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[109\] vccd vssd la_buf\[109\]/TE la_buf_enable\[109\]/B _372_/A vssd
+ vccd sky130_fd_sc_hd__and2b_2
XFILLER_46_877 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_515_ _515_/Y _515_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_33_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[103\]_B mprj_logic_high_inst/HI[433] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1394 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_446_ _446_/A _446_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf_enable\[98\]_B la_buf_enable\[98\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_593 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_377_ _377_/A _377_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_35_1672 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2237 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1525 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output640_A output640/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2177 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output738_A output738/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[22\]_B la_buf_enable\[22\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1261 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1963 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1414 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[89\]_B la_buf_enable\[89\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[91\]_A _354_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1892 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2233 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[13\]_B la_buf_enable\[13\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1935 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_310 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[92\]_B mprj_logic_high_inst/HI[422] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[45\] vccd vssd user_to_mprj_in_gates\[45\]/B mprj_logic_high_inst/HI[375]
+ input327/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_43_836 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_357 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[23\] la_buf\[23\]/TE _615_/A la_buf_enable\[23\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_19_1667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_755 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[82\]_A _345_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input469_A la_oenb_mprj[58] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input371_A la_iena_mprj[85] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input65_A la_data_out_core[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1307 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_910 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_497 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1445 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[83\]_B mprj_logic_high_inst/HI[413] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_34_825 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_429_ _429_/A _429_/Y vssd vccd vssd vccd sky130_fd_sc_hd__inv_8
XANTENNA_output688_A output688/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2181 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[73\]_A _336_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1705 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[0\]_A input550/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1367 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput1 vssd vccd _391_/A caravel_clk vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_37_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[109\] user_to_mprj_in_gates\[109\]/Y user_to_mprj_in_gates\[109\]/B
+ input14/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[74\]_B mprj_logic_high_inst/HI[404] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_313 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[0\]_A input4/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[116\]_TE mprj_logic_high_inst/HI[318] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[64\]_A _656_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_217 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[119\] _382_/Y la_oenb_core[119] mprj_logic_high_inst/HI[321]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_47_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_917 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2319 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[49\] _641_/Y la_oenb_core[49] mprj_logic_high_inst/HI[251]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_19_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[65\]_B mprj_logic_high_inst/HI[395] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input217_A la_data_out_mprj[61] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[30\]_TE la_buf\[30\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[15\]_TE mprj_logic_high_inst/HI[217] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input586_A mprj_dat_o_core[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[55\]_A _647_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_501 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_73 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[100\] vccd vssd user_to_mprj_in_gates\[100\]/B mprj_logic_high_inst/HI[430]
+ input261/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_7_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[0\] user_wb_dat_gates\[0\]/Y input550/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_48_1115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__403__A _403_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[107\]_A_N _370_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[106\] user_to_mprj_in_gates\[106\]/Y output634/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_43_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_641 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[72\] user_to_mprj_in_gates\[72\]/Y output724/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_in_ena_buf\[56\]_B mprj_logic_high_inst/HI[386] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_47_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[30\] user_wb_dat_gates\[30\]/Y input573/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_33_2129 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_305 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[46\]_A _638_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[5\] _437_/Y mprj_dat_o_user[5] mprj_dat_buf\[5\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[47\]_B mprj_logic_high_inst/HI[377] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[53\]_TE la_buf\[53\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_953 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_116 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_105 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[38\]_TE mprj_logic_high_inst/HI[240] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XPHY_138 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_127 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_165 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_327 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[37\]_A _629_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input167_A la_data_out_mprj[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[90\] la_buf\[90\]/TE _353_/A la_buf_enable\[90\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xinput622 vssd vccd input622/X user_irq_core[1] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput611 vccd vssd _439_/A mprj_dat_o_core[7] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_7_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput600 mprj_dat_o_core[26] _458_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_27_1799 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input334_A la_iena_mprj[51] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input28_A la_data_out_core[121] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[38\]_B mprj_logic_high_inst/HI[368] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input501_A la_oenb_mprj[87] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[76\] _540_/Y la_data_in_core[76] la_buf\[76\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_441 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_7 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[28\]_A _620_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2209 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output720_A output720/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[76\]_TE la_buf\[76\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_725 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[24\]_A _424_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[29\]_B mprj_logic_high_inst/HI[359] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[65\] user_to_mprj_in_gates\[65\]/Y user_to_mprj_in_gates\[65\]/B
+ input93/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_6_1359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1072 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_249 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_953 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[5\]_A_N _597_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2062 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1815 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1935 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1394 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1225 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[19\]_A _611_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[1\]_A _593_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput81 vccd vssd input81/X la_data_out_core[54] vssd vccd sky130_fd_sc_hd__buf_4
Xinput70 input70/X la_data_out_core[44] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1534 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput92 vccd vssd input92/X la_data_out_core[64] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_44_1365 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_202 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1939 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[15\]_A _415_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[25\]_TE mprj_dat_buf\[25\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_901 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_934 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2026 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[4\]_TE mprj_logic_high_inst/HI[206] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_40_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_53 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input284_A la_iena_mprj[121] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input451_A la_oenb_mprj[41] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[99\]_TE la_buf\[99\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input549_A mprj_cyc_o_core vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput430 la_oenb_mprj[22] _614_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_48_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput463 la_oenb_mprj[52] _644_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput452 _634_/A la_oenb_mprj[42] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput441 vccd vssd _624_/A la_oenb_mprj[32] vssd vccd sky130_fd_sc_hd__buf_2
Xinput474 vccd vssd _654_/A la_oenb_mprj[62] vssd vccd sky130_fd_sc_hd__buf_2
Xinput485 vccd vssd _335_/A la_oenb_mprj[72] vssd vccd sky130_fd_sc_hd__buf_2
Xinput496 _345_/A la_oenb_mprj[82] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_35_205 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1289 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1534 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[35\] user_to_mprj_in_gates\[35\]/Y output683/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output670_A output670/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output768_A output768/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1870 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1589 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_588 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_238 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_761 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1743 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_466 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1033 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1618 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1055 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[75\] vccd vssd user_to_mprj_in_gates\[75\]/B mprj_logic_high_inst/HI[405]
+ input360/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA__501__A _501_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[101\] _364_/Y la_oenb_core[101] mprj_logic_high_inst/HI[303]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1955 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1015 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_600_ _600_/A _600_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
X_531_ _531_/A _531_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[31\] _623_/Y la_oenb_core[31] mprj_logic_high_inst/HI[233]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_18_739 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[53\] la_buf\[53\]/TE _645_/A la_buf_enable\[53\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_33_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1576 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_462_ _462_/Y _462_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_6
XANTENNA_la_buf_enable\[50\]_A_N _642_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_400 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_393_ _393_/Y _393_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_6
XANTENNA_input499_A la_oenb_mprj[85] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input95_A la_data_out_core[67] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[65\]_A_N _657_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[39\] _503_/Y la_data_in_core[39] la_buf\[39\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_51_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_665 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__411__A _411_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[28\]_A _460_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_893 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1869 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2261 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xinput260 vssd vccd input260/X la_iena_mprj[0] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput271 la_iena_mprj[10] input271/X vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_49_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput282 input282/X la_iena_mprj[11] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput293 vssd vccd input293/X la_iena_mprj[14] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_51_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[18\]_A_N _610_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_742 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[28\] user_to_mprj_in_gates\[28\]/Y user_to_mprj_in_gates\[28\]/B
+ input52/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_1_1097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2054 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1943 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[101\]_TE la_buf\[101\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[0\]_A _400_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[16\]_TE mprj_adr_buf\[16\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput701 vccd vssd la_data_in_mprj[51] output701/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput712 vccd vssd la_data_in_mprj[61] output712/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1684 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput723 vccd vssd la_data_in_mprj[71] output723/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput734 vccd vssd la_data_in_mprj[81] output734/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput745 vccd vssd la_data_in_mprj[91] output745/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput756 vccd vssd mprj_dat_i_core[0] output756/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput778 vccd vssd mprj_dat_i_core[2] output778/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput767 vccd vssd mprj_dat_i_core[1] output767/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_mprj_adr_buf\[0\]_TE mprj_adr_buf\[0\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput789 vccd vssd user1_vdd_powergood output789/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_mprj_dat_buf\[19\]_A _451_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[26\]_A user_wb_dat_gates\[26\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_45_1493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_385 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1841 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1420 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_602 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[79\] _342_/Y la_oenb_core[79] mprj_logic_high_inst/HI[281]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_49_105 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[27\] _459_/Y mprj_dat_o_user[27] mprj_dat_buf\[27\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_24_2223 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[4\]_TE mprj_dat_buf\[4\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input247_A la_data_out_mprj[89] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2317 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[0\]_B mprj_logic_high_inst/HI[330] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input414_A la_oenb_mprj[123] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[17\]_A user_wb_dat_gates\[17\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XANTENNA_input10_A la_data_out_core[105] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_514_ _514_/Y _514_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_2_1373 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[124\]_TE la_buf\[124\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1916 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_445_ _445_/A _445_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
X_376_ _376_/A _376_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA__406__A _406_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[22\] _422_/Y mprj_adr_o_user[22] mprj_adr_buf\[22\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_5_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output633_A output633/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[121\]_B la_buf_enable\[121\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_580 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_550 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[71\]_TE mprj_logic_high_inst/HI[273] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1735 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[7\] la_buf\[7\]/TE _599_/A la_buf_enable\[7\]/B vssd vccd vssd vccd
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_1779 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[90\]_A input121/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2289 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1820 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_609 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1831 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input2_A caravel_clk2 vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1947 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_322 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[112\]_B la_buf_enable\[112\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[38\] vccd vssd user_to_mprj_in_gates\[38\]/B mprj_logic_high_inst/HI[368]
+ input319/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_19_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_550 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1679 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_723 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[16\] la_buf\[16\]/TE _608_/A la_buf_enable\[16\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_11_767 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input197_A la_data_out_mprj[43] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_266 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[3\]_A user_wb_dat_gates\[3\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[81\]_A input111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input364_A la_iena_mprj[79] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_922 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input58_A la_data_out_core[33] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_432 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input531_A mprj_adr_o_core[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1953 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[121\] la_buf\[121\]/TE _384_/A la_buf_enable\[121\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_4_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[6\]_A _470_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_311 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[94\]_TE mprj_logic_high_inst/HI[296] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[103\]_B la_buf_enable\[103\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_428_ _428_/A _428_/Y vssd vccd vssd vccd sky130_fd_sc_hd__inv_8
XFILLER_31_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_359_ _359_/A _359_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_1367 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output750_A output750/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[72\]_A input101/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1790 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[95\] user_to_mprj_in_gates\[95\]/Y input126/X user_to_mprj_in_gates\[95\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_5_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1324 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[0\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput2 vssd vccd _392_/A caravel_clk2 vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[0\]_B user_to_mprj_in_gates\[0\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1278 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[63\]_A input91/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input112_A la_data_out_core[82] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_697 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1490 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input579_A mprj_dat_i_user[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input481_A la_oenb_mprj[69] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[21\] _485_/Y la_data_in_core[21] la_buf\[21\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_32_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1643 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_557 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[54\]_A input81/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1127 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_284 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_409 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_697 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[4\]_A user_to_mprj_in_gates\[4\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[65\] output716/A user_to_mprj_in_gates\[65\]/Y vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_37_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[23\] user_wb_dat_gates\[23\]/Y input565/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_2
Xuser_to_mprj_in_gates\[10\] user_to_mprj_in_gates\[10\]/Y input15/X user_to_mprj_in_gates\[10\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_14_391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1721 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_884 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[45\]_A input71/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[20\] output768/A user_wb_dat_gates\[20\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[121\] user_to_mprj_in_gates\[121\]/Y user_to_mprj_in_gates\[121\]/B
+ input28/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_53_910 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_921 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_106 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_139 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_998 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_117 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_128 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__504__A _504_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[120\]_A input27/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[36\]_A input61/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[61\] _653_/Y la_oenb_core[61] mprj_logic_high_inst/HI[263]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[83\] la_buf\[83\]/TE _346_/A la_buf_enable\[83\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xinput612 vccd vssd _440_/A mprj_dat_o_core[8] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_5_2220 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1817 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput601 vccd vssd _459_/A mprj_dat_o_core[27] vssd vccd sky130_fd_sc_hd__buf_2
Xinput623 vssd vccd input623/X user_irq_core[2] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_5_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input327_A la_iena_mprj[45] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1438 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[69\] _533_/Y la_data_in_core[69] la_buf\[69\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XPHY_8 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_497 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_844 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[27\]_A input51/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[111\]_A input17/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__414__A _414_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[125\] _589_/Y la_data_in_core[125] la_buf\[125\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_10_1771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output713_A output713/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1305 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[106\]_TE mprj_logic_high_inst/HI[308] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[58\] user_to_mprj_in_gates\[58\]/Y user_to_mprj_in_gates\[58\]/B
+ input85/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_39_1605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[18\]_A input41/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_A input7/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput82 vccd vssd input82/X la_data_out_core[55] vssd vccd sky130_fd_sc_hd__buf_4
Xinput71 vccd vssd input71/X la_data_out_core[45] vssd vccd sky130_fd_sc_hd__buf_4
Xinput60 vccd vssd input60/X la_data_out_core[35] vssd vccd sky130_fd_sc_hd__buf_4
Xinput93 vccd vssd input93/X la_data_out_core[65] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_48_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1480 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[20\]_TE la_buf\[20\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_214 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_751 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[20\] vccd vssd user_to_mprj_in_gates\[20\]/B mprj_logic_high_inst/HI[350]
+ input300/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_53_795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_946 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[106\]_A_N _369_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2038 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1337 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input277_A la_iena_mprj[115] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_357 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input40_A la_data_out_core[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input444_A la_oenb_mprj[35] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput420 la_oenb_mprj[13] _605_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_48_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput464 vccd vssd _645_/A la_oenb_mprj[53] vssd vccd sky130_fd_sc_hd__buf_2
Xinput453 vccd vssd _635_/A la_oenb_mprj[43] vssd vccd sky130_fd_sc_hd__buf_4
Xinput431 vccd vssd _615_/A la_oenb_mprj[23] vssd vccd sky130_fd_sc_hd__buf_2
Xinput442 vccd vssd _625_/A la_oenb_mprj[33] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input611_A mprj_dat_o_core[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput475 la_oenb_mprj[63] _655_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput486 _336_/A la_oenb_mprj[73] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput497 vccd vssd _346_/A la_oenb_mprj[83] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_5_1393 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__409__A _409_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[28\] user_to_mprj_in_gates\[28\]/Y output675/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output663_A output663/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1882 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[43\]_TE la_buf\[43\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[28\]_TE mprj_logic_high_inst/HI[230] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[0\]_B la_buf_enable\[0\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1168 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2125 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[124\]_A input287/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1711 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1343 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_817 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1873 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[68\] vccd vssd user_to_mprj_in_gates\[68\]/B mprj_logic_high_inst/HI[398]
+ input352/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_40_1005 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1715 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1185 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1027 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_10 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_707 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_530_ _530_/Y _530_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_ena_buf\[115\]_A input277/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2256 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[46\] la_buf\[46\]/TE _638_/A la_buf_enable\[46\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[24\] _616_/Y la_oenb_core[24] mprj_logic_high_inst/HI[226]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[6\] _598_/Y la_oenb_core[6] mprj_logic_high_inst/HI[208]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_461_ _461_/A _461_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_41_721 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_392_ _392_/A _392_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_13_412 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_467 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[66\]_TE la_buf\[66\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input394_A la_oenb_mprj[105] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input88_A la_data_out_core[60] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input561_A mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[4\]_A_N _596_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_393 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput250 la_data_out_mprj[91] _555_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput261 vssd vccd input261/X la_iena_mprj[100] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput272 vssd vccd input272/X la_iena_mprj[110] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput294 vssd vccd input294/X la_iena_mprj[15] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput283 vssd vccd input283/X la_iena_mprj[120] vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_in_ena_buf\[106\]_A input267/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_220 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output780_A output780/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput702 vccd vssd la_data_in_mprj[52] output702/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[15\]_TE mprj_dat_buf\[15\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__602__A _602_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput713 vccd vssd la_data_in_mprj[62] output713/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput724 vccd vssd la_data_in_mprj[72] output724/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput735 vccd vssd la_data_in_mprj[82] output735/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput746 vccd vssd la_data_in_mprj[92] output746/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput757 vccd vssd mprj_dat_i_core[10] output757/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput768 vccd vssd mprj_dat_i_core[20] output768/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput779 vccd vssd mprj_dat_i_core[30] output779/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_41_1314 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_548 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1897 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[89\]_TE la_buf\[89\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_721 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1839 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_437 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_459 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__512__A _512_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_636 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input142_A la_data_out_mprj[109] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[95\]_A input382/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2053 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input407_A la_oenb_mprj[117] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_513_ _513_/Y _513_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_37_1928 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_529 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_444_ _444_/Y _444_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_35_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[51\] _515_/Y la_data_in_core[51] la_buf\[51\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_375_ _375_/A _375_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_41_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[123\] vccd vssd user_to_mprj_in_gates\[123\]/B mprj_logic_high_inst/HI[453]
+ input286/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_13_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1505 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_441 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_997 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__422__A _422_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[15\] _415_/Y mprj_adr_o_user[15] mprj_adr_buf\[15\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_5_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[95\] user_to_mprj_in_gates\[95\]/Y output749/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_49_651 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1645 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[86\]_A input372/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_301 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1910 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_805 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[40\] user_to_mprj_in_gates\[40\]/Y user_to_mprj_in_gates\[40\]/B
+ input66/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_buffers\[5\] output783/A user_wb_dat_gates\[5\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_52_849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_562 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[10\]_A input271/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[90\]_B user_to_mprj_in_gates\[90\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA__332__A _332_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[2\] user_to_mprj_in_gates\[2\]/Y user_to_mprj_in_gates\[2\]/B
+ input54/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[77\]_A input362/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[64\]_A_N _656_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_161 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1603 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[79\]_A_N _342_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__507__A _507_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1836 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[81\]_B user_to_mprj_in_gates\[81\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_40_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[91\] _354_/Y la_oenb_core[91] mprj_logic_high_inst/HI[293]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[17\]_A_N _609_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_934 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input357_A la_iena_mprj[72] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1618 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_477 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[99\] _563_/Y la_data_in_core[99] la_buf\[99\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input524_A mprj_adr_o_core[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[4\] vccd vssd user_to_mprj_in_gates\[4\]/B mprj_logic_high_inst/HI[334]
+ input332/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_ena_buf\[68\]_A input352/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[114\] la_buf\[114\]/TE _377_/A la_buf_enable\[114\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_1_37 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_805 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_838 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1160 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_427_ _427_/Y _427_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkinv_8
XANTENNA__417__A _417_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_358_ _358_/A _358_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_2069 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[10\] output638/A user_to_mprj_in_gates\[10\]/Y vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_6
XANTENNA_user_to_mprj_in_gates\[72\]_B user_to_mprj_in_gates\[72\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1379 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output743_A output743/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[88\] user_to_mprj_in_gates\[88\]/Y user_to_mprj_in_gates\[88\]/B
+ input118/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[59\]_A input342/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_109 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput3 caravel_rstn input3/X vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1795 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2261 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1268 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_510 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1593 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[63\]_B user_to_mprj_in_gates\[63\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[114\]_TE la_buf\[114\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1397 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[29\]_TE mprj_adr_buf\[29\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_109 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[50\] vccd vssd user_to_mprj_in_gates\[50\]/B mprj_logic_high_inst/HI[380]
+ input333/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_27_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input105_A la_data_out_core[76] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[2\] user_to_mprj_in_gates\[2\]/Y output677/A vccd vssd vssd
+ vccd sky130_fd_sc_hd__clkinv_4
XFILLER_42_189 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_543 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input474_A la_oenb_mprj[62] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_587 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input70_A la_data_out_core[44] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[14\] _478_/Y la_data_in_core[14] la_buf\[14\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[54\]_B user_to_mprj_in_gates\[54\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1139 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[61\]_TE mprj_logic_high_inst/HI[263] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[7\] _407_/Y mprj_adr_o_user[7] mprj_adr_buf\[7\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_4_1244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_985 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[58\] user_to_mprj_in_gates\[58\]/Y output708/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_37_2289 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[8\]_A _440_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output693_A output693/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[16\] input557/X user_wb_ack_gate/B user_wb_dat_gates\[16\]/Y vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_8
XFILLER_31_1121 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_896 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1154 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[45\]_B user_to_mprj_in_gates\[45\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[13\] output760/A user_wb_dat_gates\[13\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_2205 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1111 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__610__A _610_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[114\] user_to_mprj_in_gates\[114\]/Y user_to_mprj_in_gates\[114\]/B
+ input20/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_38_974 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[30\]_A user_to_mprj_in_gates\[30\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_37_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_602 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_107 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_129 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_118 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1390 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1953 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[120\]_B user_to_mprj_in_gates\[120\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[36\]_B user_to_mprj_in_gates\[36\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[97\]_A user_to_mprj_in_gates\[97\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[70\]_A _534_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[98\] vccd vssd user_to_mprj_in_gates\[98\]/B mprj_logic_high_inst/HI[428]
+ input385/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_21_89 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[84\]_TE mprj_logic_high_inst/HI[286] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[124\] _387_/Y la_oenb_core[124] mprj_logic_high_inst/HI[326]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__520__A _520_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput613 _441_/A mprj_dat_o_core[9] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput602 mprj_dat_o_core[28] _460_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput624 vssd vccd input624/X user_irq_ena[0] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_48_705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[54\] _646_/Y la_oenb_core[54] mprj_logic_high_inst/HI[256]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_27_1768 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1069 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[76\] la_buf\[76\]/TE _339_/A la_buf_enable\[76\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_47_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[21\]_A user_to_mprj_in_gates\[21\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input222_A la_data_out_mprj[66] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1417 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_473 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_9 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_657 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input591_A mprj_dat_o_core[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2142 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1029 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[124\]_A _588_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1441 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_333 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[27\]_B user_to_mprj_in_gates\[27\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[111\]_B user_to_mprj_in_gates\[111\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[88\]_A user_to_mprj_in_gates\[88\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[61\]_A _525_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[118\] _582_/Y la_data_in_core[118] la_buf\[118\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_10_1783 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__430__A _430_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[111\] user_to_mprj_in_gates\[111\]/Y output640/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_39_705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output706_A output706/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[12\]_A user_to_mprj_in_gates\[12\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_35_933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_473 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1617 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[20\]_A input562/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2097 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[126\]_A user_to_mprj_in_gates\[126\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[115\]_A _579_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__605__A _605_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_693 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[18\]_B user_to_mprj_in_gates\[18\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[79\]_A user_to_mprj_in_gates\[79\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_B user_to_mprj_in_gates\[102\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput72 input72/X la_data_out_core[46] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput61 input61/X la_data_out_core[36] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput50 vccd vssd input50/X la_data_out_core[26] vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_la_buf\[52\]_A _516_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput94 input94/X la_data_out_core[66] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput83 input83/X la_data_out_core[56] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[70\]_B la_buf_enable\[70\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__340__A _340_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[11\]_A input552/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1127 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2017 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_413 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[13\] vccd vssd user_to_mprj_in_gates\[13\]/B mprj_logic_high_inst/HI[343]
+ input292/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_buffers\[117\]_A user_to_mprj_in_gates\[117\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__515__A _515_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[106\]_A _570_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[43\]_A _507_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1212 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input172_A la_data_out_mprj[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[61\]_B la_buf_enable\[61\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input437_A la_oenb_mprj[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput410 la_oenb_mprj[11] _603_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput421 vccd vssd _606_/A la_oenb_mprj[14] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_7_2349 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input33_A la_data_out_core[126] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput454 vccd vssd _636_/A la_oenb_mprj[44] vssd vccd sky130_fd_sc_hd__buf_2
Xinput432 _616_/A la_oenb_mprj[24] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput443 la_oenb_mprj[34] _626_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_48_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[81\] _545_/Y la_data_in_core[81] la_buf\[81\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xinput465 la_oenb_mprj[54] _646_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput476 vccd vssd _656_/A la_oenb_mprj[64] vssd vccd sky130_fd_sc_hd__buf_2
Xinput487 vccd vssd _337_/A la_oenb_mprj[74] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input604_A mprj_dat_o_core[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1203 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput498 vccd vssd _347_/A la_oenb_mprj[84] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_28_281 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_273 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[108\]_A user_to_mprj_in_gates\[108\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_457 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__425__A _425_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1894 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[34\]_A _498_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output656_A output656/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[52\]_B la_buf_enable\[52\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1621 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[70\] user_to_mprj_in_gates\[70\]/Y user_to_mprj_in_gates\[70\]/B
+ input99/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[124\]_B mprj_logic_high_inst/HI[454] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_35_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_270 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_402 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_clk_buf _391_/Y user_clock mprj_clk_buf/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_52_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__335__A _335_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[25\]_A _489_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1311 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[43\]_B la_buf_enable\[43\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1429 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1841 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[110\]_A _373_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_22 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[115\]_B mprj_logic_high_inst/HI[445] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
X_460_ _460_/A _460_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_2_1589 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_593 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[17\] _609_/Y la_oenb_core[17] mprj_logic_high_inst/HI[219]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_391_ _391_/Y _391_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[39\] la_buf\[39\]/TE _631_/A la_buf_enable\[39\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_40_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1113 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2270 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input387_A la_iena_mprj[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[16\]_A _480_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1591 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input554_A mprj_dat_i_user[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1605 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[34\]_B la_buf_enable\[34\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[3\]_A input321/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_833 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[101\]_A _364_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput240 vccd vssd _546_/A la_data_out_mprj[82] vssd vccd sky130_fd_sc_hd__buf_2
Xinput251 la_data_out_mprj[92] _556_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput262 vssd vccd input262/X la_iena_mprj[101] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_48_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput295 vssd vccd input295/X la_iena_mprj[16] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput273 vssd vccd input273/X la_iena_mprj[111] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput284 vssd vccd input284/X la_iena_mprj[121] vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_in_ena_buf\[106\]_B mprj_logic_high_inst/HI[436] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1044 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_589_ _589_/A _589_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[10\]_TE la_buf\[10\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[40\] user_to_mprj_in_gates\[40\]/Y output689/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_53_1956 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1907 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output773_A output773/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput703 vccd vssd la_data_in_mprj[53] output703/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_8_483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[25\]_B la_buf_enable\[25\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput714 vccd vssd la_data_in_mprj[63] output714/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput725 vccd vssd la_data_in_mprj[73] output725/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput736 vccd vssd la_data_in_mprj[83] output736/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1727 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput747 vccd vssd la_data_in_mprj[93] output747/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput758 vccd vssd mprj_dat_i_core[11] output758/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput769 vccd vssd mprj_dat_i_core[21] output769/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_la_buf_enable\[105\]_A_N _368_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_516 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[119\]_TE mprj_logic_high_inst/HI[321] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[94\]_A _357_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_939 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1477 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[16\]_B la_buf_enable\[16\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[80\] vccd vssd user_to_mprj_in_gates\[80\]/B mprj_logic_high_inst/HI[410]
+ input366/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_28_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[95\]_B mprj_logic_high_inst/HI[425] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_46_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_65 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input135_A la_data_out_mprj[102] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_869 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_512_ _512_/Y _512_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf\[33\]_TE la_buf\[33\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input302_A la_iena_mprj[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_443_ _443_/Y _443_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_14_711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[18\]_TE mprj_logic_high_inst/HI[220] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_585 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[85\]_A _348_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_374_ _374_/A _374_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_2207 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[44\] _508_/Y la_data_in_core[44] la_buf\[44\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_13_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[116\] vccd vssd user_to_mprj_in_gates\[116\]/B mprj_logic_high_inst/HI[446]
+ input278/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_10_983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1995 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_497 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[100\] _564_/Y la_data_in_core[100] la_buf\[100\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_9_1507 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[86\]_B mprj_logic_high_inst/HI[416] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_663 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[88\] user_to_mprj_in_gates\[88\]/Y output741/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_36_357 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[33\] user_to_mprj_in_gates\[33\]/Y user_to_mprj_in_gates\[33\]/B
+ input58/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_17_571 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[76\]_A _339_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_574 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1141 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[1\]_TE la_buf\[1\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1759 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[10\]_B mprj_logic_high_inst/HI[340] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA__613__A _613_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[3\]_A input575/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1281 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1905 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[77\]_B mprj_logic_high_inst/HI[407] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[56\]_TE la_buf\[56\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1877 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[3\]_A input65/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[3\]_A_N _595_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[67\]_A _330_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1659 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1848 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__523__A _523_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_77 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[84\] _347_/Y la_oenb_core[84] mprj_logic_high_inst/HI[286]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_2_401 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_456 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input252_A la_data_out_mprj[93] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[68\]_B mprj_logic_high_inst/HI[398] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input517_A mprj_adr_o_core[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[107\] la_buf\[107\]/TE _370_/A la_buf_enable\[107\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_4_1437 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1027 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[58\]_A _650_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_426_ _426_/A _426_/Y vssd vccd vssd vccd sky130_fd_sc_hd__inv_12
XFILLER_41_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_357_ _357_/A _357_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_35_1483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__433__A _433_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output736_A output736/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[79\]_TE la_buf\[79\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1315 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_990 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[59\]_B mprj_logic_high_inst/HI[389] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1359 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xinput4 vccd vssd input4/X la_data_out_core[0] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_52_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__608__A _608_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[49\]_A _641_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_522 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__343__A _343_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1321 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1229 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[28\]_TE mprj_dat_buf\[28\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[43\] vccd vssd user_to_mprj_in_gates\[43\]/B mprj_logic_high_inst/HI[373]
+ input325/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_27_165 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__518__A _518_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[7\]_TE mprj_logic_high_inst/HI[209] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[21\] la_buf\[21\]/TE _613_/A la_buf_enable\[21\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_23_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_555 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1071 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input63_A la_data_out_core[38] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input467_A la_oenb_mprj[56] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_264 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_253 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1256 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_ack_buffer output755/A user_wb_ack_gate/Y vssd vccd vssd vccd sky130_fd_sc_hd__clkinv_8
XFILLER_19_677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1501 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__428__A _428_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output686_A output686/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_409_ _409_/A _409_/Y vssd vccd vssd vccd sky130_fd_sc_hd__inv_8
XFILLER_14_371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1707 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[63\]_A_N _655_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1166 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_581 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[78\]_A_N _341_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[27\]_A _427_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1156 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[2\]_TE mprj_sel_buf\[2\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[107\] user_to_mprj_in_gates\[107\]/Y user_to_mprj_in_gates\[107\]/B
+ input12/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_52_433 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__338__A _338_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_119 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[16\]_A_N _608_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_108 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[4\]_A _596_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_385 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1206 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1449 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[18\]_A _418_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[117\] _380_/Y la_oenb_core[117] mprj_logic_high_inst/HI[319]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xinput603 mprj_dat_o_core[29] _461_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput625 vssd vccd input625/X user_irq_ena[1] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_48_717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput614 vccd vssd input614/X mprj_iena_wb vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[47\] _639_/Y la_oenb_core[47] mprj_logic_high_inst/HI[249]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[69\] la_buf\[69\]/TE _332_/A la_buf_enable\[69\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_47_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input215_A la_data_out_mprj[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input584_A mprj_dat_o_core[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_868 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_buffers\[1\]_A user_irq_gates\[1\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_389 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_717 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[104\] user_to_mprj_in_gates\[104\]/Y output632/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_43_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[70\] user_to_mprj_in_gates\[70\]/Y output722/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_53_219 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_945 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_433 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[20\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_477 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1807 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[104\]_TE la_buf\[104\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_628 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_680 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[19\]_TE mprj_adr_buf\[19\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput40 vccd vssd input40/X la_data_out_core[17] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_11_1504 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput73 vccd vssd input73/X la_data_out_core[47] vssd vccd sky130_fd_sc_hd__buf_4
Xinput62 input62/X la_data_out_core[37] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput51 input51/X la_data_out_core[27] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput95 input95/X la_data_out_core[67] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput84 input84/X la_data_out_core[57] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA__621__A _621_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[3\]_TE mprj_adr_buf\[3\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[3\] _435_/Y mprj_dat_o_user[3] mprj_dat_buf\[3\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_45_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[11\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_241 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1139 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_469 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[51\]_TE mprj_logic_high_inst/HI[253] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_304 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1003 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1224 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_849 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__531__A _531_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input165_A la_data_out_mprj[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[7\]_TE mprj_dat_buf\[7\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput400 _373_/A la_oenb_mprj[110] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput411 la_oenb_mprj[120] _383_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_48_525 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput455 la_oenb_mprj[45] _637_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_input332_A la_iena_mprj[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput422 la_oenb_mprj[15] _607_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput433 vccd vssd _617_/A la_oenb_mprj[25] vssd vccd sky130_fd_sc_hd__buf_2
Xinput444 la_oenb_mprj[35] _627_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_5_2041 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1649 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input26_A la_data_out_core[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput466 vccd vssd _647_/A la_oenb_mprj[55] vssd vccd sky130_fd_sc_hd__buf_2
Xinput477 la_oenb_mprj[65] _657_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput488 vccd vssd _338_/A la_oenb_mprj[75] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_5_2085 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1777 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_219 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput499 vccd vssd _348_/A la_oenb_mprj[85] vssd vccd sky130_fd_sc_hd__buf_4
Xla_buf\[74\] _538_/Y la_data_in_core[74] la_buf\[74\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[127\]_TE la_buf\[127\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_422 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1640 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_676 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__441__A _441_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output649_A output649/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2345 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[63\] user_to_mprj_in_gates\[63\]/Y user_to_mprj_in_gates\[63\]/B
+ input91/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_50_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[74\]_TE mprj_logic_high_inst/HI[276] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_753 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_414 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__616__A _616_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_609 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1003 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[3\]_A _403_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1979 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1334 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__351__A _351_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1903 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[29\]_A user_wb_dat_gates\[29\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_2_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_34 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2269 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_390_ _390_/A _390_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA__526__A _526_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_277 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_480 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1169 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_613 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input282_A la_iena_mprj[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_189 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input547_A mprj_adr_o_core[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[3\]_B mprj_logic_high_inst/HI[333] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2125 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_874 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput230 vccd vssd _537_/A la_data_out_mprj[73] vssd vccd sky130_fd_sc_hd__buf_2
Xinput241 _547_/A la_data_out_mprj[83] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput252 la_data_out_mprj[93] _557_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput263 vssd vccd input263/X la_iena_mprj[102] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_48_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[97\]_TE mprj_logic_high_inst/HI[299] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xinput296 vssd vccd input296/X la_iena_mprj[17] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput274 vssd vccd input274/X la_iena_mprj[112] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput285 vssd vccd input285/X la_iena_mprj[122] vssd vccd sky130_fd_sc_hd__clkbuf_1
X_657_ _657_/A _657_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
X_588_ _588_/Y _588_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__436__A _436_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[33\] user_to_mprj_in_gates\[33\]/Y output681/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output766_A output766/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_495 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput704 vccd vssd la_data_in_mprj[54] output704/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput715 vccd vssd la_data_in_mprj[64] output715/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput726 vccd vssd la_data_in_mprj[74] output726/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput737 vccd vssd la_data_in_mprj[84] output737/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput748 vccd vssd la_data_in_mprj[94] output748/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput759 vccd vssd mprj_dat_i_core[12] output759/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_28_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1305 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_333 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[124\]_B la_buf_enable\[124\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_528 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__346__A _346_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_907 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[93\]_A input124/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1205 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[73\] vccd vssd user_to_mprj_in_gates\[73\]/B mprj_logic_high_inst/HI[403]
+ input358/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_4_1608 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[115\]_B la_buf_enable\[115\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input128_A la_data_out_core[97] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1490 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2066 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_358 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_511_ _511_/Y _511_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[51\] la_buf\[51\]/TE _643_/A la_buf_enable\[51\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_2_1354 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
X_442_ _442_/A _442_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_14_723 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_553 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1621 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_373_ _373_/A _373_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_input497_A la_oenb_mprj[83] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input93_A la_data_out_core[65] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[6\]_A user_wb_dat_gates\[6\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[84\]_A input114/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[37\] _501_/Y la_data_in_core[37] la_buf\[37\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[109\] vccd vssd user_to_mprj_in_gates\[109\]/B mprj_logic_high_inst/HI[439]
+ input270/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_10_951 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[9\] user_wb_dat_gates\[9\]/Y input581/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_10_995 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_977 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1519 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1761 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[9\]_A _473_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[106\]_B la_buf_enable\[106\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[26\] user_to_mprj_in_gates\[26\]/Y user_to_mprj_in_gates\[26\]/B
+ input50/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_20_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[75\]_A input104/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1175 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[3\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1569 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1007 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1709 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_837 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1652 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[3\]_B user_to_mprj_in_gates\[3\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[66\]_A input94/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1242 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1985 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2230 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_218 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[77\] _340_/Y la_oenb_core[77] mprj_logic_high_inst/HI[279]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[99\] la_buf\[99\]/TE _362_/A la_buf_enable\[99\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_28_2181 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xmprj_dat_buf\[25\] _457_/Y mprj_dat_o_user[25] mprj_dat_buf\[25\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input245_A la_data_out_mprj[87] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_303 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input412_A la_oenb_mprj[121] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_358 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1716 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1705 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_425_ _425_/A _425_/Y vssd vccd vssd vccd sky130_fd_sc_hd__inv_12
XANTENNA_la_buf_enable\[104\]_A_N _367_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_356_ _356_/A _356_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[57\]_A input84/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[20\] _420_/Y mprj_adr_o_user[20] mprj_adr_buf\[20\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_48_1801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[119\]_A_N _382_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[109\]_TE mprj_logic_high_inst/HI[311] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1266 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output729_A output729/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output631_A output631/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2189 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1422 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xinput5 input5/X la_data_out_core[100] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_49_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_100 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[7\]_A user_to_mprj_in_gates\[7\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_637 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1551 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__624__A _624_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[48\]_A input74/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[5\] la_buf\[5\]/TE _597_/A la_buf_enable\[5\]/B vssd vccd vssd vccd
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[23\]_TE la_buf\[23\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1208 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1653 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1675 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[36\] vccd vssd user_to_mprj_in_gates\[36\]/B mprj_logic_high_inst/HI[366]
+ input317/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_42_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_309 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__534__A _534_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[14\] la_buf\[14\]/TE _606_/A la_buf_enable\[14\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_gates\[39\]_A input64/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[123\]_A input30/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1083 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input195_A la_data_out_mprj[41] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input362_A la_iena_mprj[77] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_210 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input56_A la_data_out_core[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_243 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_777 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_645 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_626 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_689 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_408_ _408_/Y _408_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkinv_16
XFILLER_14_383 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__444__A _444_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output679_A output679/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[114\]_A input20/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_339_ _339_/A _339_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_15_1855 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[46\]_TE la_buf\[46\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1134 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1877 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[93\] user_to_mprj_in_gates\[93\]/Y user_to_mprj_in_gates\[93\]/B
+ input124/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_48_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1041 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[2\]_A_N _594_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1168 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1285 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__619__A _619_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_497 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_626 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_109 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__354__A _354_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[105\]_A input10/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1218 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput604 vccd vssd _434_/A mprj_dat_o_core[2] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_5_2212 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xinput626 vssd vccd input626/X user_irq_ena[2] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput615 vccd vssd mprj_sel_o_core[0] _396_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_217 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_921 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__529__A _529_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2289 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_77 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input110_A la_data_out_core[80] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_968 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input208_A la_data_out_mprj[53] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1811 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[69\]_TE la_buf\[69\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_331 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input577_A mprj_dat_i_user[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1421 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_585 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_729 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__439__A _439_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[63\] user_to_mprj_in_gates\[63\]/Y output714/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_1_1942 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_692 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[21\] user_wb_dat_gates\[21\]/Y input563/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_50_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput30 input30/X la_data_out_core[123] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_15_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1565 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xinput63 input63/X la_data_out_core[38] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput52 input52/X la_data_out_core[28] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput41 vccd vssd input41/X la_data_out_core[18] vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_mprj_dat_buf\[18\]_TE mprj_dat_buf\[18\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput96 input96/X la_data_out_core[68] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput85 vccd vssd input85/X la_data_out_core[58] vssd vccd sky130_fd_sc_hd__buf_4
Xinput74 vccd vssd input74/X la_data_out_core[48] vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_la_buf_enable\[3\]_B la_buf_enable\[3\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2037 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[127\]_A input290/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__349__A _349_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1717 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_286 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_651 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_684 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1785 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[81\] la_buf\[81\]/TE _344_/A la_buf_enable\[81\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xinput401 vccd vssd _374_/A la_oenb_mprj[111] vssd vccd sky130_fd_sc_hd__buf_4
Xinput412 _384_/A la_oenb_mprj[121] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_input158_A la_data_out_mprj[123] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[118\]_A input280/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput445 la_oenb_mprj[36] _628_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput423 la_oenb_mprj[16] _608_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput434 la_oenb_mprj[26] _618_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput467 la_oenb_mprj[56] _648_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput456 vccd vssd _638_/A la_oenb_mprj[46] vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_input325_A la_iena_mprj[43] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput478 vccd vssd _329_/A la_oenb_mprj[66] vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_input19_A la_data_out_core[113] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[62\]_A_N _654_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput489 _339_/A la_oenb_mprj[76] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xla_buf\[67\] _531_/Y la_data_in_core[67] la_buf\[67\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_16_434 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[77\]_A_N _340_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_611 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_688 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_165 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[123\] _587_/Y la_data_in_core[123] la_buf\[123\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[15\]_A_N _607_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[109\]_A input270/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output711_A output711/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[56\] user_to_mprj_in_gates\[56\]/Y user_to_mprj_in_gates\[56\]/B
+ input83/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_35_721 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_253 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_297 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[40\]_A input322/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2030 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1173 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__632__A _632_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1959 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2248 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_46 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[31\]_A input312/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_245 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__542__A _542_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_492 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input275_A la_iena_mprj[113] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[98\]_A input385/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_853 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input442_A la_oenb_mprj[33] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_301 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xinput220 la_data_out_mprj[64] _528_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1425 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput231 vccd vssd _538_/A la_data_out_mprj[74] vssd vccd sky130_fd_sc_hd__buf_2
Xinput242 vccd vssd _548_/A la_data_out_mprj[84] vssd vccd sky130_fd_sc_hd__buf_4
Xinput253 vccd vssd _558_/A la_data_out_mprj[94] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_7_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput297 vssd vccd input297/X la_iena_mprj[18] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput264 vssd vccd input264/X la_iena_mprj[103] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput275 vssd vccd input275/X la_iena_mprj[113] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput286 vssd vccd input286/X la_iena_mprj[123] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_48_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2298 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_656_ _656_/A _656_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
X_587_ _587_/Y _587_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_16_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[22\]_A input302/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[26\] user_to_mprj_in_gates\[26\]/Y output673/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output661_A output661/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__452__A _452_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output759_A output759/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput705 vccd vssd la_data_in_mprj[55] output705/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput716 vccd vssd la_data_in_mprj[65] output716/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput727 vccd vssd la_data_in_mprj[75] output727/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_28_1117 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput738 vccd vssd la_data_in_mprj[85] output738/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput749 vccd vssd la_data_in_mprj[95] output749/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_ena_buf\[89\]_A input375/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2029 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2007 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[41\]_TE mprj_logic_high_inst/HI[243] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__627__A _627_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[13\]_A input292/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_289 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[93\]_B user_to_mprj_in_gates\[93\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__362__A _362_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[117\]_TE la_buf\[117\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1143 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[66\] vccd vssd user_to_mprj_in_gates\[66\]/B mprj_logic_high_inst/HI[396]
+ input350/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_6_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_510_ _510_/Y _510_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_2_1322 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[0\]_A input624/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[4\] _596_/Y la_oenb_core[4] mprj_logic_high_inst/HI[206]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__537__A _537_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[22\] _614_/Y la_oenb_core[22] mprj_logic_high_inst/HI[224]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_441_ _441_/A _441_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
Xla_buf_enable\[44\] la_buf\[44\]/TE _636_/A la_buf_enable\[44\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_2_1399 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_381 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
X_372_ _372_/A _372_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[84\]_B user_to_mprj_in_gates\[84\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input392_A la_oenb_mprj[103] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input86_A la_data_out_core[59] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[64\]_TE mprj_logic_high_inst/HI[266] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2349 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_193 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_329 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_639_ _639_/Y _639_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA__447__A _447_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[19\] user_to_mprj_in_gates\[19\]/Y input42/X user_to_mprj_in_gates\[19\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_2
XANTENNA_user_to_mprj_in_gates\[75\]_B user_to_mprj_in_gates\[75\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1029 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_buffers\[29\] output777/A user_wb_dat_gates\[29\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_47_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_93 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1019 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[60\]_A user_to_mprj_in_gates\[60\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1169 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__357__A _357_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[66\]_B user_to_mprj_in_gates\[66\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2242 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[87\]_TE mprj_logic_high_inst/HI[289] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1481 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xmprj_dat_buf\[18\] _450_/Y mprj_dat_o_user[18] mprj_dat_buf\[18\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_24_2079 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input238_A la_data_out_mprj[80] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[51\]_A user_to_mprj_in_gates\[51\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input140_A la_data_out_mprj[107] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input405_A la_oenb_mprj[115] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_329 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_424_ _424_/Y _424_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkinv_16
XFILLER_37_1728 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_355_ _355_/Y _355_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
Xuser_to_mprj_in_ena_buf\[121\] vccd vssd user_to_mprj_in_gates\[121\]/B mprj_logic_high_inst/HI[451]
+ input284/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_50_1906 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[57\]_B user_to_mprj_in_gates\[57\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[91\]_A _555_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1813 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[13\] _413_/Y mprj_adr_o_user[13] mprj_adr_buf\[13\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_48_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[127\] user_to_mprj_in_gates\[127\]/Y output657/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_46_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1278 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[93\] user_to_mprj_in_gates\[93\]/Y output747/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_42_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[42\]_A user_to_mprj_in_gates\[42\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput6 input6/X la_data_out_core[101] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_49_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[3\] output781/A user_wb_dat_gates\[3\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_51_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_189 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1683 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[48\]_B user_to_mprj_in_gates\[48\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[82\]_A _546_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__640__A _640_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[0\] user_to_mprj_in_gates\[0\]/Y user_to_mprj_in_gates\[0\]/B
+ input4/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_buffers\[33\]_A user_to_mprj_in_gates\[33\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_613 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_635 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1450 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_57 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[29\] vccd vssd user_to_mprj_in_gates\[29\]/B mprj_logic_high_inst/HI[359]
+ input309/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_42_137 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1761 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[39\]_B user_to_mprj_in_gates\[39\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[123\]_B user_to_mprj_in_gates\[123\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[73\]_A _537_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input188_A la_data_out_mprj[35] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[91\]_B la_buf_enable\[91\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__550__A _550_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input355_A la_iena_mprj[70] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input49_A la_data_out_core[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input522_A mprj_adr_o_core[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[24\]_A user_to_mprj_in_gates\[24\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[112\] la_buf\[112\]/TE _375_/A la_buf_enable\[112\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xla_buf\[97\] _561_/Y la_data_in_core[97] la_buf\[97\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[2\] vccd vssd user_to_mprj_in_gates\[2\]/B mprj_logic_high_inst/HI[332]
+ input310/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_8_1383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2237 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_638 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[127\]_A _591_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_90 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_407_ _407_/A _407_/Y vssd vccd vssd vccd sky130_fd_sc_hd__inv_8
X_338_ _338_/Y _338_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_42_693 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1823 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[114\]_B user_to_mprj_in_gates\[114\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[64\]_A _528_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1260 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1867 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[82\]_B la_buf_enable\[82\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output741_A output741/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__460__A _460_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[86\] user_to_mprj_in_gates\[86\]/Y user_to_mprj_in_gates\[86\]/B
+ input116/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_22_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[15\]_A user_to_mprj_in_gates\[15\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_72 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[23\]_A input565/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2357 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_638 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_137 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__635__A _635_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[118\]_A _582_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_321 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[105\]_B user_to_mprj_in_gates\[105\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[55\]_A _519_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_354 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_376 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[73\]_B la_buf_enable\[73\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__370__A _370_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput616 mprj_sel_o_core[1] _397_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput605 vccd vssd _462_/A mprj_dat_o_core[30] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_25_2196 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[103\]_A_N _366_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[14\]_A input555/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[118\]_A_N _381_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input103_A la_data_out_core[74] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__545__A _545_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[109\]_A _573_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[0\] user_to_mprj_in_gates\[0\]/Y output627/A vccd vssd vssd
+ vccd sky130_fd_sc_hd__clkinv_4
XFILLER_51_490 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[46\]_A _510_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input472_A la_oenb_mprj[60] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[64\]_B la_buf_enable\[64\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[12\] _476_/Y la_data_in_core[12] la_buf\[12\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf\[8\] _472_/Y la_data_in_core[8] la_buf\[8\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_49_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_553 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[5\] _405_/Y mprj_adr_o_user[5] mprj_adr_buf\[5\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_47_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[13\]_TE la_buf\[13\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[56\] user_to_mprj_in_gates\[56\]/Y output706/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_37_1311 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__455__A _455_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output691_A output691/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output789_A output789/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[37\]_A _501_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput31 input31/X la_data_out_core[124] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput20 input20/X la_data_out_core[114] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xuser_wb_dat_gates\[14\] user_wb_dat_gates\[14\]/Y input555/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_50_1533 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput64 input64/X la_data_out_core[39] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput53 input53/X la_data_out_core[29] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput42 vccd vssd input42/X la_data_out_core[19] vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_la_buf_enable\[55\]_B la_buf_enable\[55\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput97 vccd vssd input97/X la_data_out_core[69] vssd vccd sky130_fd_sc_hd__buf_4
Xinput86 vccd vssd input86/X la_data_out_core[59] vssd vccd sky130_fd_sc_hd__buf_4
Xinput75 vccd vssd input75/X la_data_out_core[49] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_48_2141 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_wb_dat_buffers\[11\] output758/A user_wb_dat_gates\[11\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_user_to_mprj_oen_buffers\[122\]_A _385_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[127\]_B mprj_logic_high_inst/HI[457] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1832 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1793 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[112\] user_to_mprj_in_gates\[112\]/Y user_to_mprj_in_gates\[112\]/B
+ input18/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_22_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1729 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_722 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__365__A _365_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[28\]_A _492_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_641 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_696 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[46\]_B la_buf_enable\[46\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[96\] vccd vssd user_to_mprj_in_gates\[96\]/B mprj_logic_high_inst/HI[426]
+ input383/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[113\]_A _376_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[122\] _385_/Y la_oenb_core[122] mprj_logic_high_inst/HI[324]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xmprj_sel_buf\[3\] _399_/Y mprj_sel_o_user[3] mprj_sel_buf\[3\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xinput402 vccd vssd _375_/A la_oenb_mprj[112] vssd vccd sky130_fd_sc_hd__buf_2
Xuser_to_mprj_oen_buffers\[52\] _644_/Y la_oenb_core[52] mprj_logic_high_inst/HI[254]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[118\]_B mprj_logic_high_inst/HI[448] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput446 la_oenb_mprj[37] _629_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput424 vccd vssd _609_/A la_oenb_mprj[17] vssd vccd sky130_fd_sc_hd__buf_2
Xinput435 vccd vssd _619_/A la_oenb_mprj[27] vssd vccd sky130_fd_sc_hd__buf_2
Xinput413 _385_/A la_oenb_mprj[122] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[74\] la_buf\[74\]/TE _337_/A la_buf_enable\[74\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xinput457 vccd vssd _639_/A la_oenb_mprj[47] vssd vccd sky130_fd_sc_hd__buf_4
Xinput468 la_oenb_mprj[57] _649_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput479 vccd vssd _330_/A la_oenb_mprj[67] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_40_1757 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[36\]_TE la_buf\[36\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input318_A la_iena_mprj[37] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input220_A la_data_out_mprj[64] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_449 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[1\]_A_N _593_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[19\]_A _483_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1951 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[37\]_B la_buf_enable\[37\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_667 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[116\] _580_/Y la_data_in_core[116] la_buf\[116\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[6\]_A input354/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[104\]_A _367_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1613 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1602 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_clk2_buf_A _392_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[109\]_B mprj_logic_high_inst/HI[439] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1117 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_538 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1933 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output704_A output704/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1999 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[49\] user_to_mprj_in_gates\[49\]/Y user_to_mprj_in_gates\[49\]/B
+ input75/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_50_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[40\]_B mprj_logic_high_inst/HI[370] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_50_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[4\]_TE la_buf\[4\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[28\]_B la_buf_enable\[28\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[30\]_A _622_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1833 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[59\]_TE la_buf\[59\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1719 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1504 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2238 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1548 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_585 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[97\]_A _360_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[11\] vccd vssd user_to_mprj_in_gates\[11\]/B mprj_logic_high_inst/HI[341]
+ input282/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_43_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[31\]_B mprj_logic_high_inst/HI[361] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[19\]_B la_buf_enable\[19\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1001 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input170_A la_data_out_mprj[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[21\]_A _613_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2011 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input268_A la_iena_mprj[107] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[98\]_B mprj_logic_high_inst/HI[428] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput210 la_data_out_mprj[55] _519_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_input435_A la_oenb_mprj[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input31_A la_data_out_core[124] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput221 la_data_out_mprj[65] _529_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput232 vccd vssd _539_/A la_data_out_mprj[75] vssd vccd sky130_fd_sc_hd__buf_2
Xinput243 _549_/A la_data_out_mprj[85] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput254 vccd vssd _559_/A la_data_out_mprj[95] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_48_357 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xinput265 vssd vccd input265/X la_iena_mprj[104] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput276 vssd vccd input276/X la_iena_mprj[114] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput287 vssd vccd input287/X la_iena_mprj[124] vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_input602_A mprj_dat_o_core[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput298 vssd vccd input298/X la_iena_mprj[19] vssd vccd sky130_fd_sc_hd__clkbuf_1
X_655_ _655_/A _655_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[88\]_A _351_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_586_ _586_/A _586_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_16_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_257 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[22\]_B mprj_logic_high_inst/HI[352] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_9_910 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1071 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[19\] user_to_mprj_in_gates\[19\]/Y output665/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output654_A output654/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput706 vccd vssd la_data_in_mprj[56] output706/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput717 vccd vssd la_data_in_mprj[66] output717/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_oen_buffers\[12\]_A _604_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput728 vccd vssd la_data_in_mprj[76] output728/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput739 vccd vssd la_data_in_mprj[86] output739/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_45_2133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[89\]_B mprj_logic_high_inst/HI[419] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1730 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[79\]_A _342_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1225 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[13\]_B mprj_logic_high_inst/HI[343] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA__643__A _643_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1881 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[6\]_A input578/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[61\]_A_N _653_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1778 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1199 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[76\]_A_N _339_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1841 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_79 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[59\] vccd vssd user_to_mprj_in_gates\[59\]/B mprj_logic_high_inst/HI[389]
+ input342/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_6_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[6\]_A input98/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1312 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[0\]_B user_irq_ena_buf\[0\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_440_ _440_/A _440_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
X_371_ _371_/A _371_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[15\] _607_/Y la_oenb_core[15] mprj_logic_high_inst/HI[217]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[37\] la_buf\[37\]/TE _629_/A la_buf_enable\[37\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf_enable\[14\]_A_N _606_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__553__A _553_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1921 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input385_A la_iena_mprj[98] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[29\]_A_N _621_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input79_A la_data_out_core[52] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input552_A mprj_dat_i_user[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1449 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1201 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_638_ _638_/Y _638_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_533 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_569_ _569_/Y _569_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA__463__A _463_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output771_A output771/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__638__A _638_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1582 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1022 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[30\]_A _462_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1077 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_739 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__373__A _373_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1597 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_448 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input133_A la_data_out_mprj[100] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__548__A _548_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input300_A la_iena_mprj[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_423_ _423_/A _423_/Y vssd vccd vssd vccd sky130_fd_sc_hd__inv_8
XFILLER_35_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[21\]_A _453_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_385 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[42\] _506_/Y la_data_in_core[42] la_buf\[42\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_354_ _354_/Y _354_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_50_1918 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[114\] vccd vssd user_to_mprj_in_gates\[114\]/B mprj_logic_high_inst/HI[444]
+ input276/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[31\]_TE mprj_logic_high_inst/HI[233] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_721 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_242 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2261 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1869 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1307 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_441 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput7 vccd vssd input7/X la_data_out_core[102] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_49_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[86\] user_to_mprj_in_gates\[86\]/Y output739/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_36_124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__458__A _458_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[107\]_TE la_buf\[107\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_831 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[31\] user_to_mprj_in_gates\[31\]/Y user_to_mprj_in_gates\[31\]/B
+ input56/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_53_2232 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[12\]_A _444_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_897 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1564 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1895 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1873 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[6\]_TE mprj_adr_buf\[6\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1313 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2069 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__368__A _368_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_669 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[7\]_A _599_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[10\]_A user_wb_dat_gates\[10\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[54\]_TE mprj_logic_high_inst/HI[256] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_503 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_529 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1924 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[82\] _345_/Y la_oenb_core[82] mprj_logic_high_inst/HI[284]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_2_223 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xmprj_dat_buf\[30\] _462_/Y mprj_dat_o_user[30] mprj_dat_buf\[30\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_4_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input250_A la_data_out_mprj[91] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input348_A la_iena_mprj[64] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input515_A la_oenb_mprj[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1395 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[105\] la_buf\[105\]/TE _368_/A la_buf_enable\[105\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_33_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1559 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_91 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_80 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_406_ _406_/Y _406_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkinv_8
X_337_ _337_/Y _337_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_41_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1272 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output734_A output734/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1699 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[79\] user_to_mprj_in_gates\[79\]/Y user_to_mprj_in_gates\[79\]/B
+ input108/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_la_buf\[92\]_TE la_buf\[92\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[23\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[77\]_TE mprj_logic_high_inst/HI[279] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_617 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2002 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__651__A _651_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput617 mprj_sel_o_core[2] _398_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_5_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput606 mprj_dat_o_core[31] _463_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_21_2006 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[14\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[41\] vccd vssd user_to_mprj_in_gates\[41\]/B mprj_logic_high_inst/HI[371]
+ input323/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_44_937 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_cyc_buf_TE mprj_cyc_buf/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input298_A la_iena_mprj[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__561__A _561_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input61_A la_data_out_core[36] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input465_A la_oenb_mprj[54] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1953 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1023 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_403 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1323 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[49\] user_to_mprj_in_gates\[49\]/Y output698/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_50_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output684_A output684/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput21 input21/X la_data_out_core[115] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput10 vccd vssd input10/X la_data_out_core[105] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_15_1643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput32 input32/X la_data_out_core[125] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput43 vccd vssd input43/X la_data_out_core[1] vssd vccd sky130_fd_sc_hd__buf_4
Xinput54 vccd vssd input54/X la_data_out_core[2] vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA__471__A _471_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput98 input98/X la_data_out_core[6] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput87 vccd vssd input87/X la_data_out_core[5] vssd vccd sky130_fd_sc_hd__buf_2
Xinput76 input76/X la_data_out_core[4] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput65 input65/X la_data_out_core[3] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1844 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1073 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[105\] user_to_mprj_in_gates\[105\]/Y user_to_mprj_in_gates\[105\]/B
+ input10/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_53_767 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_233 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__646__A _646_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj2_logic_high_inst mprj2_pwrgood/A vccd2 vssd2 mprj2_logic_high
XANTENNA_mprj_adr_buf\[6\]_A _406_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__381__A _381_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[89\] vccd vssd user_to_mprj_in_gates\[89\]/B mprj_logic_high_inst/HI[419]
+ input375/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_7_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[115\] _378_/Y la_oenb_core[115] mprj_logic_high_inst/HI[317]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xinput403 _376_/A la_oenb_mprj[113] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput425 la_oenb_mprj[18] _610_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput436 _620_/A la_oenb_mprj[28] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput414 _386_/A la_oenb_mprj[123] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput458 vccd vssd _640_/A la_oenb_mprj[48] vssd vccd sky130_fd_sc_hd__buf_2
Xinput447 la_oenb_mprj[38] _630_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput469 vccd vssd _650_/A la_oenb_mprj[58] vssd vccd sky130_fd_sc_hd__buf_2
Xuser_to_mprj_oen_buffers\[45\] _637_/Y la_oenb_core[45] mprj_logic_high_inst/HI[247]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[67\] la_buf\[67\]/TE _330_/A la_buf_enable\[67\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_29_742 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input213_A la_data_out_mprj[58] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1229 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__556__A _556_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input582_A mprj_dat_o_core[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1963 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1865 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_rstn_buf_TE mprj_rstn_buf/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[6\]_B mprj_logic_high_inst/HI[336] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[109\] _573_/Y la_data_in_core[109] la_buf\[109\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_2061 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[102\] user_to_mprj_in_gates\[102\]/Y output630/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_43_1393 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__466__A _466_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1730 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1738 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[102\]_A_N _365_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[117\]_A_N _380_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[127\]_B la_buf_enable\[127\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[1\] _433_/Y mprj_dat_o_user[1] mprj_dat_buf\[1\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xmprj_logic_high_inst mprj_rstn_buf/TE la_buf_enable\[26\]/B la_buf_enable\[27\]/B
+ la_buf_enable\[28\]/B la_buf_enable\[29\]/B la_buf_enable\[30\]/B la_buf_enable\[31\]/B
+ la_buf_enable\[32\]/B la_buf_enable\[33\]/B la_buf_enable\[34\]/B la_buf_enable\[35\]/B
+ mprj_adr_buf\[0\]/TE la_buf_enable\[36\]/B la_buf_enable\[37\]/B la_buf_enable\[38\]/B
+ la_buf_enable\[39\]/B la_buf_enable\[40\]/B la_buf_enable\[41\]/B la_buf_enable\[42\]/B
+ la_buf_enable\[43\]/B la_buf_enable\[44\]/B la_buf_enable\[45\]/B mprj_adr_buf\[1\]/TE
+ la_buf_enable\[46\]/B la_buf_enable\[47\]/B la_buf_enable\[48\]/B la_buf_enable\[49\]/B
+ la_buf_enable\[50\]/B la_buf_enable\[51\]/B la_buf_enable\[52\]/B la_buf_enable\[53\]/B
+ la_buf_enable\[54\]/B la_buf_enable\[55\]/B mprj_adr_buf\[2\]/TE la_buf_enable\[56\]/B
+ la_buf_enable\[57\]/B la_buf_enable\[58\]/B la_buf_enable\[59\]/B la_buf_enable\[60\]/B
+ la_buf_enable\[61\]/B la_buf_enable\[62\]/B la_buf_enable\[63\]/B la_buf_enable\[64\]/B
+ la_buf_enable\[65\]/B mprj_adr_buf\[3\]/TE la_buf_enable\[66\]/B la_buf_enable\[67\]/B
+ la_buf_enable\[68\]/B la_buf_enable\[69\]/B la_buf_enable\[70\]/B la_buf_enable\[71\]/B
+ la_buf_enable\[72\]/B la_buf_enable\[73\]/B la_buf_enable\[74\]/B la_buf_enable\[75\]/B
+ mprj_adr_buf\[4\]/TE la_buf_enable\[76\]/B la_buf_enable\[77\]/B la_buf_enable\[78\]/B
+ la_buf_enable\[79\]/B la_buf_enable\[80\]/B la_buf_enable\[81\]/B la_buf_enable\[82\]/B
+ la_buf_enable\[83\]/B la_buf_enable\[84\]/B la_buf_enable\[85\]/B mprj_adr_buf\[5\]/TE
+ la_buf_enable\[86\]/B la_buf_enable\[87\]/B la_buf_enable\[88\]/B la_buf_enable\[89\]/B
+ la_buf_enable\[90\]/B la_buf_enable\[91\]/B la_buf_enable\[92\]/B la_buf_enable\[93\]/B
+ la_buf_enable\[94\]/B la_buf_enable\[95\]/B mprj_adr_buf\[6\]/TE la_buf_enable\[96\]/B
+ la_buf_enable\[97\]/B la_buf_enable\[98\]/B la_buf_enable\[99\]/B la_buf_enable\[100\]/B
+ la_buf_enable\[101\]/B la_buf_enable\[102\]/B la_buf_enable\[103\]/B la_buf_enable\[104\]/B
+ la_buf_enable\[105\]/B mprj_adr_buf\[7\]/TE la_buf_enable\[106\]/B la_buf_enable\[107\]/B
+ la_buf_enable\[108\]/B la_buf_enable\[109\]/B la_buf_enable\[110\]/B la_buf_enable\[111\]/B
+ la_buf_enable\[112\]/B la_buf_enable\[113\]/B la_buf_enable\[114\]/B la_buf_enable\[115\]/B
+ mprj_adr_buf\[8\]/TE la_buf_enable\[116\]/B la_buf_enable\[117\]/B la_buf_enable\[118\]/B
+ la_buf_enable\[119\]/B la_buf_enable\[120\]/B la_buf_enable\[121\]/B la_buf_enable\[122\]/B
+ la_buf_enable\[123\]/B la_buf_enable\[124\]/B la_buf_enable\[125\]/B mprj_adr_buf\[9\]/TE
+ mprj_clk_buf/TE la_buf_enable\[126\]/B la_buf_enable\[127\]/B mprj_logic_high_inst/HI[202]
+ mprj_logic_high_inst/HI[203] mprj_logic_high_inst/HI[204] mprj_logic_high_inst/HI[205]
+ mprj_logic_high_inst/HI[206] mprj_logic_high_inst/HI[207] mprj_logic_high_inst/HI[208]
+ mprj_logic_high_inst/HI[209] mprj_adr_buf\[10\]/TE mprj_logic_high_inst/HI[210]
+ mprj_logic_high_inst/HI[211] mprj_logic_high_inst/HI[212] mprj_logic_high_inst/HI[213]
+ mprj_logic_high_inst/HI[214] mprj_logic_high_inst/HI[215] mprj_logic_high_inst/HI[216]
+ mprj_logic_high_inst/HI[217] mprj_logic_high_inst/HI[218] mprj_logic_high_inst/HI[219]
+ mprj_adr_buf\[11\]/TE mprj_logic_high_inst/HI[220] mprj_logic_high_inst/HI[221]
+ mprj_logic_high_inst/HI[222] mprj_logic_high_inst/HI[223] mprj_logic_high_inst/HI[224]
+ mprj_logic_high_inst/HI[225] mprj_logic_high_inst/HI[226] mprj_logic_high_inst/HI[227]
+ mprj_logic_high_inst/HI[228] mprj_logic_high_inst/HI[229] mprj_adr_buf\[12\]/TE
+ mprj_logic_high_inst/HI[230] mprj_logic_high_inst/HI[231] mprj_logic_high_inst/HI[232]
+ mprj_logic_high_inst/HI[233] mprj_logic_high_inst/HI[234] mprj_logic_high_inst/HI[235]
+ mprj_logic_high_inst/HI[236] mprj_logic_high_inst/HI[237] mprj_logic_high_inst/HI[238]
+ mprj_logic_high_inst/HI[239] mprj_adr_buf\[13\]/TE mprj_logic_high_inst/HI[240]
+ mprj_logic_high_inst/HI[241] mprj_logic_high_inst/HI[242] mprj_logic_high_inst/HI[243]
+ mprj_logic_high_inst/HI[244] mprj_logic_high_inst/HI[245] mprj_logic_high_inst/HI[246]
+ mprj_logic_high_inst/HI[247] mprj_logic_high_inst/HI[248] mprj_logic_high_inst/HI[249]
+ mprj_adr_buf\[14\]/TE mprj_logic_high_inst/HI[250] mprj_logic_high_inst/HI[251]
+ mprj_logic_high_inst/HI[252] mprj_logic_high_inst/HI[253] mprj_logic_high_inst/HI[254]
+ mprj_logic_high_inst/HI[255] mprj_logic_high_inst/HI[256] mprj_logic_high_inst/HI[257]
+ mprj_logic_high_inst/HI[258] mprj_logic_high_inst/HI[259] mprj_adr_buf\[15\]/TE
+ mprj_logic_high_inst/HI[260] mprj_logic_high_inst/HI[261] mprj_logic_high_inst/HI[262]
+ mprj_logic_high_inst/HI[263] mprj_logic_high_inst/HI[264] mprj_logic_high_inst/HI[265]
+ mprj_logic_high_inst/HI[266] mprj_logic_high_inst/HI[267] mprj_logic_high_inst/HI[268]
+ mprj_logic_high_inst/HI[269] mprj_adr_buf\[16\]/TE mprj_logic_high_inst/HI[270]
+ mprj_logic_high_inst/HI[271] mprj_logic_high_inst/HI[272] mprj_logic_high_inst/HI[273]
+ mprj_logic_high_inst/HI[274] mprj_logic_high_inst/HI[275] mprj_logic_high_inst/HI[276]
+ mprj_logic_high_inst/HI[277] mprj_logic_high_inst/HI[278] mprj_logic_high_inst/HI[279]
+ mprj_adr_buf\[17\]/TE mprj_logic_high_inst/HI[280] mprj_logic_high_inst/HI[281]
+ mprj_logic_high_inst/HI[282] mprj_logic_high_inst/HI[283] mprj_logic_high_inst/HI[284]
+ mprj_logic_high_inst/HI[285] mprj_logic_high_inst/HI[286] mprj_logic_high_inst/HI[288]
+ mprj_logic_high_inst/HI[289] mprj_adr_buf\[18\]/TE mprj_logic_high_inst/HI[290]
+ mprj_logic_high_inst/HI[291] mprj_logic_high_inst/HI[292] mprj_logic_high_inst/HI[293]
+ mprj_logic_high_inst/HI[294] mprj_logic_high_inst/HI[295] mprj_logic_high_inst/HI[296]
+ mprj_logic_high_inst/HI[297] mprj_logic_high_inst/HI[298] mprj_logic_high_inst/HI[299]
+ mprj_adr_buf\[19\]/TE mprj_clk2_buf/TE mprj_logic_high_inst/HI[300] mprj_logic_high_inst/HI[301]
+ mprj_logic_high_inst/HI[302] mprj_logic_high_inst/HI[303] mprj_logic_high_inst/HI[304]
+ mprj_logic_high_inst/HI[305] mprj_logic_high_inst/HI[306] mprj_logic_high_inst/HI[307]
+ mprj_logic_high_inst/HI[308] mprj_logic_high_inst/HI[309] mprj_adr_buf\[20\]/TE
+ mprj_logic_high_inst/HI[310] mprj_logic_high_inst/HI[311] mprj_logic_high_inst/HI[312]
+ mprj_logic_high_inst/HI[313] mprj_logic_high_inst/HI[314] mprj_logic_high_inst/HI[315]
+ mprj_logic_high_inst/HI[316] mprj_logic_high_inst/HI[317] mprj_logic_high_inst/HI[318]
+ mprj_logic_high_inst/HI[319] mprj_adr_buf\[21\]/TE mprj_logic_high_inst/HI[320]
+ mprj_logic_high_inst/HI[321] mprj_logic_high_inst/HI[322] mprj_logic_high_inst/HI[323]
+ mprj_logic_high_inst/HI[324] mprj_logic_high_inst/HI[325] mprj_logic_high_inst/HI[326]
+ mprj_logic_high_inst/HI[327] mprj_logic_high_inst/HI[328] mprj_logic_high_inst/HI[329]
+ mprj_adr_buf\[22\]/TE mprj_logic_high_inst/HI[330] mprj_logic_high_inst/HI[331]
+ mprj_logic_high_inst/HI[332] mprj_logic_high_inst/HI[333] mprj_logic_high_inst/HI[334]
+ mprj_logic_high_inst/HI[335] mprj_logic_high_inst/HI[336] mprj_logic_high_inst/HI[337]
+ mprj_logic_high_inst/HI[338] mprj_logic_high_inst/HI[339] mprj_adr_buf\[23\]/TE
+ mprj_logic_high_inst/HI[340] mprj_logic_high_inst/HI[341] mprj_logic_high_inst/HI[342]
+ mprj_logic_high_inst/HI[343] mprj_logic_high_inst/HI[344] mprj_logic_high_inst/HI[345]
+ mprj_logic_high_inst/HI[346] mprj_logic_high_inst/HI[347] mprj_logic_high_inst/HI[348]
+ mprj_logic_high_inst/HI[349] mprj_adr_buf\[24\]/TE mprj_logic_high_inst/HI[350]
+ mprj_logic_high_inst/HI[351] mprj_logic_high_inst/HI[352] mprj_logic_high_inst/HI[353]
+ mprj_logic_high_inst/HI[354] mprj_logic_high_inst/HI[355] mprj_logic_high_inst/HI[356]
+ mprj_logic_high_inst/HI[357] mprj_logic_high_inst/HI[358] mprj_logic_high_inst/HI[359]
+ mprj_adr_buf\[25\]/TE mprj_logic_high_inst/HI[360] mprj_logic_high_inst/HI[361]
+ mprj_logic_high_inst/HI[362] mprj_logic_high_inst/HI[363] mprj_logic_high_inst/HI[364]
+ mprj_logic_high_inst/HI[365] mprj_logic_high_inst/HI[366] mprj_logic_high_inst/HI[367]
+ mprj_logic_high_inst/HI[368] mprj_logic_high_inst/HI[369] mprj_adr_buf\[26\]/TE
+ mprj_logic_high_inst/HI[370] mprj_logic_high_inst/HI[371] mprj_logic_high_inst/HI[372]
+ mprj_logic_high_inst/HI[373] mprj_logic_high_inst/HI[374] mprj_logic_high_inst/HI[375]
+ mprj_logic_high_inst/HI[376] mprj_logic_high_inst/HI[377] mprj_logic_high_inst/HI[378]
+ mprj_logic_high_inst/HI[379] mprj_adr_buf\[27\]/TE mprj_logic_high_inst/HI[380]
+ mprj_logic_high_inst/HI[381] mprj_logic_high_inst/HI[382] mprj_logic_high_inst/HI[383]
+ mprj_logic_high_inst/HI[384] mprj_logic_high_inst/HI[385] mprj_logic_high_inst/HI[386]
+ mprj_logic_high_inst/HI[387] mprj_logic_high_inst/HI[388] mprj_logic_high_inst/HI[389]
+ mprj_adr_buf\[28\]/TE mprj_logic_high_inst/HI[390] mprj_logic_high_inst/HI[391]
+ mprj_logic_high_inst/HI[392] mprj_logic_high_inst/HI[393] mprj_logic_high_inst/HI[394]
+ mprj_logic_high_inst/HI[395] mprj_logic_high_inst/HI[396] mprj_logic_high_inst/HI[397]
+ mprj_logic_high_inst/HI[398] mprj_logic_high_inst/HI[399] mprj_adr_buf\[29\]/TE
+ mprj_cyc_buf/TE mprj_logic_high_inst/HI[400] mprj_logic_high_inst/HI[401] mprj_logic_high_inst/HI[402]
+ mprj_logic_high_inst/HI[403] mprj_logic_high_inst/HI[404] mprj_logic_high_inst/HI[405]
+ mprj_logic_high_inst/HI[406] mprj_logic_high_inst/HI[407] mprj_logic_high_inst/HI[408]
+ mprj_logic_high_inst/HI[409] mprj_adr_buf\[30\]/TE mprj_logic_high_inst/HI[410]
+ mprj_logic_high_inst/HI[411] mprj_logic_high_inst/HI[412] mprj_logic_high_inst/HI[413]
+ mprj_logic_high_inst/HI[414] mprj_logic_high_inst/HI[415] mprj_logic_high_inst/HI[416]
+ mprj_logic_high_inst/HI[417] mprj_logic_high_inst/HI[418] mprj_logic_high_inst/HI[419]
+ mprj_adr_buf\[31\]/TE mprj_logic_high_inst/HI[420] mprj_logic_high_inst/HI[421]
+ mprj_logic_high_inst/HI[422] mprj_logic_high_inst/HI[423] mprj_logic_high_inst/HI[424]
+ mprj_logic_high_inst/HI[425] mprj_logic_high_inst/HI[426] mprj_logic_high_inst/HI[427]
+ mprj_logic_high_inst/HI[428] mprj_dat_buf\[0\]/TE mprj_logic_high_inst/HI[430] mprj_logic_high_inst/HI[431]
+ mprj_logic_high_inst/HI[432] mprj_logic_high_inst/HI[433] mprj_logic_high_inst/HI[434]
+ mprj_logic_high_inst/HI[435] mprj_logic_high_inst/HI[436] mprj_logic_high_inst/HI[437]
+ mprj_logic_high_inst/HI[438] mprj_logic_high_inst/HI[439] mprj_dat_buf\[1\]/TE mprj_logic_high_inst/HI[440]
+ mprj_logic_high_inst/HI[441] mprj_logic_high_inst/HI[442] mprj_logic_high_inst/HI[443]
+ mprj_logic_high_inst/HI[444] mprj_logic_high_inst/HI[445] mprj_logic_high_inst/HI[446]
+ mprj_logic_high_inst/HI[447] mprj_logic_high_inst/HI[448] mprj_logic_high_inst/HI[449]
+ mprj_dat_buf\[2\]/TE mprj_logic_high_inst/HI[450] mprj_logic_high_inst/HI[451] mprj_logic_high_inst/HI[452]
+ mprj_logic_high_inst/HI[453] mprj_logic_high_inst/HI[454] mprj_logic_high_inst/HI[455]
+ mprj_logic_high_inst/HI[456] mprj_logic_high_inst/HI[457] user_irq_ena_buf\[0\]/B
+ user_irq_ena_buf\[1\]/B mprj_dat_buf\[3\]/TE user_irq_ena_buf\[2\]/B mprj_pwrgood/A
+ user_to_mprj_wb_ena_buf/B mprj_dat_buf\[4\]/TE mprj_dat_buf\[5\]/TE mprj_dat_buf\[6\]/TE
+ mprj_dat_buf\[7\]/TE mprj_stb_buf/TE mprj_dat_buf\[8\]/TE mprj_dat_buf\[9\]/TE mprj_dat_buf\[10\]/TE
+ mprj_dat_buf\[11\]/TE mprj_dat_buf\[12\]/TE mprj_dat_buf\[13\]/TE mprj_dat_buf\[14\]/TE
+ mprj_dat_buf\[15\]/TE mprj_dat_buf\[16\]/TE mprj_dat_buf\[17\]/TE mprj_we_buf/TE
+ mprj_dat_buf\[18\]/TE mprj_dat_buf\[19\]/TE mprj_dat_buf\[20\]/TE mprj_dat_buf\[21\]/TE
+ mprj_dat_buf\[22\]/TE mprj_dat_buf\[23\]/TE mprj_dat_buf\[24\]/TE mprj_dat_buf\[25\]/TE
+ mprj_dat_buf\[26\]/TE mprj_dat_buf\[27\]/TE mprj_sel_buf\[0\]/TE mprj_dat_buf\[28\]/TE
+ mprj_dat_buf\[29\]/TE mprj_dat_buf\[30\]/TE mprj_dat_buf\[31\]/TE la_buf_enable\[0\]/B
+ la_buf_enable\[1\]/B la_buf_enable\[2\]/B la_buf_enable\[3\]/B la_buf_enable\[4\]/B
+ la_buf_enable\[5\]/B mprj_sel_buf\[1\]/TE la_buf_enable\[6\]/B la_buf_enable\[7\]/B
+ la_buf_enable\[8\]/B la_buf_enable\[9\]/B la_buf_enable\[10\]/B la_buf_enable\[11\]/B
+ la_buf_enable\[12\]/B la_buf_enable\[13\]/B la_buf_enable\[14\]/B la_buf_enable\[15\]/B
+ mprj_sel_buf\[2\]/TE la_buf_enable\[16\]/B la_buf_enable\[17\]/B la_buf_enable\[18\]/B
+ la_buf_enable\[19\]/B la_buf_enable\[20\]/B la_buf_enable\[21\]/B la_buf_enable\[22\]/B
+ la_buf_enable\[23\]/B la_buf_enable\[24\]/B la_buf_enable\[25\]/B mprj_sel_buf\[3\]/TE
+ vccd1 mprj_logic_high_inst/HI[287] mprj_logic_high_inst/HI[429] vssd1 mprj_logic_high
XFILLER_26_1591 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1516 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__376__A _376_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_A input127/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_605 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1860 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1057 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input163_A la_data_out_mprj[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2201 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[118\]_B la_buf_enable\[118\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[20\]_A input44/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput211 la_data_out_mprj[56] _520_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput200 la_data_out_mprj[46] _510_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_46_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input330_A la_iena_mprj[48] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input428_A la_oenb_mprj[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput222 la_data_out_mprj[66] _530_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput233 _540_/A la_data_out_mprj[76] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput244 _550_/A la_data_out_mprj[86] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_input24_A la_data_out_core[118] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput255 la_data_out_mprj[96] _560_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput266 vssd vccd input266/X la_iena_mprj[105] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput277 vssd vccd input277/X la_iena_mprj[115] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput288 vssd vccd input288/X la_iena_mprj[125] vssd vccd sky130_fd_sc_hd__clkbuf_1
X_654_ _654_/Y _654_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_29_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput299 vssd vccd input299/X la_iena_mprj[1] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1173 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[72\] _536_/Y la_data_in_core[72] la_buf\[72\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_40_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_585_ _585_/A _585_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_user_wb_dat_buffers\[9\]_A user_wb_dat_gates\[9\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[87\]_A input117/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_792 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1673 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1083 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput707 vccd vssd la_data_in_mprj[57] output707/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput718 vccd vssd la_data_in_mprj[67] output718/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput729 vccd vssd la_data_in_mprj[77] output729/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_output647_A output647/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_693 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[109\]_B la_buf_enable\[109\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[11\]_A input26/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1742 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[61\] user_to_mprj_in_gates\[61\]/Y user_to_mprj_in_gates\[61\]/B
+ input89/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_7_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[78\]_A input107/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[6\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1757 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[26\]_TE la_buf\[26\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2321 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1653 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[0\]_A_N _592_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_2207 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1697 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2150 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1747 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_807 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2058 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[6\]_B user_to_mprj_in_gates\[6\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1897 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_564 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_370_ _370_/A _370_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_39_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[69\]_A input97/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1911 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_903 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input280_A la_iena_mprj[118] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1392 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input378_A la_iena_mprj[91] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1999 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input545_A mprj_adr_o_core[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1753 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_133 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1257 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1904 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2097 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_637_ _637_/A _637_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
X_568_ _568_/Y _568_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf\[49\]_TE la_buf\[49\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[31\] user_to_mprj_in_gates\[31\]/Y output679/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
X_499_ _499_/Y _499_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_51_2160 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output764_A output764/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1951 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_807 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1594 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1034 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__654__A _654_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_427 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1016 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2151 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[71\] vccd vssd user_to_mprj_in_gates\[71\]/B mprj_logic_high_inst/HI[401]
+ input356/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_49_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2059 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input126_A la_data_out_core[95] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_637 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_422_ _422_/Y _422_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_6
XFILLER_39_2291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__564__A _564_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[126\]_A input33/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_353_ _353_/Y _353_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input495_A la_oenb_mprj[81] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input91_A la_data_out_core[63] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[35\] _499_/Y la_data_in_core[35] la_buf\[35\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[107\] vccd vssd user_to_mprj_in_gates\[107\]/B mprj_logic_high_inst/HI[437]
+ input268/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_10_751 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[7\] input579/X user_wb_ack_gate/B user_wb_dat_gates\[7\]/Y vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_8
XFILLER_5_221 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_254 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput8 vccd vssd input8/X la_data_out_core[103] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_7_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_497 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1870 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1723 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[79\] user_to_mprj_in_gates\[79\]/Y output731/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_la_buf_enable\[60\]_A_N _652_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__474__A _474_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[117\]_A input23/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[24\] user_to_mprj_in_gates\[24\]/Y user_to_mprj_in_gates\[24\]/B
+ input48/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_la_buf_enable\[75\]_A_N _338_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[13\]_A_N _605_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_2335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__649__A _649_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1981 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[28\]_A_N _620_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1474 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__384__A _384_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[108\]_A input13/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2317 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2085 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1936 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[75\] _338_/Y la_oenb_core[75] mprj_logic_high_inst/HI[277]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_2_235 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[97\] vccd vssd la_buf\[97\]/TE la_buf_enable\[97\]/B _360_/A vssd
+ vccd sky130_fd_sc_hd__and2b_2
XFILLER_2_279 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1892 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xmprj_dat_buf\[23\] _455_/Y mprj_dat_o_user[23] mprj_dat_buf\[23\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input243_A la_data_out_mprj[85] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1756 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__559__A _559_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_946 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input410_A la_oenb_mprj[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input508_A la_oenb_mprj[93] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_150 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_92 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_81 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_70 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_405_ _405_/Y _405_/A vssd vccd vssd vccd sky130_fd_sc_hd__inv_16
X_336_ _336_/Y _336_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_30_824 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1983 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1705 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1284 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1645 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1033 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1689 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output727_A output727/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1138 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__469__A _469_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[122\]_TE mprj_logic_high_inst/HI[324] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_63 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1761 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1772 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[70\]_A input355/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_183 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[6\]_B la_buf_enable\[6\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[3\] la_buf\[3\]/TE _595_/A la_buf_enable\[3\]/B vssd vccd vssd vccd
+ sky130_fd_sc_hd__and2b_1
XFILLER_21_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1693 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput607 vccd vssd _435_/A mprj_dat_o_core[3] vssd vccd sky130_fd_sc_hd__buf_2
Xinput618 mprj_sel_o_core[3] _399_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA__379__A _379_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2237 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[21\]_TE mprj_logic_high_inst/HI[223] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_445 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[34\] vccd vssd user_to_mprj_in_gates\[34\]/B mprj_logic_high_inst/HI[364]
+ input315/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_ena_buf\[61\]_A input345/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1869 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2125 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_150 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_305 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[12\] la_buf\[12\]/TE _604_/A la_buf_enable\[12\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_32_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input193_A la_data_out_mprj[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_839 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_378 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1468 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input360_A la_iena_mprj[75] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input458_A la_oenb_mprj[48] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input54_A la_data_out_core[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input625_A user_irq_ena[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_721 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_445 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2003 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xpowergood_check mprj2_vdd_pwrgood/A mprj_vdd_pwrgood/A vccd vssd vdda1 vdda2 dw_193520_8662#
+ vssa1 dw_201140_8600# vssa2 mgmt_protect_hv
XFILLER_34_448 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[52\]_A input335/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1978 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1335 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output677_A output677/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput22 input22/X la_data_out_core[116] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput11 vccd vssd input11/X la_data_out_core[106] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_15_1655 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xinput33 input33/X la_data_out_core[126] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput55 vccd vssd input55/X la_data_out_core[30] vssd vccd sky130_fd_sc_hd__buf_4
Xinput44 input44/X la_data_out_core[20] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_15_1699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput88 input88/X la_data_out_core[60] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput77 vccd vssd input77/X la_data_out_core[50] vssd vccd sky130_fd_sc_hd__buf_4
Xinput66 input66/X la_data_out_core[40] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput99 vccd vssd input99/X la_data_out_core[70] vssd vccd sky130_fd_sc_hd__buf_4
Xuser_to_mprj_in_gates\[91\] user_to_mprj_in_gates\[91\]/Y user_to_mprj_in_gates\[91\]/B
+ input122/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_48_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[44\]_TE mprj_logic_high_inst/HI[246] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[0\]_A _396_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[43\]_A input325/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_278 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1007 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2227 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput426 la_oenb_mprj[19] _611_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput437 vccd vssd _621_/A la_oenb_mprj[29] vssd vccd sky130_fd_sc_hd__buf_2
Xinput404 _377_/A la_oenb_mprj[114] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput415 _387_/A la_oenb_mprj[124] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xuser_to_mprj_oen_buffers\[108\] _371_/Y la_oenb_core[108] mprj_logic_high_inst/HI[310]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xinput459 _641_/A la_oenb_mprj[49] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput448 vccd vssd la_oenb_mprj[39] _631_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_754 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1208 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[38\] _630_/Y la_oenb_core[38] mprj_logic_high_inst/HI[240]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2209 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input206_A la_data_out_mprj[51] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[34\]_A input315/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1390 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1221 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__572__A _572_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input575_A mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[82\]_TE la_buf\[82\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[1\]_A _433_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[67\]_TE mprj_logic_high_inst/HI[269] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_529 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_253 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_297 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[61\] output712/A user_to_mprj_in_gates\[61\]/Y vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_output794_A output794/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[25\]_A input305/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_749 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1619 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1165 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2066 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__482__A _482_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1365 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[31\]_TE mprj_dat_buf\[31\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1283 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[90\]_A user_to_mprj_in_gates\[90\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2207 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__657__A _657_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[16\]_A input295/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_B user_to_mprj_in_gates\[96\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__392__A _392_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2297 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[20\]_B user_to_mprj_in_gates\[20\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput201 la_data_out_mprj[47] _511_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_buffers\[81\]_A user_to_mprj_in_gates\[81\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input156_A la_data_out_mprj[121] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput212 la_data_out_mprj[57] _521_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput223 la_data_out_mprj[67] _531_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput234 la_data_out_mprj[77] _541_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput245 la_data_out_mprj[87] _551_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1512 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input323_A la_iena_mprj[41] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput256 vccd vssd _561_/A la_data_out_mprj[97] vssd vccd sky130_fd_sc_hd__buf_2
Xinput267 vssd vccd input267/X la_iena_mprj[106] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput278 vssd vccd input278/X la_iena_mprj[116] vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_input17_A la_data_out_core[111] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_653_ _653_/A _653_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
Xinput289 vssd vccd input289/X la_iena_mprj[126] vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA__567__A _567_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1589 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_584_ _584_/Y _584_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf\[65\] _529_/Y la_data_in_core[65] la_buf\[65\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_565 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[87\]_B user_to_mprj_in_gates\[87\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_440 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_934 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_495 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_956 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[121\] _585_/Y la_data_in_core[121] la_buf\[121\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xmprj_adr_buf\[29\] _429_/Y mprj_adr_o_user[29] mprj_adr_buf\[29\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xoutput708 vccd vssd la_data_in_mprj[58] output708/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput719 vccd vssd la_data_in_mprj[68] output719/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_45_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1109 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[72\]_A user_to_mprj_in_gates\[72\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[11\]_B user_to_mprj_in_gates\[11\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_39_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__477__A _477_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1754 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[54\] user_to_mprj_in_gates\[54\]/Y user_to_mprj_in_gates\[54\]/B
+ input81/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_48_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1583 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_226 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[78\]_B user_to_mprj_in_gates\[78\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_17_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1135 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_609 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[110\]_A user_to_mprj_in_gates\[110\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1621 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2219 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[63\]_A user_to_mprj_in_gates\[63\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input9_A la_data_out_core[104] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2090 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__387__A _387_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_329 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[69\]_B user_to_mprj_in_gates\[69\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input273_A la_iena_mprj[111] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2119 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[101\]_A user_to_mprj_in_gates\[101\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1721 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input440_A la_oenb_mprj[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_653 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[54\]_A user_to_mprj_in_gates\[54\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input538_A mprj_adr_o_core[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[101\]_A_N _364_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_189 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_636_ _636_/A _636_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf_enable\[116\]_A_N _379_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_567_ _567_/Y _567_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_mprj_adr_buf\[22\]_TE mprj_adr_buf\[22\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[94\]_A _558_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_498_ _498_/Y _498_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_53_1769 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[24\] user_to_mprj_in_gates\[24\]/Y output671/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_51_1493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output757_A output757/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_491 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[45\]_A user_to_mprj_in_gates\[45\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_833 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1046 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_877 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1956 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[85\]_A _549_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1989 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1028 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[36\]_A user_to_mprj_in_gates\[36\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[64\] vccd vssd user_to_mprj_in_gates\[64\]/B mprj_logic_high_inst/HI[394]
+ input348/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_8_1567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input119_A la_data_out_core[89] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[42\] la_buf\[42\]/TE _634_/A la_buf_enable\[42\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[2\] _594_/Y la_oenb_core[2] mprj_logic_high_inst/HI[204]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[20\] _612_/Y la_oenb_core[20] mprj_logic_high_inst/HI[222]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_421_ _421_/A _421_/Y vssd vccd vssd vccd sky130_fd_sc_hd__inv_12
XFILLER_53_181 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_844 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_352_ _352_/Y _352_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_gates\[126\]_B user_to_mprj_in_gates\[126\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[76\]_A _540_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input390_A la_oenb_mprj[101] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input84_A la_data_out_core[57] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[94\]_B la_buf_enable\[94\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input488_A la_oenb_mprj[75] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_763 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__580__A _580_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[28\] _492_/Y la_data_in_core[28] la_buf\[28\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_13_1731 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_60 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_266 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_93 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[27\]_A user_to_mprj_in_gates\[27\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2149 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1022 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput9 vccd vssd input9/X la_data_out_core[104] vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_la_buf\[16\]_TE la_buf\[16\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_619_ _619_/Y _619_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_17_351 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[67\]_A _531_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[117\]_B user_to_mprj_in_gates\[117\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_32_387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[17\] user_to_mprj_in_gates\[17\]/Y user_to_mprj_in_gates\[17\]/B
+ input40/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_la_buf_enable\[85\]_B la_buf_enable\[85\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_550 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__490__A _490_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[27\] output775/A user_wb_dat_gates\[27\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_25_2347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[18\]_A user_to_mprj_in_gates\[18\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[26\]_A input568/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2110 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1729 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2165 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_181 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[58\]_A _522_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[108\]_B user_to_mprj_in_gates\[108\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_51_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[76\]_B la_buf_enable\[76\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1341 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1959 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_737 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[68\] _331_/Y la_oenb_core[68] mprj_logic_high_inst/HI[270]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_8_1320 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[17\]_A input558/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1768 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[16\] _448_/Y mprj_dat_o_user[16] mprj_dat_buf\[16\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input236_A la_data_out_mprj[79] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[39\]_TE la_buf\[39\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_413 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input403_A la_oenb_mprj[113] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2229 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2218 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__575__A _575_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_82 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[49\]_A _513_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_71 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_60 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_404_ _404_/A _404_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
X_335_ _335_/Y _335_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_41_162 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_93 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_836 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[67\]_B la_buf_enable\[67\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[11\] _411_/Y mprj_adr_o_user[11] mprj_adr_buf\[11\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[125\] user_to_mprj_in_gates\[125\]/Y output655/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_38_903 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[91\] user_to_mprj_in_gates\[91\]/Y output745/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_49_273 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_424 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_939 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__485__A _485_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1784 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[1\] output767/A user_wb_dat_gates\[1\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_user_to_mprj_in_ena_buf\[70\]_B mprj_logic_high_inst/HI[400] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_663 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[7\]_TE la_buf\[7\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2097 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[58\]_B la_buf_enable\[58\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[60\]_A _652_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[125\]_A _388_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput619 vccd vssd _394_/A mprj_stb_o_core vssd vccd sky130_fd_sc_hd__buf_4
Xinput608 vccd vssd _436_/A mprj_dat_o_core[4] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_9_1651 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1504 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_917 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__395__A _395_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[27\] vccd vssd user_to_mprj_in_gates\[27\]/B mprj_logic_high_inst/HI[357]
+ input307/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_ena_buf\[61\]_B mprj_logic_high_inst/HI[391] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_52_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_162 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[49\]_B la_buf_enable\[49\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[51\]_A _643_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[116\]_A _379_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input186_A la_data_out_mprj[33] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input353_A la_iena_mprj[69] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input47_A la_data_out_core[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input520_A mprj_adr_o_core[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[110\] la_buf\[110\]/TE _373_/A la_buf_enable\[110\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf_enable\[74\]_A_N _337_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[95\] _559_/Y la_data_in_core[95] la_buf\[95\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[0\] vccd vssd user_to_mprj_in_gates\[0\]/B mprj_logic_high_inst/HI[330]
+ input260/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_input618_A mprj_sel_o_core[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_777 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[89\]_A_N _352_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1957 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[52\]_B mprj_logic_high_inst/HI[382] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_43_983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[12\]_A_N _604_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput12 input12/X la_data_out_core[107] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput34 input34/X la_data_out_core[127] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput23 input23/X la_data_out_core[117] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput45 input45/X la_data_out_core[21] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_ena_buf\[9\]_A input387/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_891 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput89 vccd vssd input89/X la_data_out_core[61] vssd vccd sky130_fd_sc_hd__buf_4
Xinput78 vccd vssd input78/X la_data_out_core[51] vssd vccd sky130_fd_sc_hd__buf_4
Xinput67 vccd vssd input67/X la_data_out_core[41] vssd vccd sky130_fd_sc_hd__buf_4
Xinput56 input56/X la_data_out_core[31] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_oen_buffers\[107\]_A _370_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[42\]_A _634_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1421 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[27\]_A_N _619_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[84\] user_to_mprj_in_gates\[84\]/Y user_to_mprj_in_gates\[84\]/B
+ input114/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_6_1813 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_232 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1868 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_257 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[43\]_B mprj_logic_high_inst/HI[373] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_21_611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_165 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[33\]_A _625_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1019 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2239 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput427 vccd vssd _593_/A la_oenb_mprj[1] vssd vccd sky130_fd_sc_hd__buf_2
Xinput405 _378_/A la_oenb_mprj[115] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput416 _388_/A la_oenb_mprj[125] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput449 la_oenb_mprj[3] _595_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput438 vccd vssd _594_/A la_oenb_mprj[2] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_5_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input101_A la_data_out_core[72] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[34\]_B mprj_logic_high_inst/HI[364] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_942 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1845 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input470_A la_oenb_mprj[59] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input568_A mprj_dat_i_user[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[112\]_TE mprj_logic_high_inst/HI[314] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[24\]_A _616_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[6\] _470_/Y la_data_in_core[6] la_buf\[6\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_7_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[10\] _474_/Y la_data_in_core[10] la_buf\[10\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_49_1785 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[3\] _403_/Y mprj_adr_o_user[3] mprj_adr_buf\[3\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_47_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_we_buf_TE mprj_we_buf/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[20\]_A _420_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[25\]_B mprj_logic_high_inst/HI[355] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[54\] user_to_mprj_in_gates\[54\]/Y output704/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output787_A output787/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1177 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_953 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_430 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[12\] user_wb_dat_gates\[12\]/Y input553/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_50_2078 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[11\]_TE mprj_logic_high_inst/HI[213] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[15\]_A _607_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1295 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[110\] user_to_mprj_in_gates\[110\]/Y user_to_mprj_in_gates\[110\]/B
+ input16/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_6_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[11\]_A _411_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_585 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1932 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[16\]_B mprj_logic_high_inst/HI[346] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_43_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_268 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[9\]_A input581/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[94\] vccd vssd user_to_mprj_in_gates\[94\]/B mprj_logic_high_inst/HI[424]
+ input381/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_46_1925 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[120\] _383_/Y la_oenb_core[120] mprj_logic_high_inst/HI[322]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_sel_buf\[1\] _397_/Y mprj_sel_o_user[1] mprj_sel_buf\[1\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xinput202 la_data_out_mprj[48] _512_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_40_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[9\]_A input131/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput213 la_data_out_mprj[58] _522_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput224 la_data_out_mprj[68] _532_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput235 vccd vssd _542_/A la_data_out_mprj[78] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_7_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input149_A la_data_out_mprj[115] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[72\] la_buf\[72\]/TE _335_/A la_buf_enable\[72\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_40_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1524 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[50\] _642_/Y la_oenb_core[50] mprj_logic_high_inst/HI[252]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_29_530 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput246 vccd vssd _552_/A la_data_out_mprj[88] vssd vccd sky130_fd_sc_hd__buf_2
Xinput257 vccd vssd _562_/A la_data_out_mprj[98] vssd vccd sky130_fd_sc_hd__buf_2
Xinput268 vssd vccd input268/X la_iena_mprj[107] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput279 vssd vccd input279/X la_iena_mprj[117] vssd vccd sky130_fd_sc_hd__clkbuf_1
X_652_ _652_/A _652_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_input316_A la_iena_mprj[35] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_583_ _583_/A _583_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
Xla_buf\[58\] _522_/Y la_data_in_core[58] la_buf\[58\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__583__A _583_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_249 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1620 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[34\]_TE mprj_logic_high_inst/HI[236] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_946 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput709 vccd vssd la_data_in_mprj[59] output709/A vssd vccd sky130_fd_sc_hd__buf_2
Xla_buf\[114\] _578_/Y la_data_in_core[114] la_buf\[114\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_45_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1711 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output702_A output702/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1766 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1985 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1799 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[47\] user_to_mprj_in_gates\[47\]/Y user_to_mprj_in_gates\[47\]/B
+ input73/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_50_525 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__493__A _493_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_238 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[9\]_TE mprj_adr_buf\[9\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1141 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1147 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[9\] user_to_mprj_in_gates\[9\]/Y input131/X user_to_mprj_in_gates\[9\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_1_109 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1727 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[72\]_TE la_buf\[72\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[57\]_TE mprj_logic_high_inst/HI[259] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_739 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1648 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[98\] _361_/Y la_oenb_core[98] mprj_logic_high_inst/HI[300]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input266_A la_iena_mprj[105] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_632 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input433_A la_oenb_mprj[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__578__A _578_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input600_A mprj_dat_o_core[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_831 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1365 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_635_ _635_/Y _635_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_mprj_dat_buf\[24\]_A _456_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[31\]_A user_wb_dat_gates\[31\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_45_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_566_ _566_/A _566_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_mprj_dat_buf\[21\]_TE mprj_dat_buf\[21\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1737 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1261 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_497_ _497_/Y _497_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_oen_buffers\[0\]_TE mprj_logic_high_inst/HI[202] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_8_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[17\] user_to_mprj_in_gates\[17\]/Y output663/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_47_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output652_A output652/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[95\]_TE la_buf\[95\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__488__A _488_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2314 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[15\]_A _447_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[22\]_A user_wb_dat_gates\[22\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_50_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1058 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_385 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2213 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1589 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1917 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__398__A _398_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1485 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[57\] vccd vssd user_to_mprj_in_gates\[57\]/B mprj_logic_high_inst/HI[387]
+ input340/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_2_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[13\]_A user_wb_dat_gates\[13\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_2_1178 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_420_ _420_/Y _420_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkinv_8
XFILLER_14_503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[13\] _605_/Y la_oenb_core[13] mprj_logic_high_inst/HI[215]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_351_ _351_/A _351_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
Xla_buf_enable\[35\] la_buf\[35\]/TE _627_/A la_buf_enable\[35\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_39_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[9\] output754/A user_to_mprj_in_gates\[9\]/Y vccd vssd vssd
+ vccd sky130_fd_sc_hd__inv_6
XANTENNA_input383_A la_iena_mprj[96] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1743 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_713 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_775 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input77_A la_data_out_core[50] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input550_A mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_72 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_985 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1089 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_618_ _618_/A _618_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_300 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_549_ _549_/Y _549_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_9_562 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2326 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1811 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_29 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1855 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[26\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_617 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_609 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[100\]_A_N _363_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_215 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[12\]_TE mprj_adr_buf\[12\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1861 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[115\]_A_N _378_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[17\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input131_A la_data_out_core[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_926 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input229_A la_data_out_mprj[72] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_469 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_403_ _403_/A _403_/Y vssd vccd vssd vccd sky130_fd_sc_hd__inv_12
XANTENNA_la_buf\[2\]_A _466_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_83 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_804 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_50 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_72 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_61 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input598_A mprj_dat_o_core[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[40\] _504_/Y la_data_in_core[40] la_buf\[40\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_334_ _334_/Y _334_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_30_848 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_94 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__591__A _591_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[112\] vccd vssd user_to_mprj_in_gates\[112\]/B mprj_logic_high_inst/HI[442]
+ input274/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_31_1117 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[118\] user_to_mprj_in_gates\[118\]/Y output647/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_irq_gates\[2\]_A input623/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_915 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_281 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1257 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[84\] user_to_mprj_in_gates\[84\]/Y output737/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_37_436 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[0\]_TE mprj_dat_buf\[0\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_981 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1796 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_152 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[120\]_TE la_buf\[120\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1673 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1102 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput609 _437_/A mprj_dat_o_core[5] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1251 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[9\]_A _409_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_973 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_303 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[80\] _343_/Y la_oenb_core[80] mprj_logic_high_inst/HI[282]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input179_A la_data_out_mprj[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1978 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[50\]_A input77/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input346_A la_iena_mprj[62] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2289 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input513_A la_oenb_mprj[98] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[88\] _552_/Y la_data_in_core[88] la_buf\[88\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__586__A _586_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1048 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[103\] la_buf\[103\]/TE _366_/A la_buf_enable\[103\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_46_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2205 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1771 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1602 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[0\]_A user_to_mprj_in_gates\[0\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2249 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xinput13 vccd vssd input13/X la_data_out_core[108] vssd vccd sky130_fd_sc_hd__buf_4
Xinput24 input24/X la_data_out_core[118] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput46 vccd vssd input46/X la_data_out_core[22] vssd vccd sky130_fd_sc_hd__buf_4
Xinput35 la_data_out_core[12] input35/X vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_ena_buf\[9\]_B mprj_logic_high_inst/HI[339] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_7_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput79 vccd vssd input79/X la_data_out_core[52] vssd vccd sky130_fd_sc_hd__buf_4
Xinput68 input68/X la_data_out_core[42] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput57 vccd vssd input57/X la_data_out_core[32] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_48_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_391 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output732_A output732/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[41\]_A input67/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1308 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[77\] user_to_mprj_in_gates\[77\]/Y user_to_mprj_in_gates\[77\]/B
+ input106/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_38_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__496__A _496_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2261 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_266 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_491 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_973 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[90\]_TE mprj_logic_high_inst/HI[292] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1172 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[29\]_TE la_buf\[29\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[32\]_A input57/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput428 la_oenb_mprj[20] _612_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput406 _379_/A la_oenb_mprj[116] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput417 _389_/A la_oenb_mprj[126] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput439 vccd vssd _622_/A la_oenb_mprj[30] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_5_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2314 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_277 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[99\]_A input130/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1613 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_954 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_627 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input296_A la_iena_mprj[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_667 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_137 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input463_A la_oenb_mprj[52] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_844 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[23\]_A input47/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_365 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_553 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_781 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_921 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_932 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1719 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[47\] user_to_mprj_in_gates\[47\]/Y output696/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_output682_A output682/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_987 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_442 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[14\]_A input37/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1127 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[103\] user_to_mprj_in_gates\[103\]/Y user_to_mprj_in_gates\[103\]/B
+ input8/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_39_1922 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1944 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[9\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[73\]_A_N _336_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[88\]_A_N _351_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[87\] vccd vssd user_to_mprj_in_gates\[87\]/B mprj_logic_high_inst/HI[417]
+ input373/X vssd vccd sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[113\] _376_/Y la_oenb_core[113] mprj_logic_high_inst/HI[315]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xmprj_clk2_buf _392_/Y user_clock2 mprj_clk2_buf/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xinput203 la_data_out_mprj[49] _513_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_gates\[9\]_B user_to_mprj_in_gates\[9\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput214 la_data_out_mprj[59] _523_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput225 la_data_out_mprj[69] _533_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput236 _543_/A la_data_out_mprj[79] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[11\]_A_N _603_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput247 vccd vssd la_data_out_mprj[89] _553_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput258 la_data_out_mprj[99] _563_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput269 vssd vccd input269/X la_iena_mprj[108] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xuser_to_mprj_oen_buffers\[43\] _635_/Y la_oenb_core[43] mprj_logic_high_inst/HI[245]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[65\] la_buf\[65\]/TE _657_/A la_buf_enable\[65\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_40_1536 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_651_ _651_/A _651_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_5_1165 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_irq_buffers\[1\] user_irq_gates\[1\]/Y output793/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_44_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_582_ _582_/A _582_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_input211_A la_data_out_mprj[56] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[26\]_A_N _618_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input309_A la_iena_mprj[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2322 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input580_A mprj_dat_i_user[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1627 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2273 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1561 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[107\] _571_/Y la_data_in_core[107] la_buf\[107\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_45_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[100\] user_to_mprj_in_gates\[100\]/Y output628/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_3_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_545 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[120\]_A input283/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1197 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_991 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1981 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2028 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[102\]_TE mprj_logic_high_inst/HI[304] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_523 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1485 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_545 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[111\]_A input273/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2339 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1785 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_924 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1701 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input259_A la_data_out_mprj[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input161_A la_data_out_mprj[126] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input426_A la_oenb_mprj[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input22_A la_data_out_core[116] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2089 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
X_634_ _634_/A _634_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
Xla_buf\[70\] _534_/Y la_data_in_core[70] la_buf\[70\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_45_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__594__A _594_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_565_ _565_/Y _565_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_53_1705 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_496_ _496_/Y _496_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_18_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[102\]_A input263/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_581 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_755 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_788 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output645_A output645/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[125\]_TE mprj_logic_high_inst/HI[327] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1761 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2326 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1625 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_301 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1925 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1453 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[24\]_TE mprj_logic_high_inst/HI[226] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[91\]_A input378/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_802 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
X_350_ _350_/A _350_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_14_515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[28\] la_buf\[28\]/TE _620_/A la_buf_enable\[28\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_13_1755 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_747 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input376_A la_iena_mprj[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1206 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input543_A mprj_adr_o_core[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1553 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__589__A _589_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_975 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1715 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1737 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[82\]_A input368/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_109 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_617_ _617_/Y _617_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_53_2203 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_548_ _548_/Y _548_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_17_375 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_479_ _479_/A _479_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_53_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output762_A output762/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_574 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[62\]_TE la_buf\[62\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[47\]_TE mprj_logic_high_inst/HI[249] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__499__A _499_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1867 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[73\]_A input358/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_161 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_665 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1733 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_378 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[9\]_B la_buf_enable\[9\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[11\]_TE mprj_dat_buf\[11\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1261 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_938 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input124_A la_data_out_core[93] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[64\]_A input348/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_402_ _402_/A _402_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XPHY_40 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_62 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_51 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_73 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_333_ _333_/Y _333_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XPHY_95 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_84 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input493_A la_oenb_mprj[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[85\]_TE la_buf\[85\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[33\] _497_/Y la_data_in_core[33] la_buf\[33\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_6_511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[105\] vccd vssd user_to_mprj_in_gates\[105\]/B mprj_logic_high_inst/HI[435]
+ input266/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_10_551 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[5\] user_wb_dat_gates\[5\]/Y input577/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_48_2305 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_gates\[2\]_B user_irq_gates\[2\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_33 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[55\]_A input338/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[77\] user_to_mprj_in_gates\[77\]/Y output729/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_46_971 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_109 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1029 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[22\] user_to_mprj_in_gates\[22\]/Y user_to_mprj_in_gates\[22\]/B
+ input46/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_33_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_197 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1114 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1642 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2179 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[3\]_A _399_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_949 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[46\]_A input328/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_440 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_359 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1449 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[50\]_B user_to_mprj_in_gates\[50\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[73\] _336_/Y la_oenb_core[73] mprj_logic_high_inst/HI[275]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[95\] la_buf\[95\]/TE _358_/A la_buf_enable\[95\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xoutput690 vccd vssd la_data_in_mprj[41] output690/A vssd vccd sky130_fd_sc_hd__buf_2
Xmprj_dat_buf\[21\] _453_/Y mprj_dat_o_user[21] mprj_dat_buf\[21\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input339_A la_iena_mprj[56] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input241_A la_data_out_mprj[83] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1005 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_245 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[37\]_A input318/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input506_A la_oenb_mprj[91] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_61 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[4\]_A _436_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput25 input25/X la_data_out_core[119] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput14 input14/X la_data_out_core[109] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput36 vccd vssd input36/X la_data_out_core[13] vssd vccd sky130_fd_sc_hd__buf_4
Xinput69 input69/X la_data_out_core[43] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput58 input58/X la_data_out_core[33] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput47 vccd vssd input47/X la_data_out_core[23] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_48_2113 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2146 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[41\]_B user_to_mprj_in_gates\[41\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1456 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output725_A output725/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1033 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_256 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[28\]_A input308/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_429 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[114\]_A_N _377_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[1\] la_buf\[1\]/TE _593_/A la_buf_enable\[1\]/B vssd vccd vssd vccd
+ sky130_fd_sc_hd__and2b_1
XFILLER_31_1493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[32\]_B user_to_mprj_in_gates\[32\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[93\]_A user_to_mprj_in_gates\[93\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput407 _380_/A la_oenb_mprj[117] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput418 _390_/A la_oenb_mprj[127] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput429 vccd vssd _613_/A la_oenb_mprj[21] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_5_2059 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[19\]_A input298/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_749 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[32\] vccd vssd user_to_mprj_in_gates\[32\]/B mprj_logic_high_inst/HI[362]
+ input313/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_43_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[99\]_B user_to_mprj_in_gates\[99\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_52_793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_966 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_105 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[10\] la_buf\[10\]/TE _602_/A la_buf_enable\[10\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_22_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input191_A la_data_out_mprj[38] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input289_A la_iena_mprj[126] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[120\]_A _584_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input456_A la_oenb_mprj[46] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[84\]_A user_to_mprj_in_gates\[84\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[23\]_B user_to_mprj_in_gates\[23\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input52_A la_data_out_core[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input623_A user_irq_core[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[110\]_TE la_buf\[110\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__597__A _597_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[25\]_TE mprj_adr_buf\[25\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1712 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1113 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_944 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output675_A output675/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_999 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[122\]_A user_to_mprj_in_gates\[122\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[111\]_A _575_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[14\]_B user_to_mprj_in_gates\[14\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[75\]_A user_to_mprj_in_gates\[75\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1117 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1139 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_215 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1956 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2289 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[113\]_A user_to_mprj_in_gates\[113\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1599 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[102\]_A _566_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[66\]_A user_to_mprj_in_gates\[66\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_837 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput226 la_data_out_mprj[6] _470_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput215 la_data_out_mprj[5] _469_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput204 la_data_out_mprj[4] _468_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_40_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[106\] _369_/Y la_oenb_core[106] mprj_logic_high_inst/HI[308]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xinput259 la_data_out_mprj[9] _473_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput248 vccd vssd la_data_out_mprj[8] _472_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput237 la_data_out_mprj[7] _471_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
X_650_ _650_/Y _650_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
X_581_ _581_/Y _581_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[58\] la_buf\[58\]/TE _650_/A la_buf_enable\[58\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_44_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[36\] _628_/Y la_oenb_core[36] mprj_logic_high_inst/HI[238]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_29_576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_557 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input204_A la_data_out_mprj[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2334 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1477 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_403 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input573_A mprj_dat_i_user[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[104\]_A user_to_mprj_in_gates\[104\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2105 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[57\]_A user_to_mprj_in_gates\[57\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[30\]_A _494_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[80\]_TE mprj_logic_high_inst/HI[282] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[19\]_TE la_buf\[19\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[97\]_A _561_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output792_A output792/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[120\]_B mprj_logic_high_inst/HI[450] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_31_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1853 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_785 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[48\]_A user_to_mprj_in_gates\[48\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1061 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[21\]_A _485_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1317 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[88\]_A _552_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[111\]_B mprj_logic_high_inst/HI[441] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_947 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1959 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[39\]_A user_to_mprj_in_gates\[39\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[12\]_A _476_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input154_A la_data_out_mprj[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[30\]_B la_buf_enable\[30\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2057 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input321_A la_iena_mprj[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input15_A la_data_out_core[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_633_ _633_/A _633_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_input419_A la_oenb_mprj[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[79\]_A _543_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_888 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_877 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_564_ _564_/A _564_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
Xla_buf\[63\] _527_/Y la_data_in_core[63] la_buf\[63\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_2_1884 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_538 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_495_ _495_/Y _495_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_ena_buf\[102\]_B mprj_logic_high_inst/HI[432] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2120 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_590 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[97\]_B la_buf_enable\[97\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_767 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[27\] _427_/Y mprj_adr_o_user[27] mprj_adr_buf\[27\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_output638_A output638/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_ack_gate user_wb_ack_gate/Y input516/X user_wb_ack_gate/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_49_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[21\]_B la_buf_enable\[21\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2338 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[72\]_A_N _335_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1565 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[52\] user_to_mprj_in_gates\[52\]/Y user_to_mprj_in_gates\[52\]/B
+ input79/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
Xinput590 mprj_dat_o_core[17] _449_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_47_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[87\]_A_N _350_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_2004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1205 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_357 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[88\]_B la_buf_enable\[88\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2204 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[10\]_A_N _602_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[90\]_A _353_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[25\]_A_N _617_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[29\]_A input571/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2019 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input7_A la_data_out_core[102] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[12\]_B la_buf_enable\[12\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1559 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1621 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1272 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[91\]_B mprj_logic_high_inst/HI[421] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_26_365 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_825 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_398 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[79\]_B la_buf_enable\[79\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_700 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[81\]_A _344_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1767 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_225 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input271_A la_iena_mprj[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input369_A la_iena_mprj[83] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_85 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input536_A mprj_adr_o_core[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_486 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[126\] la_buf\[126\]/TE _389_/A la_buf_enable\[126\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_4_1913 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1979 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[82\]_B mprj_logic_high_inst/HI[412] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_45_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_616_ _616_/Y _616_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_40_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_547_ _547_/Y _547_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_17_387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_478_ _478_/A _478_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_9_531 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[72\]_A _335_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[22\] user_to_mprj_in_gates\[22\]/Y output669/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_51_1271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output755_A output755/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_781 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1785 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2293 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1445 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[73\]_B mprj_logic_high_inst/HI[403] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_50_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[63\]_A _655_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2045 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_729 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1841 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1727 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[62\] vccd vssd user_to_mprj_in_gates\[62\]/B mprj_logic_high_inst/HI[392]
+ input346/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_41_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[64\]_B mprj_logic_high_inst/HI[394] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input117_A la_data_out_core[87] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[40\] la_buf\[40\]/TE _632_/A la_buf_enable\[40\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[0\] _592_/Y la_oenb_core[0] mprj_logic_high_inst/HI[202]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_27_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_401_ _401_/A _401_/Y vssd vccd vssd vccd sky130_fd_sc_hd__inv_12
XPHY_30 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_74 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_63 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_52 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_41 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_332_ _332_/A _332_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XPHY_96 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_85 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1233 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input82_A la_data_out_core[55] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[115\]_TE mprj_logic_high_inst/HI[317] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[119\]_A _382_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[54\]_A _646_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_390 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input486_A la_oenb_mprj[73] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[26\] _490_/Y la_data_in_core[26] la_buf\[26\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_13_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_523 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2052 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1958 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_795 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_89 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[55\]_B mprj_logic_high_inst/HI[385] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2045 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_305 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_wb_dat_gates\[28\] user_wb_dat_gates\[28\]/Y input570/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_33_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[15\] user_to_mprj_in_gates\[15\]/Y input38/X user_to_mprj_in_gates\[15\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_53_1377 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[45\]_A _637_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[14\]_TE mprj_logic_high_inst/HI[216] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_372 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[25\] output773/A user_wb_dat_gates\[25\]/Y vccd vssd vssd vccd
+ sky130_fd_sc_hd__inv_6
XFILLER_29_2250 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[126\] user_to_mprj_in_gates\[126\]/Y user_to_mprj_in_gates\[126\]/B
+ input33/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_9_1687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[46\]_B mprj_logic_high_inst/HI[376] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[36\]_A _628_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1851 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1704 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput680 vccd vssd la_data_in_mprj[32] output680/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_43_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[66\] _329_/Y la_oenb_core[66] mprj_logic_high_inst/HI[268]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[88\] la_buf\[88\]/TE _351_/A la_buf_enable\[88\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xoutput691 vccd vssd la_data_in_mprj[42] output691/A vssd vccd sky130_fd_sc_hd__buf_2
Xmprj_dat_buf\[14\] _446_/Y mprj_dat_o_user[14] mprj_dat_buf\[14\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_19_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input234_A la_data_out_mprj[77] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1164 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1175 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1811 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1281 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1855 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[37\]_B mprj_logic_high_inst/HI[367] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_19_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1916 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[52\]_TE la_buf\[52\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input401_A la_oenb_mprj[111] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_600 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_633 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[37\]_TE mprj_logic_high_inst/HI[239] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1751 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_61 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput37 vccd vssd input37/X la_data_out_core[14] vssd vccd sky130_fd_sc_hd__buf_4
Xinput26 la_data_out_core[11] input26/X vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput15 input15/X la_data_out_core[10] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_oen_buffers\[27\]_A _619_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput59 input59/X la_data_out_core[34] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput48 vccd vssd input48/X la_data_out_core[24] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_48_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1468 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[123\] user_to_mprj_in_gates\[123\]/Y output653/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_46_1181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output718_A output718/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[23\]_A _423_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2191 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[28\]_B mprj_logic_high_inst/HI[358] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_34_920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_249 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1704 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[18\]_A _610_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[0\]_A _592_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2151 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2195 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput419 vccd vssd _604_/A la_oenb_mprj[12] vssd vccd sky130_fd_sc_hd__buf_2
Xinput408 _381_/A la_oenb_mprj[118] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1451 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1877 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[75\]_TE la_buf\[75\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1337 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[14\]_A _414_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[19\]_B mprj_logic_high_inst/HI[349] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_43_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[25\] vccd vssd user_to_mprj_in_gates\[25\]/B mprj_logic_high_inst/HI[355]
+ input305/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_24_441 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1902 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input184_A la_data_out_mprj[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input449_A la_oenb_mprj[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input351_A la_iena_mprj[67] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input45_A la_data_out_core[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[93\] _557_/Y la_data_in_core[93] la_buf\[93\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input616_A mprj_sel_o_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[24\]_TE mprj_dat_buf\[24\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[3\]_TE mprj_logic_high_inst/HI[205] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_30_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_466 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output668_A output668/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1817 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[98\]_TE la_buf\[98\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2242 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_890 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[82\] user_to_mprj_in_gates\[82\]/Y user_to_mprj_in_gates\[82\]/B
+ input112/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_26_2275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_205 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2093 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_547 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2257 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1843 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput205 la_data_out_mprj[50] _514_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput216 la_data_out_mprj[60] _524_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput227 vccd vssd _534_/A la_data_out_mprj[70] vssd vccd sky130_fd_sc_hd__buf_2
Xinput238 _544_/A la_data_out_mprj[80] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput249 vssd vccd _554_/A la_data_out_mprj[90] vssd vccd sky130_fd_sc_hd__clkbuf_1
X_580_ _580_/A _580_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_29_588 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_525 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[29\] _621_/Y la_oenb_core[29] mprj_logic_high_inst/HI[231]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_31_208 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2346 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1309 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_293 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_63 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_426 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input399_A la_oenb_mprj[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_96 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input566_A mprj_dat_i_user[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[4\] _468_/Y la_data_in_core[4] la_buf\[4\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_49_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1449 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[113\]_A_N _376_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__401__A _401_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1883 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[1\] _401_/Y mprj_adr_o_user[1] mprj_adr_buf\[1\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_7_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[27\]_A _459_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_385 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1521 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[52\] user_to_mprj_in_gates\[52\]/Y output702/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_output785_A output785/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[10\] user_wb_dat_gates\[10\]/Y input551/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_28_2304 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[18\]_A _450_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[25\]_A user_wb_dat_gates\[25\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_41_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[100\]_TE la_buf\[100\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[15\]_TE mprj_adr_buf\[15\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1651 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[92\] vccd vssd user_to_mprj_in_gates\[92\]/B mprj_logic_high_inst/HI[422]
+ input379/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_0_145 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_639 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2025 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1229 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input147_A la_data_out_mprj[113] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[70\] la_buf\[70\]/TE _333_/A la_buf_enable\[70\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_28_41 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_632_ _632_/Y _632_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_29_341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[16\]_A user_wb_dat_gates\[16\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_28_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input314_A la_iena_mprj[33] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_563_ _563_/Y _563_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf\[56\] _520_/Y la_data_in_core[56] la_buf\[56\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_494_ _494_/Y _494_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_38_1253 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2154 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_wb_ena_buf user_wb_ack_gate/B user_to_mprj_wb_ena_buf/B input614/X vssd
+ vccd vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_9_735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1453 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_779 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1901 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[112\] _576_/Y la_data_in_core[112] la_buf\[112\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_49_1393 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[3\]_TE mprj_dat_buf\[3\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output700_A output700/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput580 mprj_dat_i_user[8] input580/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
Xinput591 mprj_dat_o_core[18] _450_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_la_buf_enable\[120\]_B la_buf_enable\[120\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[45\] user_to_mprj_in_gates\[45\]/Y input71/X user_to_mprj_in_gates\[45\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_23_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[123\]_TE la_buf\[123\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[7\] user_to_mprj_in_gates\[7\]/Y input109/X user_to_mprj_in_gates\[7\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_4
XANTENNA_user_wb_dat_gates\[29\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2345 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1677 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_303 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[111\]_B la_buf_enable\[111\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[70\]_TE mprj_logic_high_inst/HI[272] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_712 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[2\]_A user_wb_dat_gates\[2\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[96\] _359_/Y la_oenb_core[96] mprj_logic_high_inst/HI[298]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[80\]_A input110/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input264_A la_iena_mprj[103] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1533 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_443 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input431_A la_oenb_mprj[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1588 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[9\] vccd vssd user_to_mprj_in_gates\[9\]/B mprj_logic_high_inst/HI[339]
+ input387/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_7_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input529_A mprj_adr_o_core[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[119\] vccd vssd la_buf\[119\]/TE la_buf_enable\[119\]/B _382_/A vssd
+ vccd sky130_fd_sc_hd__and2b_2
XFILLER_40_1132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_95 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_609 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1728 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1969 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[5\]_A _469_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_615_ _615_/A _615_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_546_ _546_/Y _546_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf_enable\[102\]_B la_buf_enable\[102\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_477_ _477_/Y _477_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_358 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_881 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1283 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[15\] user_to_mprj_in_gates\[15\]/Y output661/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output748_A output748/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output650_A output650/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[71\]_A input100/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1457 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[93\]_TE mprj_logic_high_inst/HI[295] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_133 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_881 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[62\]_A input90/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj2_pwrgood mprj2_pwrgood/A output790/A vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
XFILLER_8_1335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[55\] vccd vssd user_to_mprj_in_gates\[55\]/B mprj_logic_high_inst/HI[385]
+ input338/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_41_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_697 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_400_ _400_/Y _400_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XPHY_31 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_20 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[11\] _603_/Y la_oenb_core[11] mprj_logic_high_inst/HI[213]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_331_ _331_/A _331_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XPHY_64 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_53 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_42 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_97 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_86 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[33\] la_buf\[33\]/TE _625_/A la_buf_enable\[33\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XPHY_75 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[7\] user_to_mprj_in_gates\[7\]/Y output732/A vccd vssd vssd
+ vccd sky130_fd_sc_hd__clkinv_4
XFILLER_19_1999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1109 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input381_A la_iena_mprj[94] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[71\]_A_N _334_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input479_A la_oenb_mprj[67] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input75_A la_data_out_core[49] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[19\] _483_/Y la_data_in_core[19] la_buf\[19\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_13_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[53\]_A input80/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1005 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2064 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[86\]_A_N _349_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1915 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1205 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1249 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_409 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1569 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[24\]_A_N _616_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[3\]_A user_to_mprj_in_gates\[3\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_output698_A output698/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_529_ _529_/Y _529_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_133 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1345 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1621 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_395 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[39\]_A_N _631_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[44\]_A input70/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2262 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2104 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_buffers\[18\] output765/A user_wb_dat_gates\[18\]/Y vccd vssd vssd vccd
+ sky130_fd_sc_hd__inv_6
XFILLER_29_1561 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_vdd_pwrgood_A mprj_vdd_pwrgood/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1699 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_417 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[119\] user_to_mprj_in_gates\[119\]/Y user_to_mprj_in_gates\[119\]/B
+ input25/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_52_921 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_634 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[35\]_A input60/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1716 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput670 vccd vssd la_data_in_mprj[23] output670/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput681 vccd vssd la_data_in_mprj[33] output681/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2237 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput692 vccd vssd la_data_in_mprj[43] output692/A vssd vccd sky130_fd_sc_hd__buf_2
Xuser_to_mprj_oen_buffers\[59\] _651_/Y la_oenb_core[59] mprj_logic_high_inst/HI[261]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_417 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input227_A la_data_out_mprj[70] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1867 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_965 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1763 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input596_A mprj_dat_o_core[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1053 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[110\] vccd vssd user_to_mprj_in_gates\[110\]/B mprj_logic_high_inst/HI[440]
+ input272/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_11_851 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput27 input27/X la_data_out_core[120] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput16 input16/X la_data_out_core[110] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_7_833 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput49 vccd vssd input49/X la_data_out_core[25] vssd vccd sky130_fd_sc_hd__buf_4
Xinput38 vccd vssd input38/X la_data_out_core[15] vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_user_to_mprj_in_gates\[26\]_A input50/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[110\]_A input16/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__404__A _404_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[116\] user_to_mprj_in_gates\[116\]/Y output645/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_46_1193 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[82\] user_to_mprj_in_gates\[82\]/Y output735/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_4_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_rstn_buf_A input3/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_497 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[17\]_A input40/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_A input6/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1981 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput409 _382_/A la_oenb_mprj[119] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[105\]_TE mprj_logic_high_inst/HI[307] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_217 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2063 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_464 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[18\] vccd vssd user_to_mprj_in_gates\[18\]/B mprj_logic_high_inst/HI[348]
+ input297/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_51_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1373 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_659 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input177_A la_data_out_mprj[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_379 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input344_A la_iena_mprj[60] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input38_A la_data_out_core[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input511_A la_oenb_mprj[96] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[86\] _550_/Y la_data_in_core[86] la_buf\[86\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_21_1631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input609_A mprj_dat_o_core[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[101\] la_buf\[101\]/TE _364_/A la_buf_enable\[101\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_35_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_258 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_486 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_641 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output730_A output730/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[75\] user_to_mprj_in_gates\[75\]/Y user_to_mprj_in_gates\[75\]/B
+ input104/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_6_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1914 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[123\]_A input286/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1991 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[42\]_TE la_buf\[42\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1281 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1899 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2321 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[27\]_TE mprj_logic_high_inst/HI[229] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_828 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput206 la_data_out_mprj[51] _515_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput217 la_data_out_mprj[61] _525_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_48_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput228 la_data_out_mprj[71] _535_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput239 _545_/A la_data_out_mprj[81] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1984 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[114\]_A input276/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_581 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_438 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input294_A la_iena_mprj[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2221 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2265 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input559_A mprj_dat_i_user[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input461_A la_oenb_mprj[50] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2287 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_irq_ena_buf\[1\] vccd vssd user_irq_gates\[1\]/B user_irq_ena_buf\[1\]/B input625/X
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_3_165 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1901 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_865 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2223 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1544 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[105\]_A input266/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_721 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_209 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[45\] user_to_mprj_in_gates\[45\]/Y output694/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output680_A output680/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output778_A output778/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[65\]_TE la_buf\[65\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_798 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1107 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2349 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2051 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1973 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1477 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[101\] user_to_mprj_in_gates\[101\]/Y user_to_mprj_in_gates\[101\]/B
+ input6/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_41_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1733 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1939 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[14\]_TE mprj_dat_buf\[14\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__502__A _502_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[85\] vccd vssd user_to_mprj_in_gates\[85\]/B mprj_logic_high_inst/HI[415]
+ input371/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_44_2151 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[111\] _374_/Y la_oenb_core[111] mprj_logic_high_inst/HI[313]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[94\]_A input381/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[41\] _633_/Y la_oenb_core[41] mprj_logic_high_inst/HI[243]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[63\] la_buf\[63\]/TE _655_/A la_buf_enable\[63\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_29_353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_631_ _631_/A _631_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_44_301 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_562_ _562_/Y _562_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_44_334 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input307_A la_iena_mprj[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_493_ _493_/Y _493_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_44_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[88\]_TE la_buf\[88\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[49\] _513_/Y la_data_in_core[49] la_buf\[49\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_12_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2177 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_747 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__412__A _412_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[105\] _569_/Y la_data_in_core[105] la_buf\[105\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_45_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[85\]_A input371/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput570 mprj_dat_i_user[28] input570/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
Xinput581 mprj_dat_i_user[9] input581/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_36_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_161 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xinput592 mprj_dat_o_core[19] _451_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_1_1341 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_529 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[38\] user_to_mprj_in_gates\[38\]/Y user_to_mprj_in_gates\[38\]/B
+ input63/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_30_1527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[76\]_A input361/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_109 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1116 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1149 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1741 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_893 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[112\]_A_N _375_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[127\]_A_N _390_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[80\]_B user_to_mprj_in_gates\[80\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[89\] _352_/Y la_oenb_core[89] mprj_logic_high_inst/HI[291]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_1_411 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input257_A la_data_out_mprj[98] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1005 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1049 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input20_A la_data_out_core[114] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1854 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input424_A la_oenb_mprj[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[67\]_A input351/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1144 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_614_ _614_/A _614_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_665 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_545_ _545_/Y _545_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_2_1672 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1073 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_476_ _476_/Y _476_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_18_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__407__A _407_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_893 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1961 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[71\]_B user_to_mprj_in_gates\[71\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_5_761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output643_A output643/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[58\]_A input341/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_109 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_189 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1059 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1313 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[62\]_B user_to_mprj_in_gates\[62\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2121 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[49\]_A input331/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1453 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[48\] vccd vssd user_to_mprj_in_gates\[48\]/B mprj_logic_high_inst/HI[378]
+ input330/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_6_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_665 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_21 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_10 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_330_ _330_/Y _330_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XPHY_54 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_65 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_43 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_32 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_98 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_87 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_76 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2261 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1393 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1967 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[26\] la_buf\[26\]/TE _618_/A la_buf_enable\[26\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_6_569 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input374_A la_iena_mprj[88] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[53\]_B user_to_mprj_in_gates\[53\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input68_A la_data_out_core[42] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input541_A mprj_adr_o_core[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2076 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[113\]_TE la_buf\[113\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_764 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_775 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[28\]_TE mprj_adr_buf\[28\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1701 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1745 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1313 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1302 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_528_ _528_/Y _528_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_mprj_dat_buf\[7\]_A _439_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2058 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_459_ _459_/Y _459_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_6
XANTENNA_output760_A output760/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_363 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[44\]_B user_to_mprj_in_gates\[44\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2274 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__600__A _600_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[60\]_TE mprj_logic_high_inst/HI[262] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1233 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_613 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_454 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1533 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[35\]_B user_to_mprj_in_gates\[35\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[96\]_A user_to_mprj_in_gates\[96\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1728 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput660 vccd vssd la_data_in_mprj[14] output660/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput671 vccd vssd la_data_in_mprj[24] output671/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__510__A _510_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput693 vccd vssd la_data_in_mprj[44] output693/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput682 vccd vssd la_data_in_mprj[34] output682/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_43_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1982 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input122_A la_data_out_core[91] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1824 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_53 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[20\]_A user_to_mprj_in_gates\[20\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1879 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_624 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1731 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_668 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input491_A la_oenb_mprj[78] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input589_A mprj_dat_o_core[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput28 input28/X la_data_out_core[121] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput17 input17/X la_data_out_core[111] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_la_buf\[123\]_A _587_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1087 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[31\] _495_/Y la_data_in_core[31] la_buf\[31\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_32_1920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[103\] vccd vssd user_to_mprj_in_gates\[103\]/B mprj_logic_high_inst/HI[433]
+ input264/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_11_863 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_wb_dat_gates\[3\] user_wb_dat_gates\[3\]/Y input575/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
Xinput39 input39/X la_data_out_core[16] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_gates\[26\]_B user_to_mprj_in_gates\[26\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_6_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[87\]_A user_to_mprj_in_gates\[87\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[110\]_B user_to_mprj_in_gates\[110\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_6_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_878 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[60\]_A _524_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[83\]_TE mprj_logic_high_inst/HI[285] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__420__A _420_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[109\] user_to_mprj_in_gates\[109\]/Y output637/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_38_749 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[75\] user_to_mprj_in_gates\[75\]/Y output727/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_4_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[11\]_A user_to_mprj_in_gates\[11\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1597 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1820 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[20\] user_to_mprj_in_gates\[20\]/Y user_to_mprj_in_gates\[20\]/B
+ input44/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_53_1143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1897 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[125\]_A user_to_mprj_in_gates\[125\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[114\]_A _578_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2175 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[17\]_B user_to_mprj_in_gates\[17\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[30\] output779/A user_wb_dat_gates\[30\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_user_to_mprj_in_gates\[101\]_B user_to_mprj_in_gates\[101\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[78\]_A user_to_mprj_in_gates\[78\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[51\]_A _515_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1813 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__330__A _330_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[8\] _440_/Y mprj_dat_o_user[8] mprj_dat_buf\[8\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1475 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[70\]_A_N _333_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2020 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[10\]_A input551/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_273 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[85\]_A_N _348_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_925 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1817 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[116\]_A user_to_mprj_in_gates\[116\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1828 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[105\]_A _569_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__505__A _505_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_693 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_77 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[69\]_A user_to_mprj_in_gates\[69\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1503 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[42\]_A _506_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_859 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[60\]_B la_buf_enable\[60\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[71\] _334_/Y la_oenb_core[71] mprj_logic_high_inst/HI[273]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[23\]_A_N _615_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[93\] la_buf\[93\]/TE _356_/A la_buf_enable\[93\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_43_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input337_A la_iena_mprj[54] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[38\]_A_N _630_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[79\] _543_/Y la_data_in_core[79] la_buf\[79\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_21_1643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input504_A la_oenb_mprj[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_413 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2006 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_498 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[107\]_A user_to_mprj_in_gates\[107\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__415__A _415_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[33\]_A _497_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_697 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[51\]_B la_buf_enable\[51\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output723_A output723/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_391 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_380 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2349 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1615 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2073 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[68\] user_to_mprj_in_gates\[68\]/Y user_to_mprj_in_gates\[68\]/B
+ input96/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_53_505 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[123\]_B mprj_logic_high_inst/HI[453] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_273 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[24\]_A _488_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[42\]_B la_buf_enable\[42\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput207 la_data_out_mprj[52] _516_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput218 la_data_out_mprj[62] _526_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput229 la_data_out_mprj[72] _536_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_9_1283 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1996 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[114\]_B mprj_logic_high_inst/HI[444] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[30\] vccd vssd user_to_mprj_in_gates\[30\]/B mprj_logic_high_inst/HI[360]
+ input311/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_38_2137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input287_A la_iena_mprj[124] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[15\]_A _479_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input454_A la_oenb_mprj[44] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1587 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input50_A la_data_out_core[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[33\]_B la_buf_enable\[33\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input621_A user_irq_core[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[2\]_A input310/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[100\]_A _363_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1957 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[105\]_B mprj_logic_high_inst/HI[435] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_1_2257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1845 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_777 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[38\] user_to_mprj_in_gates\[38\]/Y output686/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_30_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output673_A output673/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[24\]_B la_buf_enable\[24\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1649 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2063 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1412 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2157 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_833 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[93\]_A _356_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1945 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1989 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1675 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[15\]_B la_buf_enable\[15\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[78\] vccd vssd user_to_mprj_in_gates\[78\]/B mprj_logic_high_inst/HI[408]
+ input363/X vssd vccd sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[104\] _367_/Y la_oenb_core[104] mprj_logic_high_inst/HI[306]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[94\]_B mprj_logic_high_inst/HI[424] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
X_630_ _630_/A _630_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
Xla_buf_enable\[56\] la_buf\[56\]/TE _648_/A la_buf_enable\[56\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[34\] _626_/Y la_oenb_core[34] mprj_logic_high_inst/HI[236]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_29_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1821 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
X_561_ _561_/A _561_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_44_346 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_492_ _492_/A _492_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_input202_A la_data_out_mprj[48] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2145 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[84\]_A _347_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[118\]_TE mprj_logic_high_inst/HI[320] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input98_A la_data_out_core[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input571_A mprj_dat_i_user[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_932 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1936 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_69 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1204 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput571 input571/X mprj_dat_i_user[29] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_16
Xinput560 mprj_dat_i_user[19] input560/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
Xinput582 _432_/A mprj_dat_o_core[0] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_8
XFILLER_7_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[85\]_B mprj_logic_high_inst/HI[415] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput593 _433_/A mprj_dat_o_core[1] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_36_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[32\]_TE la_buf\[32\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_2098 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output790_A output790/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_571 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[75\]_A _338_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[17\]_TE mprj_logic_high_inst/HI[219] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1951 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__603__A _603_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[2\]_A input572/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1507 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_641 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[76\]_B mprj_logic_high_inst/HI[406] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1253 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[2\]_A input54/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_850 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[66\]_A _329_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1704 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[0\]_TE la_buf\[0\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__513__A _513_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_55 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1483 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_456 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input152_A la_data_out_mprj[118] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[67\]_B mprj_logic_high_inst/HI[397] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[55\]_TE la_buf\[55\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_613_ _613_/Y _613_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input417_A la_oenb_mprj[126] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input13_A la_data_out_core[108] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[61\] _525_/Y la_data_in_core[61] la_buf\[61\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_544_ _544_/Y _544_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
X_475_ _475_/Y _475_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_2_1695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1506 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[57\]_A _649_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_523 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1837 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[25\] _425_/Y mprj_adr_o_user[25] mprj_adr_buf\[25\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA__423__A _423_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_773 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1001 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output636_A output636/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1619 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2252 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1089 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[58\]_B mprj_logic_high_inst/HI[388] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1437 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[50\] user_to_mprj_in_gates\[50\]/Y user_to_mprj_in_gates\[50\]/B
+ input77/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
Xinput390 _364_/A la_oenb_mprj[101] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_52_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_861 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[48\]_A _640_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2037 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__333__A _333_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[78\]_TE la_buf\[78\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input5_A la_data_out_core[100] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1590 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[49\]_B mprj_logic_high_inst/HI[379] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2177 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_11 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_22 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_102 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2084 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__508__A _508_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_55 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_44 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_327 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_33 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_88 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_77 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_66 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_99 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1225 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[39\]_A _631_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[19\] la_buf\[19\]/TE _611_/A la_buf_enable\[19\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_13_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input367_A la_iena_mprj[81] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_irq_gates\[2\] user_irq_gates\[2\]/Y user_irq_gates\[2\]/B input623/X vssd vccd
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_46_2088 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input534_A mprj_adr_o_core[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1365 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2331 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[124\] la_buf\[124\]/TE _387_/A la_buf_enable\[124\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_8_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[27\]_TE mprj_dat_buf\[27\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_441 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2182 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_527_ _527_/Y _527_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_2_1481 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__418__A _418_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[6\]_TE mprj_logic_high_inst/HI[208] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
X_458_ _458_/Y _458_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_4
XFILLER_31_2324 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_389_ _389_/A _389_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_9_331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[20\] user_to_mprj_in_gates\[20\]/Y output667/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output753_A output753/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[98\] user_to_mprj_in_gates\[98\]/Y user_to_mprj_in_gates\[98\]/B
+ input129/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_29_2286 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[26\]_A _426_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[111\]_A_N _374_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1267 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[126\]_A_N _389_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_669 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_466 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[3\]_A _595_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1589 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput661 vccd vssd la_data_in_mprj[15] output661/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput672 vccd vssd la_data_in_mprj[25] output672/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput650 vccd vssd la_data_in_mprj[120] output650/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_43_1505 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput694 vccd vssd la_data_in_mprj[45] output694/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput683 vccd vssd la_data_in_mprj[35] output683/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_8_1123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[17\]_A _417_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1549 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[60\] vccd vssd user_to_mprj_in_gates\[60\]/B mprj_logic_high_inst/HI[390]
+ input344/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_mprj_sel_buf\[1\]_TE mprj_sel_buf\[1\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1994 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input115_A la_data_out_core[85] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput18 input18/X la_data_out_core[112] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_input80_A la_data_out_core[53] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1099 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_190 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_301 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input484_A la_oenb_mprj[71] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_802 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput29 input29/X la_data_out_core[122] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xla_buf\[24\] _488_/Y la_data_in_core[24] la_buf\[24\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_32_1965 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_buffers\[0\]_A user_irq_gates\[0\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_584 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[68\] user_to_mprj_in_gates\[68\]/Y output719/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_45_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1832 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[26\] user_wb_dat_gates\[26\]/Y input568/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_33_1729 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[13\] user_to_mprj_in_gates\[13\]/Y user_to_mprj_in_gates\[13\]/B
+ input36/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_buffers\[23\] output771/A user_wb_dat_gates\[23\]/Y vccd vssd vssd vccd
+ sky130_fd_sc_hd__inv_6
XANTENNA__611__A _611_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1393 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1869 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[124\] user_to_mprj_in_gates\[124\]/Y user_to_mprj_in_gates\[124\]/B
+ input31/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_3_80 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_761 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_249 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1031 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2032 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[10\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2076 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[103\]_TE la_buf\[103\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[18\]_TE mprj_adr_buf\[18\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1559 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__521__A _521_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[2\]_TE mprj_adr_buf\[2\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[64\] _656_/Y la_oenb_core[64] mprj_logic_high_inst/HI[266]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[86\] la_buf\[86\]/TE _349_/A la_buf_enable\[86\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_43_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[12\] _444_/Y mprj_dat_o_user[12] mprj_dat_buf\[12\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input232_A la_data_out_mprj[75] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_cyc_buf_A _393_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1841 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_411 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2018 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[50\]_TE mprj_logic_high_inst/HI[252] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_694 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_197 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__431__A _431_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[121\] user_to_mprj_in_gates\[121\]/Y output651/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_mprj_dat_buf\[6\]_TE mprj_dat_buf\[6\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2317 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output716_A output716/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[126\]_TE la_buf\[126\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1905 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__606__A _606_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1673 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[2\]_A _402_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__341__A _341_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_819 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2209 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput208 la_data_out_mprj[53] _517_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_wb_dat_buffers\[28\]_A user_wb_dat_gates\[28\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
Xinput219 la_data_out_mprj[63] _527_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_9_1251 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1295 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2149 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[73\]_TE mprj_logic_high_inst/HI[275] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[23\] vccd vssd user_to_mprj_in_gates\[23\]/B mprj_logic_high_inst/HI[353]
+ input303/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA__516__A _516_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1047 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input182_A la_data_out_mprj[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input447_A la_oenb_mprj[38] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input43_A la_data_out_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1831 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_buffers\[19\]_A user_wb_dat_gates\[19\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_43_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[2\]_B mprj_logic_high_inst/HI[332] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xla_buf\[91\] _555_/Y la_data_in_core[91] la_buf\[91\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input614_A mprj_iena_wb vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__426__A _426_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_233 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output666_A output666/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_473 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[80\] user_to_mprj_in_gates\[80\]/Y user_to_mprj_in_gates\[80\]/B
+ input110/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_6_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1953 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[84\]_A_N _347_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2075 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1424 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[123\]_B la_buf_enable\[123\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_889 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[96\]_TE mprj_logic_high_inst/HI[298] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_325 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[99\]_A_N _362_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[22\]_A_N _614_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__336__A _336_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_907 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1979 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[92\]_A input123/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[37\]_A_N _629_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_137 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[114\]_B la_buf_enable\[114\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_560_ _560_/Y _560_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_2_1833 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_358 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[27\] _619_/Y la_oenb_core[27] mprj_logic_high_inst/HI[229]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[49\] la_buf\[49\]/TE _641_/A la_buf_enable\[49\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[9\] _601_/Y la_oenb_core[9] mprj_logic_high_inst/HI[211]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_25_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_491_ _491_/Y _491_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_53_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[5\]_A user_wb_dat_gates\[5\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input397_A la_oenb_mprj[108] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1445 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[83\]_A input113/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input564_A mprj_dat_i_user[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[2\] _466_/Y la_data_in_core[2] la_buf\[2\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_49_2053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_944 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1142 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1175 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1733 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2309 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput572 mprj_dat_i_user[2] input572/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
Xinput561 mprj_dat_i_user[1] input561/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
Xinput550 mprj_dat_i_user[0] input550/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_la_buf\[8\]_A _472_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1788 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[105\]_B la_buf_enable\[105\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput583 _442_/A mprj_dat_o_core[10] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput594 mprj_dat_o_core[20] _452_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_39_1009 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[50\] user_to_mprj_in_gates\[50\]/Y output700/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output783_A output783/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1632 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1621 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[74\]_A input103/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1963 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1425 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[2\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_130 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2233 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[2\]_B user_to_mprj_in_gates\[2\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1565 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_862 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[65\]_A input93/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[90\] vccd vssd user_to_mprj_in_gates\[90\]/B mprj_logic_high_inst/HI[420]
+ input377/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_46_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_925 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input145_A la_data_out_mprj[111] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_612_ _612_/A _612_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_29_163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input312_A la_iena_mprj[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_133 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_543_ _543_/Y _543_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_53_2219 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_474_ _474_/Y _474_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf\[54\] _518_/Y la_data_in_core[54] la_buf\[54\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[126\] vccd vssd user_to_mprj_in_gates\[126\]/B mprj_logic_high_inst/HI[456]
+ input289/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_13_531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1974 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[56\]_A input83/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[110\] _574_/Y la_data_in_core[110] la_buf\[110\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xmprj_adr_buf\[18\] _418_/Y mprj_adr_o_user[18] mprj_adr_buf\[18\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_5_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1057 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[98\] user_to_mprj_in_gates\[98\]/Y output752/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output629_A output629/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2264 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput380 vssd vccd input380/X la_iena_mprj[93] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1416 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[6\]_A user_to_mprj_in_gates\[6\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput391 _365_/A la_oenb_mprj[102] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xuser_to_mprj_in_gates\[43\] user_to_mprj_in_gates\[43\]/Y input69/X user_to_mprj_in_gates\[43\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_buffers\[8\] output786/A user_wb_dat_gates\[8\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_16_391 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2185 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[47\]_A input73/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__614__A _614_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1771 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[5\] user_to_mprj_in_gates\[5\]/Y input87/X user_to_mprj_in_gates\[5\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_45_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[108\]_TE mprj_logic_high_inst/HI[310] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1051 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_12 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1972 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_637 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_56 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_45 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_34 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_89 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_78 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_67 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[38\]_A input63/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__524__A _524_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[122\]_A input29/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[94\] _357_/Y la_oenb_core[94] mprj_logic_high_inst/HI[296]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_2_733 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input262_A la_iena_mprj[101] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[22\]_TE la_buf\[22\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1907 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_221 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1631 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input527_A mprj_adr_o_core[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[7\] vccd vssd user_to_mprj_in_gates\[7\]/B mprj_logic_high_inst/HI[337]
+ input365/X vssd vccd sky130_fd_sc_hd__and2_1
Xla_buf_enable\[117\] la_buf\[117\]/TE _380_/A la_buf_enable\[117\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_8_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_667 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_526_ _526_/Y _526_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_45_497 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_457_ _457_/A _457_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_20_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2336 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_388_ _388_/Y _388_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_gates\[29\]_A input53/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1613 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[113\]_A input19/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__434__A _434_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[13\] user_to_mprj_in_gates\[13\]/Y output659/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_29_2210 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output746_A output746/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_409 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_943 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1213 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__609__A _609_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_478 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_681 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__344__A _344_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_A input9/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1134 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[45\]_TE la_buf\[45\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput662 vccd vssd la_data_in_mprj[16] output662/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput640 vccd vssd la_data_in_mprj[111] output640/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput651 vccd vssd la_data_in_mprj[121] output651/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput695 vccd vssd la_data_in_mprj[46] output695/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput673 vccd vssd la_data_in_mprj[26] output673/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput684 vccd vssd la_data_in_mprj[36] output684/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_8_1135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[53\] vccd vssd user_to_mprj_in_gates\[53\]/B mprj_logic_high_inst/HI[383]
+ input336/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_28_921 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1909 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__519__A _519_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input108_A la_data_out_core[79] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[31\] la_buf\[31\]/TE _623_/A la_buf_enable\[31\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_in_buffers\[5\] user_to_mprj_in_gates\[5\]/Y output710/A vccd vssd vssd
+ vccd sky130_fd_sc_hd__clkinv_4
XFILLER_19_1799 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1619 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xinput19 input19/X la_data_out_core[113] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_32_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input477_A la_oenb_mprj[65] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input73_A la_data_out_core[47] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[17\] _481_/Y la_data_in_core[17] la_buf\[17\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_6_357 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1141 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2195 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__429__A _429_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1844 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_509_ _509_/A _509_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_21_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output696_A output696/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[68\]_TE la_buf\[68\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[19\] user_wb_dat_gates\[19\]/Y input560/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_6_891 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[2\]_B la_buf_enable\[2\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[16\] user_wb_dat_gates\[16\]/Y output763/A vccd vssd vssd vccd
+ sky130_fd_sc_hd__clkinv_4
XFILLER_29_2095 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2009 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_92 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[126\]_A input289/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[117\] user_to_mprj_in_gates\[117\]/Y user_to_mprj_in_gates\[117\]/B
+ input23/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_42_1583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__339__A _339_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1043 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_607 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2088 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[17\]_TE mprj_dat_buf\[17\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_349 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[127\] _390_/Y la_oenb_core[127] mprj_logic_high_inst/HI[329]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[79\] la_buf\[79\]/TE _342_/A la_buf_enable\[79\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[57\] _649_/Y la_oenb_core[57] mprj_logic_high_inst/HI[259]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[117\]_A input279/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input225_A la_data_out_mprj[69] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1897 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_721 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_467 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input594_A mprj_dat_o_core[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[110\]_A_N _373_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[125\]_A_N _388_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[114\] user_to_mprj_in_gates\[114\]/Y output643/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_38_537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[80\] user_to_mprj_in_gates\[80\]/Y output733/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_output709_A output709/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[108\]_A input269/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_529 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_518 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_581 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2217 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__622__A _622_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput209 la_data_out_mprj[54] _518_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_42_2081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[16\] vccd vssd user_to_mprj_in_gates\[16\]/B mprj_logic_high_inst/HI[346]
+ input295/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_16_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_768 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_757 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[30\]_A input311/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1059 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__532__A _532_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input175_A la_data_out_mprj[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_157 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input342_A la_iena_mprj[59] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[97\]_A input384/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input36_A la_data_out_core[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[84\] _548_/Y la_data_in_core[84] la_buf\[84\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_1_2237 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input607_A mprj_dat_o_core[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_245 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[21\]_A input301/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2261 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_492 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1593 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__442__A _442_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output659_A output659/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[73\] user_to_mprj_in_gates\[73\]/Y user_to_mprj_in_gates\[73\]/B
+ input102/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[88\]_A input374/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1013 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1725 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__617__A _617_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1925 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[12\]_A input291/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_256 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[92\]_B user_to_mprj_in_gates\[92\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA__352__A _352_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[79\]_A input364/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[40\]_TE mprj_logic_high_inst/HI[242] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1812 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1981 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_389 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1795 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1856 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__527__A _527_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_490_ _490_/A _490_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_44_77 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_735 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input292_A la_iena_mprj[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[83\]_B user_to_mprj_in_gates\[83\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input557_A mprj_dat_i_user[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2065 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[116\]_TE la_buf\[116\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_477 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1154 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput573 mprj_dat_i_user[30] input573/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
Xinput562 input562/X mprj_dat_i_user[20] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_16
Xinput551 mprj_dat_i_user[10] input551/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_2170 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput540 vccd vssd _430_/A mprj_adr_o_core[30] vssd vccd sky130_fd_sc_hd__buf_2
Xinput584 _443_/A mprj_dat_o_core[11] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput595 mprj_dat_o_core[21] _453_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_35_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__437__A _437_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_551 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[43\] user_to_mprj_in_gates\[43\]/Y output692/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_34_1644 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output776_A output776/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[74\]_B user_to_mprj_in_gates\[74\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_8_783 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[63\]_TE mprj_logic_high_inst/HI[265] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__347__A _347_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1777 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1154 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[65\]_B user_to_mprj_in_gates\[65\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[83\] vccd vssd user_to_mprj_in_gates\[83\]/B mprj_logic_high_inst/HI[413]
+ input369/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_49_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[61\] la_buf\[61\]/TE _653_/A la_buf_enable\[61\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_45_613 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_611_ _611_/Y _611_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_buffers\[50\]_A user_to_mprj_in_gates\[50\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input138_A la_data_out_mprj[105] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_542_ _542_/Y _542_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_33_819 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_359 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input305_A la_iena_mprj[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_189 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_473_ _473_/Y _473_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_2_1686 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_543 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[47\] _511_/Y la_data_in_core[47] la_buf\[47\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_40_340 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1986 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1953 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[83\]_A_N _346_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[119\] vccd vssd user_to_mprj_in_gates\[119\]/B mprj_logic_high_inst/HI[449]
+ input281/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_13_587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[56\]_B user_to_mprj_in_gates\[56\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[90\]_A _554_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[86\]_TE mprj_logic_high_inst/HI[288] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[98\]_A_N _361_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2160 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[103\] _567_/Y la_data_in_core[103] la_buf\[103\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_42_1913 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[21\]_A_N _613_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_992 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[41\]_A user_to_mprj_in_gates\[41\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput370 vssd vccd input370/X la_iena_mprj[84] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput381 vssd vccd input381/X la_iena_mprj[94] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1428 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput392 _366_/A la_oenb_mprj[103] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_la_buf_enable\[36\]_A_N _628_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1152 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[36\] user_to_mprj_in_gates\[36\]/Y user_to_mprj_in_gates\[36\]/B
+ input61/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_52_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[47\]_B user_to_mprj_in_gates\[47\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[81\]_A _545_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__630__A _630_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2293 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_440 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1063 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[32\]_A user_to_mprj_in_gates\[32\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_39_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_13 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_46 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_35 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_24 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_79 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_68 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_57 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_693 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[99\]_A user_to_mprj_in_gates\[99\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[38\]_B user_to_mprj_in_gates\[38\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1574 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[122\]_B user_to_mprj_in_gates\[122\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[72\]_A _536_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[90\]_B la_buf_enable\[90\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__540__A _540_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[87\] _350_/Y la_oenb_core[87] mprj_logic_high_inst/HI[289]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_29_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_200 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_211 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input255_A la_data_out_mprj[96] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_39 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[23\]_A user_to_mprj_in_gates\[23\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input422_A la_oenb_mprj[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1895 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1687 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[31\]_A input574/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_525_ _525_/A _525_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_53_2028 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[126\]_A _590_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_456_ _456_/Y _456_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_4
X_387_ _387_/A _387_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_2348 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[29\]_B user_to_mprj_in_gates\[29\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_B user_to_mprj_in_gates\[113\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_9_355 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[63\]_A _527_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[30\] _430_/Y mprj_adr_o_user[30] mprj_adr_buf\[30\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[81\]_B la_buf_enable\[81\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__450__A _450_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2222 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output641_A output641/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output739_A output739/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2062 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[14\]_A user_to_mprj_in_gates\[14\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_432 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[22\]_A input564/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[117\]_A _581_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2259 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__625__A _625_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_B user_to_mprj_in_gates\[104\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[54\]_A _518_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[72\]_B la_buf_enable\[72\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_wb_ena_buf_A input614/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__360__A _360_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput663 vccd vssd la_data_in_mprj[17] output663/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput630 vccd vssd la_data_in_mprj[102] output630/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput641 vccd vssd la_data_in_mprj[112] output641/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput652 vccd vssd la_data_in_mprj[122] output652/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_28_1031 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput696 vccd vssd la_data_in_mprj[47] output696/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput685 vccd vssd la_data_in_mprj[37] output685/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput674 vccd vssd la_data_in_mprj[27] output674/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_8_1103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_stb_buf_A _394_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1147 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[46\] vccd vssd user_to_mprj_in_gates\[46\]/B mprj_logic_high_inst/HI[376]
+ input328/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_28_977 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[13\]_A input554/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1781 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[119\]_A user_to_mprj_in_gates\[119\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[108\]_A _572_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[24\] la_buf\[24\]/TE _616_/A la_buf_enable\[24\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA__535__A _535_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[45\]_A _509_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input372_A la_iena_mprj[86] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_387 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input66_A la_data_out_core[40] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[63\]_B la_buf_enable\[63\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1429 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_553 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_597 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_402 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1589 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_273 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_508_ _508_/Y _508_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA__445__A _445_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_439_ _439_/Y _439_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_output689_A output689/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[36\]_A _500_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[54\]_B la_buf_enable\[54\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_881 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[121\]_A _384_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[126\]_B mprj_logic_high_inst/HI[456] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_37_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_240 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1055 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1077 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1088 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_917 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[12\]_TE la_buf\[12\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_991 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__355__A _355_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_641 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[27\]_A _491_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[45\]_B la_buf_enable\[45\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_328 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[112\]_A _375_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1337 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_11 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[117\]_B mprj_logic_high_inst/HI[447] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input120_A la_data_out_core[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input218_A la_data_out_mprj[62] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_273 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input587_A mprj_dat_o_core[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[18\]_A _482_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[1\] input561/X user_wb_ack_gate/B user_wb_dat_gates\[1\]/Y vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_8
Xuser_to_mprj_in_ena_buf\[101\] vccd vssd user_to_mprj_in_gates\[101\]/B mprj_logic_high_inst/HI[431]
+ input262/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_7_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[36\]_B la_buf_enable\[36\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[5\]_A input343/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[103\]_A _366_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[107\] user_to_mprj_in_gates\[107\]/Y output635/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_38_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[108\]_B mprj_logic_high_inst/HI[438] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_38_549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[73\] user_to_mprj_in_gates\[73\]/Y output725/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_4_1353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[35\]_TE la_buf\[35\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[31\] user_wb_dat_gates\[31\]/Y input574/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_21_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1815 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[27\]_B la_buf_enable\[27\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[6\] _438_/Y mprj_dat_o_user[6] mprj_dat_buf\[6\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_1657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1128 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2093 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_733 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_210 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[96\]_A _359_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_416 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[30\]_B mprj_logic_high_inst/HI[360] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[3\]_TE la_buf\[3\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_482 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[18\]_B la_buf_enable\[18\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_637 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_125 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input168_A la_data_out_mprj[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[20\]_A _612_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[91\] la_buf\[91\]/TE _354_/A la_buf_enable\[91\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_7_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[97\]_B mprj_logic_high_inst/HI[427] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[58\]_TE la_buf\[58\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1719 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input335_A la_iena_mprj[52] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input29_A la_data_out_core[122] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[77\] _541_/Y la_data_in_core[77] la_buf\[77\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input502_A la_oenb_mprj[88] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[87\]_A _350_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[21\]_B mprj_logic_high_inst/HI[351] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1900 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[11\]_A _603_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output721_A output721/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[88\]_B mprj_logic_high_inst/HI[418] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_24_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[66\] user_to_mprj_in_gates\[66\]/Y user_to_mprj_in_gates\[66\]/B
+ input94/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_38_357 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[78\]_A _341_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[12\]_B mprj_logic_high_inst/HI[342] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_268 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__633__A _633_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[5\]_A input577/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[79\]_B mprj_logic_high_inst/HI[409] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1072 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1307 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_79 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[5\]_A input87/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1868 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[69\]_A _332_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[124\]_A_N _387_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_585 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__543__A _543_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input285_A la_iena_mprj[122] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input452_A la_oenb_mprj[42] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1166 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput530 vccd vssd _421_/A mprj_adr_o_core[21] vssd vccd sky130_fd_sc_hd__buf_2
Xinput563 mprj_dat_i_user[21] input563/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
Xinput552 mprj_dat_i_user[11] input552/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
Xinput541 mprj_adr_o_core[31] _431_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput574 mprj_dat_i_user[31] input574/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
XFILLER_48_677 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_305 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput585 _444_/A mprj_dat_o_core[12] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput596 mprj_dat_o_core[22] _454_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_51_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[9\]_TE mprj_logic_high_inst/HI[211] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1389 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_533 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[36\] user_to_mprj_in_gates\[36\]/Y output684/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA__453__A _453_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output671_A output671/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output769_A output769/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_751 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_600 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1785 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_113 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__628__A _628_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_157 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_872 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__363__A _363_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1133 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_739 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[76\] vccd vssd user_to_mprj_in_gates\[76\]/B mprj_logic_high_inst/HI[406]
+ input361/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_28_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1251 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[102\] _365_/Y la_oenb_core[102] mprj_logic_high_inst/HI[304]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_610_ _610_/Y _610_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA__538__A _538_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_541_ _541_/A _541_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[32\] _624_/Y la_oenb_core[32] mprj_logic_high_inst/HI[234]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_2_1643 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1632 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[54\] la_buf\[54\]/TE _646_/A la_buf_enable\[54\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
X_472_ _472_/A _472_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_input200_A la_data_out_mprj[46] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_691 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_853 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[20\]_A _452_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_190 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_352 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input96_A la_data_out_core[68] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1998 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1829 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_721 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1819 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput360 vssd vccd input360/X la_iena_mprj[75] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput371 vssd vccd input371/X la_iena_mprj[85] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1565 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__448__A _448_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput382 vssd vccd input382/X la_iena_mprj[95] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput393 vccd vssd _367_/A la_oenb_mprj[104] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_51_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_691 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[11\]_A _443_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[29\] user_to_mprj_in_gates\[29\]/Y user_to_mprj_in_gates\[29\]/B
+ input53/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_16_371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1453 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_385 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1475 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[30\]_TE mprj_logic_high_inst/HI[232] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[29\]_A _429_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1257 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__358__A _358_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_102 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1075 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[6\]_A _598_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_47 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_14 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_25 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_36 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_58 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[106\]_TE la_buf\[106\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_69 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1586 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[5\]_TE mprj_adr_buf\[5\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1283 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[28\] _460_/Y mprj_dat_o_user[28] mprj_dat_buf\[28\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input150_A la_data_out_mprj[116] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input248_A la_data_out_mprj[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input415_A la_oenb_mprj[124] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input11_A la_data_out_core[106] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[31\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_989 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_524_ _524_/A _524_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_33_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_455_ _455_/Y _455_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_6
XFILLER_53_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[53\]_TE mprj_logic_high_inst/HI[255] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_386_ _386_/Y _386_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_31_2305 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[23\] _423_/Y mprj_adr_o_user[23] mprj_adr_buf\[23\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_29_2234 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[9\]_TE mprj_dat_buf\[9\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_573 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output634_A output634/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2041 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput190 vccd vssd la_data_out_mprj[37] _501_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[22\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_617 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_691 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1840 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[8\] la_buf\[8\]/TE _600_/A la_buf_enable\[8\]/B vssd vccd vssd vccd
+ sky130_fd_sc_hd__and2b_1
XANTENNA__641__A _641_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1600 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2209 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_wb_ena_buf_B user_to_mprj_wb_ena_buf/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput631 vccd vssd la_data_in_mprj[103] output631/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput642 vccd vssd la_data_in_mprj[113] output642/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput653 vccd vssd la_data_in_mprj[123] output653/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput697 vccd vssd la_data_in_mprj[48] output697/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput686 vccd vssd la_data_in_mprj[38] output686/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput664 vccd vssd la_data_in_mprj[18] output664/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput675 vccd vssd la_data_in_mprj[28] output675/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_8_1115 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input3_A caravel_rstn vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1065 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[82\]_A_N _345_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[91\]_TE la_buf\[91\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[13\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[76\]_TE mprj_logic_high_inst/HI[278] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[39\] vccd vssd user_to_mprj_in_gates\[39\]/B mprj_logic_high_inst/HI[369]
+ input320/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_3_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[97\]_A_N _360_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2040 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_67 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[17\] la_buf\[17\]/TE _609_/A la_buf_enable\[17\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf_enable\[20\]_A_N _612_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_867 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1957 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input198_A la_data_out_mprj[44] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__551__A _551_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_399 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[35\]_A_N _627_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input365_A la_iena_mprj[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input59_A la_data_out_core[34] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_irq_gates\[0\] user_irq_gates\[0\]/Y user_irq_gates\[0\]/B input621/X vssd vccd
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_26_1739 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2203 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input532_A mprj_adr_o_core[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[122\] la_buf\[122\]/TE _385_/A la_buf_enable\[122\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_4_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_414 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_499 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_507_ _507_/Y _507_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_53_1114 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_438_ _438_/A _438_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
X_369_ _369_/Y _369_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_31_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__461__A _461_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output751_A output751/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[96\] user_to_mprj_in_gates\[96\]/Y user_to_mprj_in_gates\[96\]/B
+ input127/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_42_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[99\]_TE mprj_logic_high_inst/HI[301] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_219 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_753 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_797 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__636__A _636_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[5\]_A _405_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1378 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__371__A _371_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1698 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2164 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_23 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1051 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_753 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input113_A la_data_out_core[83] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__546__A _546_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1309 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_613 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input482_A la_oenb_mprj[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[22\] _486_/Y la_data_in_core[22] la_buf\[22\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_7_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_189 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_841 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[5\]_B mprj_logic_high_inst/HI[335] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_517 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_stb_buf_TE mprj_stb_buf/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[66\] user_to_mprj_in_gates\[66\]/Y output717/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA__456__A _456_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[24\] user_wb_dat_gates\[24\]/Y input566/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_2
Xuser_to_mprj_in_gates\[11\] user_to_mprj_in_gates\[11\]/Y input26/X user_to_mprj_in_gates\[11\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_50_1821 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_buffers\[21\] output769/A user_wb_dat_gates\[21\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1182 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[126\]_B la_buf_enable\[126\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[122\] user_to_mprj_in_gates\[122\]/Y user_to_mprj_in_gates\[122\]/B
+ input29/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_37_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1967 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__366__A _366_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_277 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_428 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_47 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[95\]_A input126/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1197 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_104 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[31\]_TE mprj_adr_buf\[31\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[62\] _654_/Y la_oenb_core[62] mprj_logic_high_inst/HI[264]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[84\] la_buf\[84\]/TE _347_/A la_buf_enable\[84\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_7_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[117\]_B la_buf_enable\[117\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[10\] _442_/Y mprj_dat_o_user[10] mprj_dat_buf\[10\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input230_A la_data_out_mprj[73] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input328_A la_iena_mprj[46] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_553 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_buffers\[8\]_A user_wb_dat_gates\[8\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_299 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[86\]_A input116/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_999 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[126\] _590_/Y la_data_in_core[126] la_buf\[126\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_28_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_682 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[108\]_B la_buf_enable\[108\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[10\]_A input15/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output714_A output714/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[59\] user_to_mprj_in_gates\[59\]/Y user_to_mprj_in_gates\[59\]/B
+ input86/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_39_1705 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_572 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2185 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[77\]_A input106/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1337 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[5\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1477 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[5\]_B user_to_mprj_in_gates\[5\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1847 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_553 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[21\] vccd vssd user_to_mprj_in_gates\[21\]/B mprj_logic_high_inst/HI[351]
+ input301/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[68\]_A input96/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[25\]_TE la_buf\[25\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_413 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input180_A la_data_out_mprj[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input278_A la_iena_mprj[116] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input41_A la_data_out_core[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input445_A la_oenb_mprj[36] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1090 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput520 vccd vssd _412_/A mprj_adr_o_core[12] vssd vccd sky130_fd_sc_hd__buf_2
Xinput553 mprj_dat_i_user[12] input553/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
Xinput564 mprj_dat_i_user[22] input564/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
XFILLER_48_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput542 vccd vssd _403_/A mprj_adr_o_core[3] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input612_A mprj_dat_o_core[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput531 mprj_adr_o_core[22] _422_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput575 vccd vssd input575/X mprj_dat_i_user[3] vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2036 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput586 _445_/A mprj_dat_o_core[13] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput597 vccd vssd _455_/A mprj_dat_o_core[23] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_29_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2069 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_501 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_A input86/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[29\] user_to_mprj_in_gates\[29\]/Y output676/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_32_2093 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output664_A output664/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_763 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_612 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[9\]_A user_to_mprj_in_gates\[9\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_38_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_884 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__644__A _644_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[48\]_TE la_buf\[48\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1281 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1855 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1167 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1590 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[69\] vccd vssd user_to_mprj_in_gates\[69\]/B mprj_logic_high_inst/HI[399]
+ input353/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_40_1105 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1859 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
X_540_ _540_/Y _540_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_40_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1594 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_339 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[47\] la_buf\[47\]/TE _639_/A la_buf_enable\[47\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[25\] _617_/Y la_oenb_core[25] mprj_logic_high_inst/HI[227]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[7\] _599_/Y la_oenb_core[7] mprj_logic_high_inst/HI[209]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_471_ _471_/Y _471_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_25_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2091 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_523 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[125\]_A input32/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__554__A _554_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input395_A la_oenb_mprj[106] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input89_A la_data_out_core[61] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input562_A mprj_dat_i_user[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[0\] _464_/Y la_data_in_core[0] la_buf\[0\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_4_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1185 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput350 vssd vccd input350/X la_iena_mprj[66] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput361 vssd vccd input361/X la_iena_mprj[76] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput372 vssd vccd input372/X la_iena_mprj[86] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_36_637 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_90 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput383 vssd vccd input383/X la_iena_mprj[96] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput394 vccd vssd _368_/A la_oenb_mprj[105] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_35_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_383 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2144 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__464__A _464_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_A input22/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output781_A output781/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[123\]_A_N _386_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1308 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1010 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__639__A _639_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1087 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_497 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_114 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1953 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_26 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_37 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_59 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_48 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__374__A _374_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[107\]_A input12/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1554 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_69 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2026 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_268 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_217 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input143_A la_data_out_mprj[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__549__A _549_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2120 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2153 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input310_A la_iena_mprj[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input408_A la_oenb_mprj[118] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_523_ _523_/Y _523_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_33_629 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
X_454_ _454_/Y _454_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_4
XFILLER_26_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[52\] _516_/Y la_data_in_core[52] la_buf\[52\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[124\] vccd vssd user_to_mprj_in_gates\[124\]/B mprj_logic_high_inst/HI[454]
+ input287/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_13_331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_662 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_385_ _385_/Y _385_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_35_1785 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1763 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1501 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[16\] _416_/Y mprj_adr_o_user[16] mprj_adr_buf\[16\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_42_1701 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output627_A output627/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[96\] user_to_mprj_in_gates\[96\]/Y output750/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_42_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__459__A _459_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1341 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2097 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xmprj_rstn_buf input3/X user_reset mprj_rstn_buf/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xinput180 vccd vssd la_data_out_mprj[28] _492_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_1789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput191 vssd vccd _502_/A la_data_out_mprj[38] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_36_456 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[41\] user_to_mprj_in_gates\[41\]/Y user_to_mprj_in_gates\[41\]/B
+ input67/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_buffers\[6\] output784/A user_wb_dat_gates\[6\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_52_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[5\]_B la_buf_enable\[5\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2324 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1612 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput632 vccd vssd la_data_in_mprj[104] output632/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput643 vccd vssd la_data_in_mprj[114] output643/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput654 vccd vssd la_data_in_mprj[124] output654/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput687 vccd vssd la_data_in_mprj[39] output687/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput665 vccd vssd la_data_in_mprj[19] output665/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput676 vccd vssd la_data_in_mprj[29] output676/A vssd vccd sky130_fd_sc_hd__buf_2
Xuser_to_mprj_in_gates\[3\] user_to_mprj_in_gates\[3\]/Y input65/X user_to_mprj_in_gates\[3\]/B
+ vssd vccd vssd vccd sky130_fd_sc_hd__nand2_2
Xoutput698 vccd vssd la_data_in_mprj[49] output698/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_25_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__369__A _369_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[121\]_TE mprj_logic_high_inst/HI[323] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_445 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_949 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[60\]_A input344/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_79 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_879 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[92\] _355_/Y la_oenb_core[92] mprj_logic_high_inst/HI[294]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_30_1682 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input260_A la_iena_mprj[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input358_A la_iena_mprj[73] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input525_A mprj_adr_o_core[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[5\] vccd vssd user_to_mprj_in_gates\[5\]/B mprj_logic_high_inst/HI[335]
+ input343/X vssd vccd sky130_fd_sc_hd__and2_1
Xla_buf_enable\[115\] la_buf\[115\]/TE _378_/A la_buf_enable\[115\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_oen_buffers\[20\]_TE mprj_logic_high_inst/HI[222] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_506_ _506_/Y _506_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_33_426 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[51\]_A input334/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_437_ _437_/A _437_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_14_651 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1159 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_368_ _368_/A _368_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_1413 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[11\] output649/A user_to_mprj_in_gates\[11\]/Y vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_6
XANTENNA_output744_A output744/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_40 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[89\] user_to_mprj_in_gates\[89\]/Y user_to_mprj_in_gates\[89\]/B
+ input119/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_42_2265 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1553 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1193 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1851 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1302 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1895 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[42\]_A input324/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__652__A _652_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2176 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[43\]_TE mprj_logic_high_inst/HI[245] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_35 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1740 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[51\] vccd vssd user_to_mprj_in_gates\[51\]/B mprj_logic_high_inst/HI[381]
+ input334/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_47_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1795 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xmprj_cyc_buf _393_/Y mprj_cyc_o_user mprj_cyc_buf/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input106_A la_data_out_core[77] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_245 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[33\]_A input314/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[3\] user_to_mprj_in_gates\[3\]/Y output688/A vccd vssd vssd
+ vccd sky130_fd_sc_hd__clkinv_4
XFILLER_42_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_470 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_632 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__562__A _562_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input475_A la_oenb_mprj[63] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input71_A la_data_out_core[45] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[119\]_TE la_buf\[119\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[15\] _479_/Y la_data_in_core[15] la_buf\[15\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_7_669 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[0\]_A _432_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_831 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_897 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_396 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2001 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[8\] _408_/Y mprj_adr_o_user[8] mprj_adr_buf\[8\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[59\] user_to_mprj_in_gates\[59\]/Y output709/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[24\]_A input304/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output694_A output694/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1811 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__472__A _472_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[17\] user_wb_dat_gates\[17\]/Y input558/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf_enable\[81\]_A_N _344_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[81\]_TE la_buf\[81\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_680 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[14\] output761/A user_wb_dat_gates\[14\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[66\]_TE mprj_logic_high_inst/HI[268] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[96\]_A_N _359_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1194 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[115\] user_to_mprj_in_gates\[115\]/Y user_to_mprj_in_gates\[115\]/B
+ input21/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA__647__A _647_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_510 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1419 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[34\]_A_N _626_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[15\]_A input294/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2309 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1608 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_749 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[95\]_B user_to_mprj_in_gates\[95\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA__382__A _382_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[49\]_A_N _641_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1739 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_clk2_buf_TE mprj_clk2_buf/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[99\] vccd vssd user_to_mprj_in_gates\[99\]/B mprj_logic_high_inst/HI[429]
+ input386/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_49_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[30\]_TE mprj_dat_buf\[30\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[125\] _388_/Y la_oenb_core[125] mprj_logic_high_inst/HI[327]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_7_1929 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[55\] _647_/Y la_oenb_core[55] mprj_logic_high_inst/HI[257]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_0_889 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[80\]_A user_to_mprj_in_gates\[80\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1169 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[77\] la_buf\[77\]/TE _340_/A la_buf_enable\[77\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_input223_A la_data_out_mprj[67] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[2\]_A input626/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__557__A _557_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1817 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input592_A mprj_dat_o_core[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[86\]_B user_to_mprj_in_gates\[86\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[89\]_TE mprj_logic_high_inst/HI[291] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_411 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[119\] _583_/Y la_data_in_core[119] la_buf\[119\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_10_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[112\] user_to_mprj_in_gates\[112\]/Y output641/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_3_694 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[10\]_B user_to_mprj_in_gates\[10\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[71\]_A user_to_mprj_in_gates\[71\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_output707_A output707/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__467__A _467_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_B user_to_mprj_in_gates\[77\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_30_793 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1647 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[62\]_A user_to_mprj_in_gates\[62\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__377__A _377_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_852 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[14\] vccd vssd user_to_mprj_in_gates\[14\]/B mprj_logic_high_inst/HI[344]
+ input293/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[68\]_B user_to_mprj_in_gates\[68\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_40_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2002 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input173_A la_data_out_mprj[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[100\]_A user_to_mprj_in_gates\[100\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_469 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input340_A la_iena_mprj[57] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input438_A la_oenb_mprj[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput510 _358_/A la_oenb_mprj[95] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_buffers\[53\]_A user_to_mprj_in_gates\[53\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput521 vccd vssd mprj_adr_o_core[13] _413_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input34_A la_data_out_core[127] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput554 mprj_dat_i_user[13] input554/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_48_635 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput543 mprj_adr_o_core[4] _404_/A vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
Xinput532 mprj_adr_o_core[23] _423_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput576 vccd vssd input576/X mprj_dat_i_user[4] vssd vccd sky130_fd_sc_hd__buf_6
Xinput565 mprj_dat_i_user[23] input565/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
Xla_buf\[82\] _546_/Y la_data_in_core[82] la_buf\[82\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_48_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput587 vccd vssd _446_/A mprj_dat_o_core[14] vssd vccd sky130_fd_sc_hd__buf_4
Xinput598 mprj_dat_o_core[24] _456_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_input605_A mprj_dat_o_core[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1314 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_893 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_B user_to_mprj_in_gates\[59\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[93\]_A _557_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_775 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output657_A output657/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[44\]_A user_to_mprj_in_gates\[44\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[71\] user_to_mprj_in_gates\[71\]/Y user_to_mprj_in_gates\[71\]/B
+ input100/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_41_1629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_189 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1525 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[21\]_TE mprj_adr_buf\[21\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_373 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1703 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1823 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[84\]_A _548_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1113 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1867 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1769 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_428 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[35\]_A user_to_mprj_in_gates\[35\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1985 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1827 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1297 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_178 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_690 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1573 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
X_470_ _470_/A _470_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[18\] _610_/Y la_oenb_core[18] mprj_logic_high_inst/HI[220]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_25_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[125\]_B user_to_mprj_in_gates\[125\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[75\]_A _539_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_579 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input388_A la_oenb_mprj[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input290_A la_iena_mprj[127] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[93\]_B la_buf_enable\[93\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input555_A mprj_dat_i_user[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__570__A _570_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1716 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[26\]_A user_to_mprj_in_gates\[26\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput340 vssd vccd input340/X la_iena_mprj[57] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput351 vssd vccd input351/X la_iena_mprj[67] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput362 vssd vccd input362/X la_iena_mprj[77] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput373 vssd vccd input373/X la_iena_mprj[87] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput384 vssd vccd input384/X la_iena_mprj[97] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput395 vccd vssd _369_/A la_oenb_mprj[106] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_35_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2281 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_599_ _599_/A _599_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_43_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[116\]_B user_to_mprj_in_gates\[116\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[41\] user_to_mprj_in_gates\[41\]/Y output690/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf\[66\]_A _530_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output774_A output774/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[84\]_B la_buf_enable\[84\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__480__A _480_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[17\]_A user_to_mprj_in_gates\[17\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1022 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[25\]_A input567/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_126 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[15\]_TE la_buf\[15\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_27 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_38 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_16 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__655__A _655_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_49 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[107\]_B user_to_mprj_in_gates\[107\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[57\]_A _521_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_1631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1090 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[75\]_B la_buf_enable\[75\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__390__A _390_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2038 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[81\] vccd vssd user_to_mprj_in_gates\[81\]/B mprj_logic_high_inst/HI[411]
+ input367/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_24_2303 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[16\]_A input557/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input136_A la_data_out_mprj[103] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_522_ _522_/A _522_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_input303_A la_iena_mprj[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__565__A _565_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_453_ _453_/Y _453_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_4
XFILLER_26_693 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[48\]_A _512_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_384_ _384_/Y _384_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf\[45\] _509_/Y la_data_in_core[45] la_buf\[45\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_51_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[117\] vccd vssd user_to_mprj_in_gates\[117\]/B mprj_logic_high_inst/HI[447]
+ input279/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_51_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[66\]_B la_buf_enable\[66\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_70 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_553 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[101\] _565_/Y la_data_in_core[101] la_buf\[101\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_9_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1757 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xinput170 vccd vssd la_data_out_mprj[19] _483_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput181 la_data_out_mprj[29] _493_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xuser_to_mprj_in_buffers\[89\] user_to_mprj_in_gates\[89\]/Y output742/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_7_1397 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[38\]_TE la_buf\[38\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput192 vssd vccd _503_/A la_data_out_mprj[39] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_36_468 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__475__A _475_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[34\] user_to_mprj_in_gates\[34\]/Y user_to_mprj_in_gates\[34\]/B
+ input59/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_51_449 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[39\]_A _503_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[57\]_B la_buf_enable\[57\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2336 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[124\]_A _387_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput633 vccd vssd la_data_in_mprj[105] output633/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput644 vccd vssd la_data_in_mprj[115] output644/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput688 vccd vssd la_data_in_mprj[3] output688/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput677 vccd vssd la_data_in_mprj[2] output677/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput666 vccd vssd la_data_in_mprj[1] output666/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput655 vccd vssd la_data_in_mprj[125] output655/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_25_1911 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput699 vccd vssd la_data_in_mprj[4] output699/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_41_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__385__A _385_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1715 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[60\]_B mprj_logic_high_inst/HI[390] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[6\]_TE la_buf\[6\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1330 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_807 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2097 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[48\]_B la_buf_enable\[48\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[115\]_A _378_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[85\] _348_/Y la_oenb_core[85] mprj_logic_high_inst/HI[287]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[50\]_A _642_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input253_A la_data_out_mprj[94] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_2111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input420_A la_oenb_mprj[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input518_A mprj_adr_o_core[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1504 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[108\] la_buf\[108\]/TE _371_/A la_buf_enable\[108\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
X_505_ _505_/Y _505_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_18_479 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1283 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_438 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[51\]_B mprj_logic_high_inst/HI[381] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_42_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[122\]_A_N _385_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_436_ _436_/Y _436_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
X_367_ _367_/Y _367_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf_enable\[39\]_B la_buf_enable\[39\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[8\]_A input376/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[41\]_A _633_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[106\]_A _369_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output737_A output737/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_766 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[42\]_B mprj_logic_high_inst/HI[372] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_32_471 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[32\]_A _624_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1752 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_47 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[99\]_A _362_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[44\] vccd vssd user_to_mprj_in_gates\[44\]/B mprj_logic_high_inst/HI[374]
+ input326/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_3_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[33\]_B mprj_logic_high_inst/HI[363] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[22\] la_buf\[22\]/TE _614_/A la_buf_enable\[22\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_23_482 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1701 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input468_A la_oenb_mprj[57] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input370_A la_iena_mprj[84] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input64_A la_data_out_core[39] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[23\]_A _615_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_821 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1491 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_854 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1367 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[24\]_B mprj_logic_high_inst/HI[354] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1509 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output687_A output687/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_419_ _419_/Y _419_/A vssd vccd vssd vccd sky130_fd_sc_hd__inv_16
XFILLER_14_471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_964 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[111\]_TE mprj_logic_high_inst/HI[313] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[14\]_A _606_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_692 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1212 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[108\] user_to_mprj_in_gates\[108\]/Y user_to_mprj_in_gates\[108\]/B
+ input13/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_37_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[10\]_A _410_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_522 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1682 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[15\]_B mprj_logic_high_inst/HI[345] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_33_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[8\]_A input580/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1505 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[10\]_TE mprj_logic_high_inst/HI[212] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[118\] _381_/Y la_oenb_core[118] mprj_logic_high_inst/HI[320]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_27_1847 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[8\]_A input120/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[48\] _640_/Y la_oenb_core[48] mprj_logic_high_inst/HI[250]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_47_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[2\]_B user_irq_ena_buf\[2\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_585 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input216_A la_data_out_mprj[60] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__573__A _573_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input585_A mprj_dat_o_core[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1575 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_445 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_673 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[105\] user_to_mprj_in_gates\[105\]/Y output633/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_43_1693 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[71\] user_to_mprj_in_gates\[71\]/Y output723/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_4_1142 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1991 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1197 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__483__A _483_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2321 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[33\]_TE mprj_logic_high_inst/HI[235] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1030 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1697 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[4\] _436_/Y mprj_dat_o_user[4] mprj_dat_buf\[4\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_29_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1170 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1722 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[109\]_TE la_buf\[109\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_897 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_525 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__393__A _393_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[8\]_TE mprj_adr_buf\[8\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input166_A la_data_out_mprj[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1655 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xinput500 vccd vssd _349_/A la_oenb_mprj[86] vssd vccd sky130_fd_sc_hd__buf_4
Xinput511 la_oenb_mprj[96] _359_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1705 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput555 mprj_dat_i_user[14] input555/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
XANTENNA__568__A _568_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2091 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input333_A la_iena_mprj[50] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput544 _405_/A mprj_adr_o_core[5] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput522 mprj_adr_o_core[14] _414_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput533 vccd vssd _424_/A mprj_adr_o_core[24] vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_input27_A la_data_out_core[120] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput566 mprj_dat_i_user[24] input566/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
Xinput577 mprj_dat_i_user[5] input577/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_48_669 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[80\]_A_N _343_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput588 vccd vssd _447_/A mprj_dat_o_core[15] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_5_2185 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[71\]_TE la_buf\[71\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input500_A la_oenb_mprj[86] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1484 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput599 vccd vssd mprj_dat_o_core[25] _457_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xla_buf\[75\] _539_/Y la_data_in_core[75] la_buf\[75\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[23\]_A _455_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[56\]_TE mprj_logic_high_inst/HI[258] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[30\]_A user_wb_dat_gates\[30\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_43_385 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[95\]_A_N _358_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_588 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[33\]_A_N _625_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1692 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[48\]_A_N _640_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_669 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__478__A _478_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[64\] user_to_mprj_in_gates\[64\]/Y user_to_mprj_in_gates\[64\]/B
+ input92/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_mprj_dat_buf\[14\]_A _446_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[21\]_A user_wb_dat_gates\[21\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_35_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_525 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[20\]_TE mprj_dat_buf\[20\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2140 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1423 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2091 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[94\]_TE la_buf\[94\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_102 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__388__A _388_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_113 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[79\]_TE mprj_logic_high_inst/HI[281] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1624 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[9\]_A _601_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[12\]_A user_wb_dat_gates\[12\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_25_385 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input283_A la_iena_mprj[120] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_245 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input450_A la_oenb_mprj[40] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1728 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_289 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input548_A mprj_adr_o_core[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput330 vssd vccd input330/X la_iena_mprj[48] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput341 vssd vccd input341/X la_iena_mprj[58] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput352 vssd vccd input352/X la_iena_mprj[68] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput363 vssd vccd input363/X la_iena_mprj[78] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_49_989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput374 vssd vccd input374/X la_iena_mprj[88] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput385 vssd vccd input385/X la_iena_mprj[98] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput396 _370_/A la_oenb_mprj[107] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_35_105 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1281 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_609 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_598_ _598_/Y _598_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_43_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_322 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[34\] user_to_mprj_in_gates\[34\]/Y output682/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output767_A output767/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_551 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_41 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_74 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_63 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_96 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[25\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_606 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_17 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_28 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_39 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1654 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_248 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[74\] vccd vssd user_to_mprj_in_gates\[74\]/B mprj_logic_high_inst/HI[404]
+ input359/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_28_1761 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1603 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[100\] _363_/Y la_oenb_core[100] mprj_logic_high_inst/HI[302]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_24_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[16\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1084 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input129_A la_data_out_core[98] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_959 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[30\] _622_/Y la_oenb_core[30] mprj_logic_high_inst/HI[232]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_18_639 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[52\] la_buf\[52\]/TE _644_/A la_buf_enable\[52\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_33_609 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_521_ _521_/A _521_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_2_1465 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2188 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_452_ _452_/Y _452_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_4
X_383_ _383_/A _383_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[1\]_A _465_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input498_A la_oenb_mprj[84] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_355 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input94_A la_data_out_core[66] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__581__A _581_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[38\] _502_/Y la_data_in_core[38] la_buf\[38\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_51_1077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[11\]_TE mprj_adr_buf\[11\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1619 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_gates\[1\]_A input622/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput171 la_data_out_mprj[1] _465_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput160 la_data_out_mprj[125] _589_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_49_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput193 la_data_out_mprj[3] _467_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput182 la_data_out_mprj[2] _466_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_51_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[27\] user_to_mprj_in_gates\[27\]/Y user_to_mprj_in_gates\[27\]/B
+ input51/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_32_697 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__491__A _491_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1898 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_196 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2348 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput634 vccd vssd la_data_in_mprj[106] output634/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput645 vccd vssd la_data_in_mprj[116] output645/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput667 vccd vssd la_data_in_mprj[20] output667/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput678 vccd vssd la_data_in_mprj[30] output678/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput656 vccd vssd la_data_in_mprj[126] output656/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput689 vccd vssd la_data_in_mprj[40] output689/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_41_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[8\]_A _408_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1342 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[78\] _341_/Y la_oenb_core[78] mprj_logic_high_inst/HI[280]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_46_1157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[26\] _458_/Y mprj_dat_o_user[26] mprj_dat_buf\[26\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_24_2123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_568 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input246_A la_data_out_mprj[88] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1630 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1516 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_403 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input413_A la_oenb_mprj[122] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__576__A _576_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_447 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
X_504_ _504_/A _504_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_42_973 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_435_ _435_/A _435_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_14_675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_366_ _366_/Y _366_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_35_1573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_830 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[21\] _421_/Y mprj_adr_o_user[21] mprj_adr_buf\[21\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[8\]_B mprj_logic_high_inst/HI[338] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_373 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output632_A output632/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[40\]_A input66/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1427 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1173 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__486__A _486_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_778 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_417 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[6\] la_buf\[6\]/TE _598_/A la_buf_enable\[6\]/B vssd vccd vssd vccd
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1993 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2009 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[31\]_A input56/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1764 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input1_A caravel_clk vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__396__A _396_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_767 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[37\] vccd vssd user_to_mprj_in_gates\[37\]/B mprj_logic_high_inst/HI[367]
+ input318/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[98\]_A input129/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[15\] la_buf\[15\]/TE _607_/A la_buf_enable\[15\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_23_494 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_605 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_667 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[28\]_TE la_buf\[28\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input196_A la_data_out_mprj[42] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_678 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_137 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input363_A la_iena_mprj[78] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2207 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input57_A la_data_out_core[32] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[22\]_A input46/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_866 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input530_A mprj_adr_o_core[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[120\] la_buf\[120\]/TE _383_/A la_buf_enable\[120\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_19_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1897 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_748 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[89\]_A input119/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_418_ _418_/A _418_/Y vssd vccd vssd vccd sky130_fd_sc_hd__inv_12
XFILLER_14_483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1911 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_349_ _349_/A _349_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_976 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1999 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1819 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1690 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[94\] user_to_mprj_in_gates\[94\]/Y user_to_mprj_in_gates\[94\]/B
+ input125/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_gates\[13\]_A input36/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1224 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1385 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1145 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_39 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[8\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[121\]_A_N _384_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2345 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[8\]_B user_to_mprj_in_gates\[8\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_48_829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1677 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input111_A la_data_out_core[81] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input209_A la_data_out_mprj[54] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1933 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1109 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input578_A mprj_dat_i_user[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input480_A la_oenb_mprj[68] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1565 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[20\] _484_/Y la_data_in_core[20] la_buf\[20\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_48_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_542 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_862 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[64\] user_to_mprj_in_gates\[64\]/Y output715/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_37_2155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[22\] user_wb_dat_gates\[22\]/Y input564/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_14_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1042 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1425 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[120\] user_to_mprj_in_gates\[120\]/Y user_to_mprj_in_gates\[120\]/B
+ input27/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_9_1087 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1734 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1182 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_309 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_501 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2253 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[110\]_A input272/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1841 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_272 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1115 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[60\] _652_/Y la_oenb_core[60] mprj_logic_high_inst/HI[262]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[82\] la_buf\[82\]/TE _345_/A la_buf_enable\[82\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xinput501 _350_/A la_oenb_mprj[87] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput512 _360_/A la_oenb_mprj[97] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_input159_A la_data_out_mprj[124] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput545 mprj_adr_o_core[6] _406_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput523 vccd vssd _415_/A mprj_adr_o_core[15] vssd vccd sky130_fd_sc_hd__buf_2
Xinput534 _425_/A mprj_adr_o_core[25] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput567 mprj_dat_i_user[25] input567/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
Xinput578 mprj_dat_i_user[6] input578/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
Xinput556 mprj_dat_i_user[15] input556/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
XFILLER_44_1981 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input326_A la_iena_mprj[44] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput589 _448_/A mprj_dat_o_core[16] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_oen_buffers\[101\]_TE mprj_logic_high_inst/HI[303] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__584__A _584_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[68\] _532_/Y la_data_in_core[68] la_buf\[68\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[101\]_A input262/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2041 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_700 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[124\] _588_/Y la_data_in_core[124] la_buf\[124\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_2181 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output712_A output712/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[57\] user_to_mprj_in_gates\[57\]/Y user_to_mprj_in_gates\[57\]/B
+ input84/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_19_361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__494__A _494_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[119\]_A input25/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_419 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1807 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[124\]_TE mprj_logic_high_inst/HI[326] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_136 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_169 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[90\]_A input377/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1693 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input276_A la_iena_mprj[114] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1177 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__579__A _579_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input443_A la_oenb_mprj[34] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2310 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput320 vccd vssd la_iena_mprj[39] input320/X vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1929 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[23\]_TE mprj_logic_high_inst/HI[225] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xinput331 vssd vccd input331/X la_iena_mprj[49] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput342 vssd vccd input342/X la_iena_mprj[59] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput353 vssd vccd input353/X la_iena_mprj[69] vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_input610_A mprj_dat_o_core[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput364 vssd vccd input364/X la_iena_mprj[79] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput375 vssd vccd input375/X la_iena_mprj[89] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput386 vssd vccd input386/X la_iena_mprj[99] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput397 vccd vssd _371_/A la_oenb_mprj[108] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_48_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[81\]_A input367/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_161 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2261 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_597_ _597_/A _597_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_32_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2169 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[27\] user_to_mprj_in_gates\[27\]/Y output674/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output662_A output662/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1181 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1788 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__489__A _489_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[72\]_A input357/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1989 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_18 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_29 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2069 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[8\]_B la_buf_enable\[8\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_1699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[61\]_TE la_buf\[61\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1866 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[46\]_TE mprj_logic_high_inst/HI[248] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__399__A _399_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[94\]_A_N _357_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[67\] vccd vssd user_to_mprj_in_gates\[67\]/B mprj_logic_high_inst/HI[397]
+ input351/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_24_1659 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_607 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_520_ _520_/Y _520_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_6_1580 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[63\]_A input347/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[5\] _597_/Y la_oenb_core[5] mprj_logic_high_inst/HI[207]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[23\] _615_/Y la_oenb_core[23] mprj_logic_high_inst/HI[225]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_451_ _451_/Y _451_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_4
XFILLER_32_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[45\] la_buf\[45\]/TE _637_/A la_buf_enable\[45\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_25_150 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_382_ _382_/Y _382_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf_enable\[32\]_A_N _624_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1001 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input393_A la_oenb_mprj[104] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input87_A la_data_out_core[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[47\]_A_N _639_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input560_A mprj_dat_i_user[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[10\]_TE mprj_dat_buf\[10\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_721 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_irq_gates\[1\]_B user_irq_gates\[1\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_916 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput172 vccd vssd la_data_out_mprj[20] _484_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput150 la_data_out_mprj[116] _580_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput161 la_data_out_mprj[126] _590_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput194 la_data_out_mprj[40] _504_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput183 la_data_out_mprj[30] _494_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_ena_buf\[54\]_A input337/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_429 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
X_649_ _649_/A _649_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_38_2080 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_632 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1811 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1975 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[84\]_TE la_buf\[84\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[69\]_TE mprj_logic_high_inst/HI[271] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xoutput635 vccd vssd la_data_in_mprj[107] output635/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput668 vccd vssd la_data_in_mprj[21] output668/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput679 vccd vssd la_data_in_mprj[31] output679/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput646 vccd vssd la_data_in_mprj[117] output646/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput657 vccd vssd la_data_in_mprj[127] output657/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_45_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1935 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1225 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[2\]_A _398_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_949 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_437 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[45\]_A input327/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_481 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_665 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2077 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1354 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_359 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2293 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2135 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xmprj_dat_buf\[19\] _451_/Y mprj_dat_o_user[19] mprj_dat_buf\[19\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_24_2179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input239_A la_data_out_mprj[81] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input141_A la_data_out_mprj[108] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1675 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1528 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[36\]_A input317/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1230 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input406_A la_oenb_mprj[116] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_503_ _503_/Y _503_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_26_470 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1296 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_434_ _434_/A _434_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_35_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[50\] _514_/Y la_data_in_core[50] la_buf\[50\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__592__A _592_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2106 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_365_ _365_/A _365_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[122\] vccd vssd user_to_mprj_in_gates\[122\]/B mprj_logic_high_inst/HI[452]
+ input285/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_14_687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2297 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[3\]_A _435_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_842 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_886 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[14\] _414_/Y mprj_adr_o_user[14] mprj_adr_buf\[14\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_29_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[40\]_B user_to_mprj_in_gates\[40\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[94\] user_to_mprj_in_gates\[94\]/Y output748/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_49_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[27\]_A input307/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_749 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_buffers\[4\] output782/A user_wb_dat_gates\[4\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_51_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1794 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[31\]_B user_to_mprj_in_gates\[31\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[1\] user_to_mprj_in_gates\[1\]/Y user_to_mprj_in_gates\[1\]/B
+ input43/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_buffers\[92\]_A user_to_mprj_in_gates\[92\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1787 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[18\]_A input297/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[98\]_B user_to_mprj_in_gates\[98\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input189_A la_data_out_mprj[36] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[90\] _353_/Y la_oenb_core[90] mprj_logic_high_inst/HI[292]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[22\]_B user_to_mprj_in_gates\[22\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input356_A la_iena_mprj[71] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[83\]_A user_to_mprj_in_gates\[83\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_3_878 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1832 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[98\] _562_/Y la_data_in_core[98] la_buf\[98\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[3\] vccd vssd user_to_mprj_in_gates\[3\]/B mprj_logic_high_inst/HI[333]
+ input321/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_input523_A mprj_adr_o_core[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__587__A _587_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[113\] la_buf\[113\]/TE _376_/A la_buf_enable\[113\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_19_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2326 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[89\]_B user_to_mprj_in_gates\[89\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1093 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_417_ _417_/Y _417_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_6
X_348_ _348_/A _348_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_15_1923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_495 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1847 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[121\]_A user_to_mprj_in_gates\[121\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output742_A output742/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[110\]_A _574_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[13\]_B user_to_mprj_in_gates\[13\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[74\]_A user_to_mprj_in_gates\[74\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1629 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[87\] user_to_mprj_in_gates\[87\]/Y user_to_mprj_in_gates\[87\]/B
+ input117/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_42_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__497__A _497_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[24\]_TE mprj_adr_buf\[24\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_705 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1870 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2161 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[112\]_A user_to_mprj_in_gates\[112\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_498 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[101\]_A _565_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[65\]_A user_to_mprj_in_gates\[65\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1117 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2252 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_329 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_543 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1901 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_727 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input104_A la_data_out_core[75] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1967 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[1\] user_to_mprj_in_gates\[1\]/Y output666/A vccd vssd vssd
+ vccd sky130_fd_sc_hd__clkinv_4
XFILLER_23_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_410 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_62 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_443 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1533 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input473_A la_oenb_mprj[61] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[103\]_A user_to_mprj_in_gates\[103\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[13\] _477_/Y la_data_in_core[13] la_buf\[13\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf\[9\] _473_/Y la_data_in_core[9] la_buf\[9\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_48_1017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[56\]_A user_to_mprj_in_gates\[56\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2027 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[6\] _406_/Y mprj_adr_o_user[6] mprj_adr_buf\[6\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_47_830 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1280 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_554 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[57\] user_to_mprj_in_gates\[57\]/Y output707/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_37_2167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2009 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_579 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[96\]_A _560_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output692_A output692/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1731 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[15\] user_wb_dat_gates\[15\]/Y input556/X user_wb_ack_gate/B vssd
+ vccd vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_50_1633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1021 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_785 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1677 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1054 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_981 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[47\]_A user_to_mprj_in_gates\[47\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[12\] output759/A user_wb_dat_gates\[12\]/Y vssd vccd vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_2127 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[20\]_A _484_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[113\] user_to_mprj_in_gates\[113\]/Y user_to_mprj_in_gates\[113\]/B
+ input19/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_9_1099 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1194 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[18\]_TE la_buf\[18\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[87\]_A _551_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[110\]_B mprj_logic_high_inst/HI[440] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[97\] vccd vssd user_to_mprj_in_gates\[97\]/B mprj_logic_high_inst/HI[427]
+ input384/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_49_1337 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[38\]_A user_to_mprj_in_gates\[38\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[123\] _386_/Y la_oenb_core[123] mprj_logic_high_inst/HI[325]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[11\]_A _475_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput502 vccd vssd _351_/A la_oenb_mprj[88] vssd vccd sky130_fd_sc_hd__buf_4
Xuser_to_mprj_oen_buffers\[53\] _645_/Y la_oenb_core[53] mprj_logic_high_inst/HI[255]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xinput513 _361_/A la_oenb_mprj[98] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput546 mprj_adr_o_core[7] _407_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput524 vccd vssd _416_/A mprj_adr_o_core[16] vssd vccd sky130_fd_sc_hd__buf_2
Xinput535 _426_/A mprj_adr_o_core[26] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput557 input557/X mprj_dat_i_user[16] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_16
Xinput579 mprj_dat_i_user[7] input579/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
Xinput568 mprj_dat_i_user[26] input568/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[75\] la_buf\[75\]/TE _338_/A la_buf_enable\[75\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_40_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input319_A la_iena_mprj[38] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input221_A la_data_out_mprj[65] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1453 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_844 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[78\]_A _542_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[101\]_B mprj_logic_high_inst/HI[431] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input590_A mprj_dat_o_core[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[96\]_B la_buf_enable\[96\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_712 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_277 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[117\] _581_/Y la_data_in_core[117] la_buf\[117\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[29\]_A user_to_mprj_in_gates\[29\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_4_962 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[110\] user_to_mprj_in_gates\[110\]/Y output639/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf_enable\[20\]_B la_buf_enable\[20\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output705_A output705/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[119\]_B user_to_mprj_in_gates\[119\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[69\]_A _533_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[120\]_A_N _383_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[87\]_B la_buf_enable\[87\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1138 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1485 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1933 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[28\]_A input570/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[11\]_B la_buf_enable\[11\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1819 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_148 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1565 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[9\]_TE la_buf\[9\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[90\]_B mprj_logic_high_inst/HI[420] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[12\] vccd vssd user_to_mprj_in_gates\[12\]/B mprj_logic_high_inst/HI[342]
+ input291/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_la_buf_enable\[78\]_B la_buf_enable\[78\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2340 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[80\]_A _343_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input171_A la_data_out_mprj[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input269_A la_iena_mprj[108] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[19\]_A input560/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input436_A la_oenb_mprj[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput321 vccd vssd la_iena_mprj[3] input321/X vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput310 vssd vccd input310/X la_iena_mprj[2] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1504 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1537 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input32_A la_data_out_core[125] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_413 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xinput354 la_iena_mprj[6] input354/X vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput343 vccd vssd input343/X la_iena_mprj[5] vssd vccd sky130_fd_sc_hd__buf_2
Xinput332 vccd vssd input332/X la_iena_mprj[4] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_48_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[80\] _544_/Y la_data_in_core[80] la_buf\[80\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xinput376 input376/X la_iena_mprj[8] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput365 input365/X la_iena_mprj[7] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput387 vccd vssd input387/X la_iena_mprj[9] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input603_A mprj_dat_o_core[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__595__A _595_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput398 _372_/A la_oenb_mprj[109] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_28_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1147 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[81\]_B mprj_logic_high_inst/HI[411] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
X_596_ _596_/A _596_/Y vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_32_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_803 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[69\]_B la_buf_enable\[69\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1425 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[71\]_A _334_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_575 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output655_A output655/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2233 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1229 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1491 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_413 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1852 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_19 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[72\]_B mprj_logic_high_inst/HI[402] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_357 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1970 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[62\]_A _654_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[127\]_A _390_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1299 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1592 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[63\]_B mprj_logic_high_inst/HI[393] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
X_450_ _450_/Y _450_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_4
Xuser_to_mprj_oen_buffers\[16\] _608_/Y la_oenb_core[16] mprj_logic_high_inst/HI[218]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
X_381_ _381_/A _381_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_25_162 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[38\] la_buf\[38\]/TE _630_/A la_buf_enable\[38\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_40_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1057 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input386_A la_iena_mprj[99] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[53\]_A _645_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[118\]_A _381_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input553_A mprj_dat_i_user[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2013 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_740 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_777 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput140 _571_/A la_data_out_mprj[107] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput151 _581_/A la_data_out_mprj[117] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput162 vccd vssd _591_/A la_data_out_mprj[127] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_48_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput195 la_data_out_mprj[41] _505_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput173 la_data_out_mprj[21] _485_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput184 la_data_out_mprj[31] _495_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1389 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[54\]_B mprj_logic_high_inst/HI[384] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
X_648_ _648_/Y _648_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_36_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2092 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
X_579_ _579_/Y _579_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_output772_A output772/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[114\]_TE mprj_logic_high_inst/HI[316] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1987 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[109\]_A _372_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[44\]_A _636_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_383 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput636 vccd vssd la_data_in_mprj[108] output636/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput658 vccd vssd la_data_in_mprj[12] output658/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput669 vccd vssd la_data_in_mprj[22] output669/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput647 vccd vssd la_data_in_mprj[118] output647/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_28_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[45\]_B mprj_logic_high_inst/HI[375] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_600 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1366 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_327 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[13\]_TE mprj_logic_high_inst/HI[215] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[35\]_A _627_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1642 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1593 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[31\]_A _431_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input134_A la_data_out_mprj[101] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[36\]_B mprj_logic_high_inst/HI[366] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_18_427 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1220 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input301_A la_iena_mprj[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_502_ _502_/A _502_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
X_433_ _433_/A _433_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_41_441 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2265 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_364_ _364_/Y _364_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf\[43\] _507_/Y la_data_in_core[43] la_buf\[43\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_31_2118 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[115\] vccd vssd user_to_mprj_in_gates\[115\]/B mprj_logic_high_inst/HI[445]
+ input277/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[26\]_A _618_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_854 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1925 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2361 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_11 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1407 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1568 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[87\] user_to_mprj_in_gates\[87\]/Y output740/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_mprj_adr_buf\[22\]_A _422_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[51\]_TE la_buf\[51\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[27\]_B mprj_logic_high_inst/HI[357] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_51_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[32\] user_to_mprj_in_gates\[32\]/Y user_to_mprj_in_gates\[32\]/B
+ input57/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_51_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[36\]_TE mprj_logic_high_inst/HI[238] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[93\]_A_N _356_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[17\]_A _609_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1085 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1659 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[31\]_A_N _623_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1001 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2241 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[13\]_A _413_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[46\]_A_N _638_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_213 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[18\]_B mprj_logic_high_inst/HI[348] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1141 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[83\] _346_/Y la_oenb_core[83] mprj_logic_high_inst/HI[285]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[31\] _463_/Y mprj_dat_o_user[31] mprj_dat_buf\[31\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_5_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_334 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input349_A la_iena_mprj[65] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input251_A la_data_out_mprj[92] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1844 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2027 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input516_A mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[74\]_TE la_buf\[74\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[106\] la_buf\[106\]/TE _369_/A la_buf_enable\[106\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_19_725 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[59\]_TE mprj_logic_high_inst/HI[261] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2338 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_205 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1615 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_416_ _416_/A _416_/Y vssd vccd vssd vccd sky130_fd_sc_hd__inv_12
X_347_ _347_/A _347_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_35_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1935 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1225 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output735_A output735/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1365 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[23\]_TE mprj_dat_buf\[23\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[2\]_TE mprj_logic_high_inst/HI[204] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[97\]_TE la_buf\[97\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_2264 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_555 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[42\] vccd vssd user_to_mprj_in_gates\[42\]/B mprj_logic_high_inst/HI[372]
+ input324/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_38_1924 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[20\] la_buf\[20\]/TE _612_/A la_buf_enable\[20\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_23_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input299_A la_iena_mprj[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_74 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input62_A la_data_out_core[37] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1990 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input466_A la_oenb_mprj[55] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1029 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_120 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2039 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_665 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2353 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__598__A _598_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_197 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_533 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_dat_buf\[26\]_A _458_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output685_A output685/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1645 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1743 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2139 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1850 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1703 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[17\]_A _449_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_1747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2222 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_buffers\[24\]_A user_wb_dat_gates\[24\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_53_823 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_886 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_385 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[106\] user_to_mprj_in_gates\[106\]/Y user_to_mprj_in_gates\[106\]/B
+ input11/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_52_344 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_720 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[116\] _379_/Y la_oenb_core[116] mprj_logic_high_inst/HI[318]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
Xinput503 vccd vssd _352_/A la_oenb_mprj[89] vssd vccd sky130_fd_sc_hd__buf_4
Xinput514 _362_/A la_oenb_mprj[99] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput525 mprj_adr_o_core[17] _417_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput536 vccd vssd _427_/A mprj_adr_o_core[27] vssd vccd sky130_fd_sc_hd__buf_2
Xinput569 mprj_dat_i_user[27] input569/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_8
Xinput558 mprj_dat_i_user[17] input558/X vssd vccd vssd vccd sky130_fd_sc_hd__buf_12
XFILLER_47_105 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1421 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput547 _408_/A mprj_adr_o_core[8] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1590 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[46\] _638_/Y la_oenb_core[46] mprj_logic_high_inst/HI[248]
+ vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_47_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[68\] la_buf\[68\]/TE _331_/A la_buf_enable\[68\]/B vssd vccd vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_28_341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1869 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input214_A la_data_out_mprj[59] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[15\]_A user_wb_dat_gates\[15\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_16_503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input583_A mprj_dat_o_core[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_234 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[14\]_TE mprj_adr_buf\[14\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1651 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_974 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[103\] user_to_mprj_in_gates\[103\]/Y output631/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_43_1493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_650 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1885 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_790 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1901 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[28\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[2\] _434_/Y mprj_dat_o_user[2] mprj_dat_buf\[2\]/TE vccd vssd vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[2\]_TE mprj_dat_buf\[2\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2306 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_193 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[110\]_B la_buf_enable\[110\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[122\]_TE la_buf\[122\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_561 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1673 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_buffers\[1\]_A user_wb_dat_gates\[1\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1113 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2167 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_97 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input164_A la_data_out_mprj[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[19\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput300 vssd vccd input300/X la_iena_mprj[20] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput311 vssd vccd input311/X la_iena_mprj[30] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_49_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input331_A la_iena_mprj[49] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput333 vssd vccd input333/X la_iena_mprj[50] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput322 vssd vccd input322/X la_iena_mprj[40] vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_input429_A la_oenb_mprj[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput344 vssd vccd input344/X la_iena_mprj[60] vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_1_999 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input25_A la_data_out_core[119] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_469 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput388 la_oenb_mprj[0] _592_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput355 vssd vccd input355/X la_iena_mprj[70] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput366 vssd vccd input366/X la_iena_mprj[80] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput377 vssd vccd input377/X la_iena_mprj[90] vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput399 la_oenb_mprj[10] _602_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_la_buf\[4\]_A _468_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[73\] _537_/Y la_data_in_core[73] la_buf\[73\]/TE vccd vssd vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[101\]_B la_buf_enable\[101\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_595_ _595_/A _595_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[70\]_A input99/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output648_A output648/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1037 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[62\] user_to_mprj_in_gates\[62\]/Y user_to_mprj_in_gates\[62\]/B
+ input90/X vssd vccd vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_48_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1864 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_653 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_193 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1050 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1802 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_892 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1982 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[61\]_A input89/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_2307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1847 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_992 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_380_ _380_/A _380_/Y vccd vssd vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[92\]_TE mprj_logic_high_inst/HI[294] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_133 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input281_A la_iena_mprj[119] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input379_A la_iena_mprj[92] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[52\]_A input79/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input546_A mprj_adr_o_core[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput130 vccd vssd input130/X la_data_out_core[99] vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_48_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput163 la_data_out_mprj[12] _476_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput141 _572_/A la_data_out_mprj[108] vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput152 la_data_out_mprj[118] _582_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_48_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_417 vccd vssd vssd vccd sky130_fd_sc_hd__decap_3
Xinput196 la_data_out_mprj[42] _506_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput174 la_data_out_mprj[22] _486_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput185 la_data_out_mprj[32] _496_/A vssd vccd vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_40_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_647_ _647_/Y _647_/A vccd vssd vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_601 vccd vssd vssd vccd sky130_fd_sc_hd__decap_6
X_578_ _578_/Y _578_/A vccd vssd vssd vccd sky130_fd_sc_hd__inv_4
XFILLER_32_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[2\]_A user_to_mprj_in_gates\[2\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[32\] user_to_mprj_in_gates\[32\]/Y output680/A vccd vssd
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output765_A output765/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_874 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[43\]_A input69/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput659 vccd vssd la_data_in_mprj[13] output659/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput637 vccd vssd la_data_in_mprj[109] output637/A vssd vccd sky130_fd_sc_hd__buf_2
Xoutput648 vccd vssd la_data_in_mprj[119] output648/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_45_2053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2097 vccd vssd vssd vccd sky130_fd_sc_hd__decap_8
.ends

